
module inc_by_2(A, Out);
    input [15:0] A;
    output [15:0] Out;

    

endmodule
