
module fulladder1_15 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4;

  INVX1 U1 ( .A(n4), .Y(n1) );
  INVX4 U2 ( .A(n2), .Y(n3) );
  INVX1 U3 ( .A(B), .Y(n2) );
  INVX1 U4 ( .A(A), .Y(n4) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U6 ( .A(n3), .B(n4), .Y(P) );
  FAX1 U7 ( .A(Cin), .B(n1), .C(n3), .YC(), .YS(S) );
endmodule


module fulladder1_14 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(n6), .Y(n3) );
  INVX1 U4 ( .A(n6), .Y(n4) );
  INVX1 U5 ( .A(A), .Y(n6) );
  XOR2X1 U6 ( .A(n2), .B(n4), .Y(n5) );
  XOR2X1 U7 ( .A(Cin), .B(n5), .Y(S) );
  AND2X2 U8 ( .A(B), .B(n3), .Y(G) );
  XNOR2X1 U9 ( .A(B), .B(n6), .Y(P) );
endmodule


module fulladder1_13 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n7;

  INVX1 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(A), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  BUFX2 U5 ( .A(P), .Y(n5) );
  INVX1 U6 ( .A(n7), .Y(P) );
  AND2X2 U7 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U8 ( .A(n4), .B(n2), .Y(n7) );
  XOR2X1 U9 ( .A(Cin), .B(n5), .Y(S) );
endmodule


module fulladder1_12 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n6;

  BUFX4 U1 ( .A(B), .Y(n4) );
  XOR2X1 U2 ( .A(n4), .B(A), .Y(P) );
  BUFX2 U3 ( .A(n4), .Y(n1) );
  INVX1 U4 ( .A(A), .Y(n6) );
  BUFX2 U5 ( .A(n6), .Y(n2) );
  INVX1 U6 ( .A(n6), .Y(n3) );
  XNOR2X1 U7 ( .A(Cin), .B(n5), .Y(S) );
  XOR2X1 U8 ( .A(n1), .B(n2), .Y(n5) );
  AND2X2 U9 ( .A(B), .B(n3), .Y(G) );
endmodule


module fulladder1_11 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3;

  XOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX8 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(P), .Y(n2) );
  INVX1 U4 ( .A(n3), .Y(P) );
  AND2X2 U5 ( .A(B), .B(A), .Y(G) );
  XNOR2X1 U6 ( .A(B), .B(A), .Y(n3) );
endmodule


module fulladder1_10 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3, n4, n5;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  XOR2X1 U2 ( .A(n4), .B(n5), .Y(n1) );
  XOR2X1 U3 ( .A(B), .B(A), .Y(P) );
  BUFX2 U4 ( .A(A), .Y(n3) );
  BUFX2 U5 ( .A(B), .Y(n4) );
  INVX1 U6 ( .A(n3), .Y(n5) );
  AND2X2 U7 ( .A(B), .B(A), .Y(G) );
endmodule


module fulladder1_9 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3;

  XOR2X1 U1 ( .A(B), .B(A), .Y(P) );
  BUFX2 U2 ( .A(P), .Y(n2) );
  XNOR2X1 U3 ( .A(Cin), .B(n3), .Y(S) );
  INVX1 U4 ( .A(n2), .Y(n3) );
  AND2X2 U5 ( .A(B), .B(A), .Y(G) );
endmodule


module fulladder1_8 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3;

  INVX1 U1 ( .A(n3), .Y(n1) );
  XNOR2X1 U2 ( .A(n2), .B(n1), .Y(S) );
  INVX1 U3 ( .A(Cin), .Y(n2) );
  XNOR2X1 U4 ( .A(B), .B(A), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(P) );
  AND2X2 U6 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_7 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XNOR2X1 U1 ( .A(Cin), .B(n2), .Y(S) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  INVX1 U3 ( .A(P), .Y(n2) );
  AND2X2 U4 ( .A(B), .B(A), .Y(G) );
endmodule


module fulladder1_6 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n6, n7;

  BUFX2 U1 ( .A(n5), .Y(n1) );
  XNOR2X1 U2 ( .A(B), .B(n5), .Y(P) );
  XNOR2X1 U3 ( .A(Cin), .B(n7), .Y(S) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(B), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  INVX1 U7 ( .A(A), .Y(n5) );
  INVX1 U8 ( .A(n1), .Y(n6) );
  XOR2X1 U9 ( .A(n4), .B(n1), .Y(n7) );
  AND2X2 U10 ( .A(n2), .B(n6), .Y(G) );
endmodule


module fulladder1_5 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  XOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  XNOR2X1 U2 ( .A(B), .B(n2), .Y(n1) );
  XOR2X1 U3 ( .A(B), .B(A), .Y(P) );
  INVX1 U4 ( .A(A), .Y(n2) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_4 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3, n4;

  INVX1 U1 ( .A(A), .Y(n3) );
  BUFX2 U2 ( .A(P), .Y(n1) );
  XNOR2X1 U3 ( .A(B), .B(n3), .Y(P) );
  XNOR2X1 U4 ( .A(n4), .B(n1), .Y(S) );
  INVX1 U5 ( .A(Cin), .Y(n4) );
  AND2X2 U6 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_3 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n4, n5, n6, n7, n8, n9;

  XOR2X1 U1 ( .A(B), .B(A), .Y(P) );
  AND2X2 U2 ( .A(n7), .B(n5), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(S) );
  AND2X2 U4 ( .A(Cin), .B(n9), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(n5) );
  AND2X2 U6 ( .A(n8), .B(P), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  INVX1 U8 ( .A(Cin), .Y(n8) );
  INVX1 U9 ( .A(P), .Y(n9) );
  AND2X2 U10 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_2 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  XOR2X1 U1 ( .A(n1), .B(n3), .Y(S) );
  INVX1 U2 ( .A(Cin), .Y(n1) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  INVX1 U4 ( .A(P), .Y(n3) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_1 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3;

  XOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX8 U2 ( .A(n2), .Y(n1) );
  BUFX2 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(n3), .Y(P) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U6 ( .A(A), .B(B), .Y(n3) );
endmodule


module fulladder1_0 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U2 ( .A(n1), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n1) );
endmodule


module demux1to4_17 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n14, n16;

  INVX1 U1 ( .A(\S<1> ), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  OR2X2 U3 ( .A(n8), .B(n2), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out1) );
  OR2X2 U5 ( .A(\S<0> ), .B(n2), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(\S<0> ), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  INVX1 U11 ( .A(n9), .Y(n11) );
  OR2X2 U12 ( .A(n10), .B(n16), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(Out3) );
  OR2X2 U14 ( .A(n11), .B(\S<0> ), .Y(n14) );
  INVX1 U15 ( .A(n14), .Y(Out2) );
  AND2X2 U16 ( .A(In), .B(n6), .Y(Out0) );
  INVX1 U17 ( .A(\S<0> ), .Y(n16) );
endmodule


module demux1to4_18 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  OR2X2 U1 ( .A(n13), .B(n15), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n12), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n10), .B(n14), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  OR2X2 U7 ( .A(\S<0> ), .B(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(\S<0> ), .B(In), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  AND2X2 U11 ( .A(In), .B(n14), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(n11), .Y(n13) );
  BUFX2 U14 ( .A(\S<1> ), .Y(n14) );
  AND2X2 U15 ( .A(n8), .B(In), .Y(Out0) );
  INVX1 U16 ( .A(\S<0> ), .Y(n15) );
endmodule


module demux1to4_19 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n13, n15;

  INVX1 U1 ( .A(n15), .Y(n1) );
  OR2X2 U2 ( .A(n10), .B(n15), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(\S<1> ), .B(\S<0> ), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(n5) );
  AND2X2 U6 ( .A(n1), .B(In), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(\S<1> ), .B(In), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  INVX1 U10 ( .A(n8), .Y(n10) );
  OR2X2 U11 ( .A(n9), .B(n1), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(Out2) );
  OR2X2 U13 ( .A(n7), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out1) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
  AND2X2 U16 ( .A(n5), .B(In), .Y(Out0) );
endmodule


module demux1to4_20 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n14;

  OR2X2 U1 ( .A(n11), .B(n14), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n10), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(\S<0> ), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(\S<0> ), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(In), .B(\S<1> ), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  INVX1 U11 ( .A(n9), .Y(n11) );
  OR2X2 U12 ( .A(n8), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(Out1) );
  AND2X2 U14 ( .A(In), .B(n6), .Y(Out0) );
  INVX1 U15 ( .A(\S<0> ), .Y(n14) );
endmodule


module demux1to4_21 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n12, n13, n14;

  OR2X2 U1 ( .A(n9), .B(n14), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n8), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  AND2X2 U5 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(\S<1> ), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  INVX1 U9 ( .A(n7), .Y(n9) );
  AND2X1 U10 ( .A(In), .B(n13), .Y(n12) );
  OR2X2 U11 ( .A(n6), .B(\S<1> ), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(Out1) );
  AND2X2 U13 ( .A(n14), .B(n12), .Y(Out0) );
  INVX1 U14 ( .A(\S<1> ), .Y(n13) );
  INVX1 U15 ( .A(\S<0> ), .Y(n14) );
endmodule


module demux1to4_22 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18;

  AND2X2 U1 ( .A(In), .B(n17), .Y(n7) );
  OR2X2 U2 ( .A(n8), .B(\S<0> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out0) );
  OR2X2 U4 ( .A(n12), .B(\S<0> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out2) );
  OR2X2 U6 ( .A(n10), .B(\S<1> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out1) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(\S<0> ), .B(n14), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  AND2X2 U11 ( .A(\S<1> ), .B(n14), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(n11), .Y(n13) );
  BUFX2 U14 ( .A(In), .Y(n14) );
  OR2X2 U15 ( .A(n13), .B(n18), .Y(n15) );
  INVX1 U16 ( .A(n15), .Y(Out3) );
  INVX1 U17 ( .A(\S<1> ), .Y(n17) );
  INVX1 U18 ( .A(\S<0> ), .Y(n18) );
endmodule


module demux1to4_23 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n14;

  OR2X2 U1 ( .A(n11), .B(n14), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n10), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(\S<0> ), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(\S<0> ), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(In), .B(\S<1> ), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  INVX1 U11 ( .A(n9), .Y(n11) );
  OR2X2 U12 ( .A(n8), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(Out1) );
  AND2X2 U14 ( .A(In), .B(n6), .Y(Out0) );
  INVX1 U15 ( .A(\S<0> ), .Y(n14) );
endmodule


module demux1to4_24 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20;

  AND2X1 U1 ( .A(In), .B(n19), .Y(n11) );
  OR2X2 U2 ( .A(\S<0> ), .B(n12), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out0) );
  OR2X2 U4 ( .A(n15), .B(n20), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out3) );
  OR2X2 U6 ( .A(n14), .B(\S<0> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out2) );
  OR2X2 U8 ( .A(n10), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  AND2X2 U10 ( .A(\S<0> ), .B(n18), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(n10) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  AND2X2 U13 ( .A(\S<1> ), .B(n16), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(n14) );
  INVX1 U15 ( .A(n13), .Y(n15) );
  INVX1 U16 ( .A(n17), .Y(n16) );
  INVX1 U17 ( .A(In), .Y(n17) );
  INVX1 U18 ( .A(n17), .Y(n18) );
  INVX1 U19 ( .A(\S<1> ), .Y(n19) );
  INVX1 U20 ( .A(\S<0> ), .Y(n20) );
endmodule


module demux1to4_25 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n14;

  OR2X2 U1 ( .A(\S<0> ), .B(\S<1> ), .Y(n10) );
  OR2X2 U2 ( .A(n9), .B(n14), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X2 U4 ( .A(n6), .B(\S<1> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out1) );
  AND2X2 U6 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  AND2X2 U8 ( .A(\S<1> ), .B(In), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(n8) );
  INVX1 U10 ( .A(n7), .Y(n9) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  OR2X2 U12 ( .A(n8), .B(\S<0> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(Out2) );
  INVX1 U14 ( .A(\S<0> ), .Y(n14) );
  AND2X2 U15 ( .A(n11), .B(In), .Y(Out0) );
endmodule


module demux1to4_26 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n5, n6, n8, n10, n11, n12, n13, n14, n16;

  INVX1 U1 ( .A(n16), .Y(n1) );
  OR2X2 U2 ( .A(n14), .B(n16), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(\S<0> ), .B(\S<1> ), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(n5) );
  OR2X2 U6 ( .A(n13), .B(n1), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(Out2) );
  OR2X2 U8 ( .A(n11), .B(\S<1> ), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(Out1) );
  AND2X2 U10 ( .A(In), .B(n1), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  AND2X2 U12 ( .A(In), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(n13) );
  INVX1 U14 ( .A(n12), .Y(n14) );
  AND2X2 U15 ( .A(n5), .B(In), .Y(Out0) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
endmodule


module demux1to4_27 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14;

  OR2X2 U1 ( .A(n10), .B(n14), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n11), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n8), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  AND2X2 U7 ( .A(\S<0> ), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(\S<1> ), .B(In), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  INVX1 U11 ( .A(n9), .Y(n11) );
  OR2X2 U12 ( .A(\S<0> ), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(n13) );
  AND2X2 U14 ( .A(n13), .B(In), .Y(Out0) );
  INVX1 U15 ( .A(\S<0> ), .Y(n14) );
endmodule


module demux1to4_28 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n12, n13, n14;

  OR2X2 U1 ( .A(n8), .B(n14), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n9), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  AND2X2 U5 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(In), .B(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  INVX1 U9 ( .A(n7), .Y(n9) );
  OR2X2 U10 ( .A(n6), .B(\S<1> ), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(Out1) );
  AND2X2 U12 ( .A(n14), .B(n12), .Y(Out0) );
  AND2X1 U13 ( .A(In), .B(n13), .Y(n12) );
  INVX1 U14 ( .A(\S<1> ), .Y(n13) );
  INVX1 U15 ( .A(\S<0> ), .Y(n14) );
endmodule


module demux1to4_29 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n15, n16;

  OR2X2 U1 ( .A(n11), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n10), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  AND2X2 U5 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(n16), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(In), .B(\S<1> ), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  INVX1 U11 ( .A(n9), .Y(n11) );
  OR2X2 U12 ( .A(n6), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(Out1) );
  INVX4 U14 ( .A(n15), .Y(Out0) );
  OR2X2 U15 ( .A(n8), .B(\S<1> ), .Y(n15) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
endmodule


module demux1to4_30 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n16;

  OR2X2 U1 ( .A(n14), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n13), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n9), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  OR2X2 U7 ( .A(n11), .B(\S<1> ), .Y(n7) );
  AND2X2 U8 ( .A(\S<0> ), .B(In), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(n16), .B(In), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  AND2X2 U12 ( .A(In), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(n13) );
  INVX1 U14 ( .A(n12), .Y(n14) );
  INVX4 U15 ( .A(n7), .Y(Out0) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
endmodule


module demux1to4_31 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n16;

  OR2X2 U1 ( .A(n14), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n13), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n9), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  OR2X2 U7 ( .A(n11), .B(\S<1> ), .Y(n7) );
  AND2X2 U8 ( .A(\S<0> ), .B(In), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(In), .B(n16), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  AND2X2 U12 ( .A(In), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(n13) );
  INVX1 U14 ( .A(n12), .Y(n14) );
  INVX4 U15 ( .A(n7), .Y(Out0) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
endmodule


module demux1to4_32 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n11, n12, n13, n14, n16;

  OR2X2 U1 ( .A(n12), .B(\S<0> ), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out2) );
  OR2X2 U3 ( .A(n6), .B(\S<1> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out1) );
  AND2X2 U5 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(n16), .B(In), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  OR2X2 U9 ( .A(n13), .B(n16), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(Out3) );
  AND2X2 U11 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(n11), .Y(n13) );
  OR2X2 U14 ( .A(n8), .B(\S<1> ), .Y(n14) );
  INVX1 U15 ( .A(n14), .Y(Out0) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
endmodule


module demux1to4_15 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17;

  INVX1 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  BUFX2 U3 ( .A(\S<0> ), .Y(n3) );
  OR2X2 U4 ( .A(n14), .B(n17), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out3) );
  OR2X2 U6 ( .A(n13), .B(n3), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(Out2) );
  OR2X2 U8 ( .A(\S<1> ), .B(\S<0> ), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(n3), .B(n2), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  AND2X2 U12 ( .A(n2), .B(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n12), .Y(n13) );
  INVX1 U14 ( .A(n12), .Y(n14) );
  OR2X2 U15 ( .A(n11), .B(\S<1> ), .Y(n15) );
  INVX1 U16 ( .A(n15), .Y(Out1) );
  INVX1 U17 ( .A(\S<0> ), .Y(n17) );
  AND2X2 U18 ( .A(n9), .B(In), .Y(Out0) );
endmodule


module demux1to4_14 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  OR2X2 U1 ( .A(n13), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n12), .B(n15), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n10), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  OR2X2 U7 ( .A(\S<1> ), .B(\S<0> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(n15), .B(n14), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  AND2X2 U11 ( .A(\S<1> ), .B(n14), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(n11), .Y(n13) );
  INVX1 U14 ( .A(\S<0> ), .Y(n16) );
  BUFX2 U15 ( .A(In), .Y(n14) );
  INVX1 U16 ( .A(n16), .Y(n15) );
  AND2X2 U17 ( .A(In), .B(n8), .Y(Out0) );
endmodule


module demux1to4_13 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  OR2X2 U1 ( .A(n10), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n9), .B(n15), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(\S<1> ), .B(\S<0> ), .Y(n5) );
  AND2X2 U6 ( .A(n15), .B(n11), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(\S<1> ), .B(n11), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  INVX1 U10 ( .A(n8), .Y(n10) );
  BUFX2 U11 ( .A(In), .Y(n11) );
  INVX1 U12 ( .A(n5), .Y(n12) );
  OR2X2 U13 ( .A(n7), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out1) );
  INVX1 U15 ( .A(n16), .Y(n15) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
  AND2X2 U17 ( .A(n12), .B(In), .Y(Out0) );
endmodule


module demux1to4_12 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15;

  BUFX2 U1 ( .A(In), .Y(n1) );
  OR2X2 U2 ( .A(n12), .B(n15), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(n11), .B(\S<0> ), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out2) );
  OR2X2 U6 ( .A(\S<1> ), .B(\S<0> ), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(\S<0> ), .B(n1), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(\S<1> ), .B(n1), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  INVX1 U12 ( .A(n10), .Y(n12) );
  OR2X2 U13 ( .A(n9), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out1) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
  AND2X2 U16 ( .A(n7), .B(In), .Y(Out0) );
endmodule


module demux1to4_11 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  BUFX2 U1 ( .A(In), .Y(n1) );
  OR2X2 U2 ( .A(n12), .B(n16), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(n11), .B(n15), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out2) );
  OR2X2 U6 ( .A(\S<1> ), .B(n15), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(n15), .B(n1), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(\S<1> ), .B(n1), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  INVX1 U12 ( .A(n10), .Y(n12) );
  INVX1 U13 ( .A(n16), .Y(n15) );
  OR2X2 U14 ( .A(n9), .B(\S<1> ), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(Out1) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
  AND2X2 U17 ( .A(In), .B(n7), .Y(Out0) );
endmodule


module demux1to4_10 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  OR2X2 U1 ( .A(n13), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n12), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n10), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  OR2X2 U7 ( .A(\S<1> ), .B(\S<0> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(\S<0> ), .B(n15), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  AND2X2 U11 ( .A(\S<1> ), .B(n15), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(n11), .Y(n13) );
  AND2X2 U14 ( .A(n8), .B(In), .Y(Out0) );
  INVX1 U15 ( .A(\S<0> ), .Y(n16) );
  BUFX2 U16 ( .A(In), .Y(n15) );
endmodule


module demux1to4_9 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  BUFX2 U1 ( .A(In), .Y(n1) );
  OR2X2 U2 ( .A(n12), .B(n15), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(n11), .B(n16), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out2) );
  OR2X2 U6 ( .A(\S<1> ), .B(\S<0> ), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(n16), .B(n1), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(n1), .B(\S<1> ), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  INVX1 U12 ( .A(n10), .Y(n12) );
  OR2X2 U13 ( .A(n9), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out1) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
  INVX1 U16 ( .A(n15), .Y(n16) );
  AND2X2 U17 ( .A(n7), .B(In), .Y(Out0) );
endmodule


module demux1to4_8 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  BUFX2 U1 ( .A(In), .Y(n1) );
  OR2X2 U2 ( .A(n12), .B(n16), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(n11), .B(n15), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out2) );
  OR2X2 U6 ( .A(\S<1> ), .B(n15), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(n15), .B(n1), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(n1), .B(\S<1> ), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  INVX1 U12 ( .A(n10), .Y(n12) );
  OR2X2 U13 ( .A(n9), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out1) );
  INVX1 U15 ( .A(n16), .Y(n15) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
  AND2X2 U17 ( .A(n7), .B(In), .Y(Out0) );
endmodule


module demux1to4_7 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  BUFX2 U1 ( .A(In), .Y(n1) );
  OR2X2 U2 ( .A(n12), .B(n15), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out2) );
  OR2X2 U4 ( .A(n9), .B(\S<1> ), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out1) );
  OR2X2 U6 ( .A(\S<1> ), .B(\S<0> ), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(n15), .B(n1), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(n1), .B(\S<1> ), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  INVX1 U12 ( .A(n10), .Y(n12) );
  INVX1 U13 ( .A(n16), .Y(n15) );
  OR2X2 U14 ( .A(n11), .B(n16), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(Out3) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
  AND2X2 U17 ( .A(In), .B(n7), .Y(Out0) );
endmodule


module demux1to4_6 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n16), .Y(n15) );
  OR2X2 U3 ( .A(n12), .B(n16), .Y(n2) );
  INVX1 U4 ( .A(n2), .Y(Out3) );
  OR2X2 U5 ( .A(n11), .B(n15), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(Out2) );
  OR2X2 U7 ( .A(\S<1> ), .B(\S<0> ), .Y(n6) );
  INVX1 U8 ( .A(n6), .Y(n7) );
  AND2X2 U9 ( .A(n1), .B(n15), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  AND2X2 U11 ( .A(n1), .B(\S<1> ), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(n11) );
  INVX1 U13 ( .A(n10), .Y(n12) );
  OR2X2 U14 ( .A(n9), .B(\S<1> ), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(Out1) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
  AND2X2 U17 ( .A(In), .B(n7), .Y(Out0) );
endmodule


module demux1to4_5 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n6, n7, n8, n9, n10, n11, n12, n13, n15;

  BUFX2 U1 ( .A(In), .Y(n1) );
  OR2X2 U2 ( .A(n12), .B(n15), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(Out3) );
  OR2X2 U4 ( .A(n9), .B(\S<1> ), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(Out1) );
  OR2X2 U6 ( .A(\S<1> ), .B(\S<0> ), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  AND2X2 U8 ( .A(n1), .B(\S<0> ), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  AND2X2 U10 ( .A(n1), .B(\S<1> ), .Y(n10) );
  INVX1 U11 ( .A(n10), .Y(n11) );
  INVX1 U12 ( .A(n10), .Y(n12) );
  OR2X2 U13 ( .A(n11), .B(\S<0> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out2) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
  AND2X2 U16 ( .A(n7), .B(In), .Y(Out0) );
endmodule


module demux1to4_4 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9, n10, n11, n12, n14;

  INVX1 U1 ( .A(\S<0> ), .Y(n14) );
  OR2X2 U2 ( .A(n10), .B(n14), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X2 U4 ( .A(\S<0> ), .B(\S<1> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  OR2X2 U6 ( .A(n11), .B(\S<0> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out2) );
  AND2X2 U8 ( .A(\S<0> ), .B(In), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(n8) );
  AND2X2 U10 ( .A(In), .B(\S<1> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(n10) );
  INVX1 U12 ( .A(n9), .Y(n11) );
  OR2X2 U13 ( .A(n8), .B(\S<1> ), .Y(n12) );
  INVX1 U14 ( .A(n12), .Y(Out1) );
  AND2X2 U15 ( .A(n4), .B(In), .Y(Out0) );
endmodule


module demux1to4_3 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n16;

  OR2X2 U1 ( .A(n13), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n8), .B(\S<1> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out0) );
  OR2X2 U5 ( .A(n12), .B(\S<0> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out2) );
  AND2X2 U7 ( .A(In), .B(n16), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  AND2X2 U9 ( .A(\S<0> ), .B(In), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  AND2X2 U11 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(n11), .Y(n13) );
  INVX1 U14 ( .A(\S<0> ), .Y(n16) );
  OR2X2 U15 ( .A(n10), .B(\S<1> ), .Y(n14) );
  INVX1 U16 ( .A(n14), .Y(Out1) );
endmodule


module demux1to4_2 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16;

  INVX1 U1 ( .A(\S<0> ), .Y(n16) );
  OR2X2 U2 ( .A(n15), .B(n16), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X2 U4 ( .A(n12), .B(\S<1> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out0) );
  OR2X2 U6 ( .A(n14), .B(\S<0> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out2) );
  OR2X2 U8 ( .A(n10), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  AND2X2 U10 ( .A(\S<0> ), .B(In), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(n10) );
  AND2X2 U12 ( .A(n16), .B(In), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(\S<1> ), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(n14) );
  INVX1 U16 ( .A(n13), .Y(n15) );
endmodule


module demux1to4_1 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n16;

  INVX1 U1 ( .A(\S<0> ), .Y(n16) );
  OR2X2 U2 ( .A(n12), .B(n16), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X2 U4 ( .A(n8), .B(\S<1> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out0) );
  OR2X2 U6 ( .A(n13), .B(\S<0> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out2) );
  AND2X2 U8 ( .A(n16), .B(In), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(n8) );
  AND2X2 U10 ( .A(\S<0> ), .B(In), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(n10) );
  AND2X2 U12 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  INVX1 U14 ( .A(n11), .Y(n13) );
  OR2X2 U15 ( .A(n10), .B(\S<1> ), .Y(n14) );
  INVX1 U16 ( .A(n14), .Y(Out1) );
endmodule


module demux1to4_0 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16;

  OR2X2 U1 ( .A(n15), .B(n16), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  OR2X2 U3 ( .A(n14), .B(\S<0> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out2) );
  OR2X2 U5 ( .A(n10), .B(\S<1> ), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out1) );
  OR2X2 U7 ( .A(n12), .B(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(Out0) );
  AND2X2 U9 ( .A(\S<0> ), .B(In), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(n10) );
  AND2X2 U11 ( .A(n16), .B(In), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  AND2X2 U13 ( .A(In), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(n14) );
  INVX1 U15 ( .A(n13), .Y(n15) );
  INVX1 U16 ( .A(\S<0> ), .Y(n16) );
endmodule


module cla4_3 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \C<1> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90;

  fulladder1_15 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n87), .G(n83) );
  fulladder1_14 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(\C<1> ), .S(\S<1> ), 
        .P(n88), .G(n84) );
  fulladder1_13 \fa[2]  ( .A(n65), .B(\B<2> ), .Cin(n49), .S(\S<2> ), .P(n89), 
        .G(n85) );
  fulladder1_12 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n81), .S(\S<3> ), .P(
        n90), .G(n86) );
  INVX1 U1 ( .A(n86), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(n90), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  INVX2 U5 ( .A(n17), .Y(n73) );
  OR2X2 U6 ( .A(n19), .B(n41), .Y(n5) );
  INVX1 U7 ( .A(n82), .Y(n71) );
  XOR2X1 U8 ( .A(n16), .B(n59), .Y(n6) );
  XOR2X1 U9 ( .A(n10), .B(n64), .Y(n7) );
  INVX1 U10 ( .A(n87), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  INVX1 U12 ( .A(n52), .Y(n10) );
  BUFX2 U13 ( .A(n54), .Y(n11) );
  INVX1 U14 ( .A(\B<1> ), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(n13) );
  INVX1 U16 ( .A(n38), .Y(n14) );
  BUFX2 U17 ( .A(n73), .Y(n15) );
  INVX1 U18 ( .A(n67), .Y(n16) );
  INVX1 U19 ( .A(\A<2> ), .Y(n61) );
  BUFX2 U20 ( .A(\A<2> ), .Y(n65) );
  INVX1 U21 ( .A(n83), .Y(n18) );
  NOR3X1 U22 ( .A(n58), .B(n67), .C(n18), .Y(n17) );
  AND2X2 U23 ( .A(\B<2> ), .B(n61), .Y(n19) );
  BUFX2 U24 ( .A(\A<3> ), .Y(n64) );
  AND2X2 U25 ( .A(n88), .B(n70), .Y(n20) );
  BUFX2 U26 ( .A(n69), .Y(n21) );
  AND2X2 U27 ( .A(n44), .B(n42), .Y(n22) );
  INVX1 U28 ( .A(n22), .Y(n23) );
  AND2X2 U29 ( .A(n14), .B(n40), .Y(n24) );
  INVX1 U30 ( .A(n24), .Y(n25) );
  INVX1 U31 ( .A(n20), .Y(n26) );
  OR2X2 U32 ( .A(n54), .B(n72), .Y(n27) );
  INVX1 U33 ( .A(n27), .Y(n28) );
  OR2X2 U34 ( .A(n73), .B(n26), .Y(n29) );
  INVX1 U35 ( .A(n29), .Y(n30) );
  BUFX2 U36 ( .A(n75), .Y(n31) );
  BUFX2 U37 ( .A(n78), .Y(n32) );
  AND2X2 U38 ( .A(n23), .B(n89), .Y(n33) );
  INVX1 U39 ( .A(n33), .Y(n34) );
  AND2X2 U40 ( .A(n7), .B(n6), .Y(n35) );
  INVX1 U41 ( .A(n35), .Y(n36) );
  BUFX2 U42 ( .A(n77), .Y(n37) );
  AND2X2 U43 ( .A(n90), .B(n7), .Y(n38) );
  INVX1 U44 ( .A(n38), .Y(n39) );
  BUFX2 U45 ( .A(n48), .Y(n40) );
  AND2X2 U46 ( .A(n60), .B(\A<2> ), .Y(n41) );
  INVX1 U47 ( .A(n41), .Y(n42) );
  BUFX2 U48 ( .A(n74), .Y(n43) );
  INVX1 U49 ( .A(n19), .Y(n44) );
  INVX1 U50 ( .A(n72), .Y(n45) );
  BUFX2 U51 ( .A(n43), .Y(n46) );
  BUFX2 U52 ( .A(\A<3> ), .Y(n47) );
  XNOR2X1 U53 ( .A(\B<1> ), .B(n55), .Y(n70) );
  NAND3X1 U54 ( .A(n53), .B(n47), .C(n2), .Y(n48) );
  OAI21X1 U55 ( .A(n50), .B(n66), .C(n46), .Y(n49) );
  INVX1 U56 ( .A(n20), .Y(n50) );
  NAND3X1 U57 ( .A(n57), .B(n62), .C(n85), .Y(n51) );
  INVX1 U58 ( .A(\B<3> ), .Y(n52) );
  INVX1 U59 ( .A(n52), .Y(n53) );
  AND2X2 U60 ( .A(n89), .B(n5), .Y(n54) );
  INVX1 U61 ( .A(n11), .Y(n63) );
  INVX1 U62 ( .A(\A<1> ), .Y(n55) );
  INVX1 U63 ( .A(n55), .Y(n56) );
  INVX1 U64 ( .A(n61), .Y(n57) );
  INVX1 U65 ( .A(\A<0> ), .Y(n58) );
  INVX1 U66 ( .A(n58), .Y(n59) );
  INVX1 U67 ( .A(n51), .Y(n72) );
  INVX1 U68 ( .A(\B<2> ), .Y(n60) );
  INVX1 U69 ( .A(n60), .Y(n62) );
  INVX1 U70 ( .A(n66), .Y(\C<1> ) );
  AND2X2 U71 ( .A(n21), .B(n15), .Y(n66) );
  INVX1 U72 ( .A(n81), .Y(n79) );
  INVX1 U73 ( .A(\B<0> ), .Y(n67) );
  BUFX2 U74 ( .A(n40), .Y(n68) );
  NAND3X1 U75 ( .A(Cin), .B(n9), .C(n6), .Y(n69) );
  NAND3X1 U76 ( .A(n56), .B(n13), .C(n84), .Y(n74) );
  OAI21X1 U77 ( .A(n50), .B(n66), .C(n46), .Y(n82) );
  OAI21X1 U78 ( .A(n63), .B(n71), .C(n45), .Y(n81) );
  NAND3X1 U79 ( .A(n47), .B(n53), .C(n86), .Y(n78) );
  NAND3X1 U80 ( .A(n45), .B(n43), .C(n32), .Y(n75) );
  OAI21X1 U81 ( .A(n30), .B(n31), .C(n25), .Y(n76) );
  AOI21X1 U82 ( .A(n68), .B(n28), .C(n76), .Y(GG) );
  NAND3X1 U83 ( .A(n20), .B(n4), .C(n87), .Y(n77) );
  NOR3X1 U84 ( .A(n34), .B(n36), .C(n37), .Y(PG) );
  OAI21X1 U85 ( .A(n39), .B(n79), .C(n68), .Y(Cout) );
endmodule


module cla4_2 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106;

  fulladder1_11 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(n78), .S(\S<0> ), .P(
        n103), .G(n99) );
  fulladder1_10 \fa[1]  ( .A(n76), .B(\B<1> ), .Cin(n13), .S(\S<1> ), .P(n104), 
        .G(n100) );
  fulladder1_9 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n15), .S(\S<2> ), .P(
        n105), .G(n101) );
  fulladder1_8 \fa[3]  ( .A(n65), .B(\B<3> ), .Cin(n98), .S(\S<3> ), .P(n106), 
        .G(n102) );
  OR2X2 U1 ( .A(n89), .B(n90), .Y(n16) );
  INVX1 U2 ( .A(n82), .Y(n1) );
  XNOR2X1 U3 ( .A(\B<2> ), .B(n66), .Y(n2) );
  INVX1 U4 ( .A(n2), .Y(n3) );
  INVX1 U5 ( .A(\B<0> ), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(n5) );
  INVX1 U7 ( .A(n97), .Y(n6) );
  INVX1 U8 ( .A(n6), .Y(n7) );
  AND2X2 U9 ( .A(n105), .B(n2), .Y(n19) );
  INVX1 U10 ( .A(n80), .Y(n94) );
  INVX1 U11 ( .A(n42), .Y(n84) );
  BUFX2 U12 ( .A(n44), .Y(n8) );
  INVX1 U13 ( .A(n50), .Y(n9) );
  XOR2X1 U14 ( .A(\B<1> ), .B(n61), .Y(n10) );
  INVX1 U15 ( .A(n50), .Y(n51) );
  OR2X2 U16 ( .A(Cin), .B(n18), .Y(n35) );
  INVX1 U17 ( .A(Cin), .Y(n67) );
  AND2X2 U18 ( .A(n32), .B(n34), .Y(PG) );
  INVX1 U19 ( .A(\B<2> ), .Y(n77) );
  BUFX2 U20 ( .A(\A<3> ), .Y(n65) );
  AND2X2 U21 ( .A(n27), .B(n59), .Y(n12) );
  INVX1 U22 ( .A(n12), .Y(n13) );
  AND2X2 U23 ( .A(n8), .B(n81), .Y(n14) );
  INVX1 U24 ( .A(n14), .Y(n15) );
  INVX1 U25 ( .A(n16), .Y(GG) );
  OR2X1 U26 ( .A(n80), .B(n93), .Y(n18) );
  AND2X2 U27 ( .A(n64), .B(n52), .Y(n20) );
  INVX1 U28 ( .A(n20), .Y(n21) );
  AND2X2 U29 ( .A(n31), .B(n29), .Y(n22) );
  INVX1 U30 ( .A(n22), .Y(n23) );
  BUFX2 U31 ( .A(n83), .Y(n24) );
  BUFX2 U32 ( .A(n87), .Y(n25) );
  AND2X2 U33 ( .A(n57), .B(Cin), .Y(n26) );
  INVX1 U34 ( .A(n26), .Y(n27) );
  AND2X2 U35 ( .A(\B<3> ), .B(n62), .Y(n28) );
  INVX1 U36 ( .A(n28), .Y(n29) );
  AND2X2 U37 ( .A(n73), .B(n65), .Y(n30) );
  INVX1 U38 ( .A(n30), .Y(n31) );
  AND2X2 U39 ( .A(n48), .B(n19), .Y(n32) );
  AND2X2 U40 ( .A(n10), .B(n104), .Y(n33) );
  AND2X2 U41 ( .A(n97), .B(n33), .Y(n34) );
  INVX1 U42 ( .A(n35), .Y(n36) );
  OR2X2 U43 ( .A(n43), .B(n71), .Y(n37) );
  INVX1 U44 ( .A(n37), .Y(n38) );
  BUFX2 U45 ( .A(n88), .Y(n39) );
  AND2X2 U46 ( .A(n55), .B(n1), .Y(n40) );
  INVX1 U47 ( .A(n40), .Y(n41) );
  BUFX2 U48 ( .A(n56), .Y(n42) );
  BUFX2 U49 ( .A(n85), .Y(n43) );
  BUFX2 U50 ( .A(n86), .Y(n44) );
  BUFX2 U51 ( .A(\A<0> ), .Y(n45) );
  AND2X2 U52 ( .A(n96), .B(n7), .Y(n46) );
  INVX1 U53 ( .A(n46), .Y(n47) );
  AND2X2 U54 ( .A(n103), .B(n91), .Y(n48) );
  INVX1 U55 ( .A(n48), .Y(n49) );
  INVX1 U56 ( .A(n53), .Y(n50) );
  BUFX2 U57 ( .A(n92), .Y(n52) );
  NAND3X1 U58 ( .A(\A<2> ), .B(n72), .C(n101), .Y(n53) );
  BUFX2 U59 ( .A(n42), .Y(n54) );
  INVX1 U60 ( .A(n3), .Y(n55) );
  NAND3X1 U61 ( .A(n60), .B(n74), .C(n102), .Y(n56) );
  INVX1 U62 ( .A(n49), .Y(n57) );
  INVX1 U63 ( .A(n43), .Y(n58) );
  INVX1 U64 ( .A(n58), .Y(n59) );
  INVX1 U65 ( .A(n62), .Y(n60) );
  INVX1 U66 ( .A(n105), .Y(n82) );
  INVX1 U67 ( .A(n75), .Y(n61) );
  INVX1 U68 ( .A(n75), .Y(n76) );
  INVX1 U69 ( .A(n79), .Y(n91) );
  INVX1 U70 ( .A(n65), .Y(n62) );
  INVX1 U71 ( .A(\B<3> ), .Y(n73) );
  INVX1 U72 ( .A(n19), .Y(n63) );
  INVX1 U73 ( .A(n63), .Y(n64) );
  INVX1 U74 ( .A(n59), .Y(n93) );
  AND2X2 U75 ( .A(n23), .B(n106), .Y(n97) );
  INVX1 U76 ( .A(\A<2> ), .Y(n66) );
  INVX1 U77 ( .A(n67), .Y(n68) );
  INVX1 U78 ( .A(\B<1> ), .Y(n69) );
  INVX1 U79 ( .A(n69), .Y(n70) );
  INVX1 U80 ( .A(n33), .Y(n71) );
  INVX1 U81 ( .A(n77), .Y(n72) );
  INVX1 U82 ( .A(n73), .Y(n74) );
  INVX1 U83 ( .A(\A<1> ), .Y(n75) );
  INVX1 U84 ( .A(n67), .Y(n78) );
  NAND3X1 U85 ( .A(n61), .B(n70), .C(n100), .Y(n86) );
  OAI21X1 U86 ( .A(n8), .B(n41), .C(n9), .Y(n80) );
  NAND3X1 U87 ( .A(n5), .B(n45), .C(n99), .Y(n85) );
  XNOR2X1 U88 ( .A(\B<0> ), .B(\A<0> ), .Y(n79) );
  AOI21X1 U89 ( .A(n59), .B(n49), .C(n71), .Y(n92) );
  AOI21X1 U90 ( .A(n94), .B(n21), .C(n36), .Y(n98) );
  OAI21X1 U91 ( .A(n68), .B(n93), .C(n52), .Y(n81) );
  NAND3X1 U92 ( .A(n9), .B(n82), .C(n42), .Y(n83) );
  OAI21X1 U93 ( .A(n7), .B(n84), .C(n24), .Y(n90) );
  NAND3X1 U94 ( .A(n51), .B(n44), .C(n42), .Y(n88) );
  NAND3X1 U95 ( .A(n3), .B(n42), .C(n51), .Y(n87) );
  OAI21X1 U96 ( .A(n39), .B(n38), .C(n25), .Y(n89) );
  OAI21X1 U97 ( .A(n93), .B(n78), .C(n52), .Y(n95) );
  OAI21X1 U98 ( .A(n95), .B(n63), .C(n94), .Y(n96) );
  NAND2X1 U99 ( .A(n54), .B(n47), .Y(Cout) );
endmodule


module cla4_1 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87, n88,
         n89, n90, n91, n92, n93;

  fulladder1_7 \fa[0]  ( .A(n66), .B(\B<0> ), .Cin(n3), .S(\S<0> ), .P(n90), 
        .G(n86) );
  fulladder1_6 \fa[1]  ( .A(n22), .B(n19), .Cin(n24), .S(\S<1> ), .P(n91), .G(
        n87) );
  fulladder1_5 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n6), .S(\S<2> ), .P(n92), 
        .G(n88) );
  fulladder1_4 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n84), .S(\S<3> ), .P(n93), .G(n89) );
  INVX1 U1 ( .A(n43), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(n11), .Y(n3) );
  AND2X2 U4 ( .A(n11), .B(n55), .Y(n4) );
  INVX1 U5 ( .A(\A<2> ), .Y(n18) );
  BUFX2 U6 ( .A(n61), .Y(n5) );
  OR2X2 U7 ( .A(n36), .B(n54), .Y(n6) );
  INVX1 U8 ( .A(\A<3> ), .Y(n9) );
  INVX1 U9 ( .A(\B<0> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(n8) );
  XNOR2X1 U11 ( .A(n9), .B(\B<3> ), .Y(n15) );
  BUFX2 U12 ( .A(n91), .Y(n10) );
  INVX1 U13 ( .A(n43), .Y(n11) );
  AND2X2 U14 ( .A(n31), .B(n40), .Y(n76) );
  BUFX2 U15 ( .A(n20), .Y(n12) );
  INVX1 U16 ( .A(n21), .Y(n22) );
  BUFX2 U17 ( .A(\B<2> ), .Y(n13) );
  XOR2X1 U18 ( .A(\B<0> ), .B(n62), .Y(n14) );
  XNOR2X1 U19 ( .A(n17), .B(\A<1> ), .Y(n20) );
  BUFX2 U20 ( .A(n19), .Y(n16) );
  INVX1 U21 ( .A(\B<1> ), .Y(n17) );
  XNOR2X1 U22 ( .A(\B<2> ), .B(n18), .Y(n67) );
  BUFX4 U23 ( .A(\B<1> ), .Y(n19) );
  INVX1 U24 ( .A(\A<1> ), .Y(n21) );
  AND2X2 U25 ( .A(n65), .B(n35), .Y(n23) );
  INVX1 U26 ( .A(n23), .Y(n24) );
  OR2X2 U27 ( .A(n38), .B(n37), .Y(n25) );
  INVX1 U28 ( .A(n25), .Y(PG) );
  AND2X2 U29 ( .A(n91), .B(n20), .Y(n27) );
  AND2X2 U30 ( .A(n15), .B(n93), .Y(n28) );
  OR2X2 U31 ( .A(n74), .B(n73), .Y(n29) );
  INVX1 U32 ( .A(n29), .Y(n30) );
  BUFX2 U33 ( .A(n75), .Y(n31) );
  AND2X2 U34 ( .A(n65), .B(n44), .Y(n32) );
  INVX1 U35 ( .A(n32), .Y(n33) );
  AND2X2 U36 ( .A(n2), .B(n49), .Y(n34) );
  INVX1 U37 ( .A(n34), .Y(n35) );
  AND2X2 U38 ( .A(n43), .B(n45), .Y(n36) );
  BUFX2 U39 ( .A(n79), .Y(n37) );
  BUFX2 U40 ( .A(n78), .Y(n38) );
  BUFX2 U41 ( .A(n71), .Y(n39) );
  BUFX2 U42 ( .A(n83), .Y(n40) );
  AND2X2 U43 ( .A(n92), .B(n67), .Y(n41) );
  INVX1 U44 ( .A(n41), .Y(n42) );
  BUFX2 U45 ( .A(Cin), .Y(n43) );
  INVX1 U46 ( .A(n49), .Y(n44) );
  AND2X2 U47 ( .A(n48), .B(n33), .Y(n45) );
  INVX1 U48 ( .A(n40), .Y(n46) );
  INVX1 U49 ( .A(n46), .Y(n47) );
  BUFX2 U50 ( .A(n27), .Y(n48) );
  AND2X2 U51 ( .A(n90), .B(n14), .Y(n49) );
  AND2X2 U52 ( .A(n82), .B(n81), .Y(n50) );
  INVX1 U53 ( .A(n50), .Y(n51) );
  AND2X2 U54 ( .A(n28), .B(n51), .Y(n52) );
  INVX1 U55 ( .A(n52), .Y(n53) );
  INVX1 U56 ( .A(n70), .Y(n54) );
  AND2X2 U57 ( .A(n82), .B(n65), .Y(n55) );
  INVX1 U58 ( .A(n74), .Y(n56) );
  AND2X2 U59 ( .A(n63), .B(n45), .Y(n57) );
  INVX1 U60 ( .A(n57), .Y(n58) );
  INVX1 U61 ( .A(n73), .Y(n59) );
  INVX1 U62 ( .A(n69), .Y(n73) );
  INVX1 U63 ( .A(n42), .Y(n63) );
  AOI21X1 U64 ( .A(n82), .B(n58), .C(n4), .Y(n84) );
  OAI21X1 U65 ( .A(n74), .B(n41), .C(n28), .Y(n77) );
  INVX1 U66 ( .A(n72), .Y(n74) );
  BUFX2 U67 ( .A(\A<2> ), .Y(n60) );
  INVX1 U68 ( .A(n11), .Y(n61) );
  BUFX2 U69 ( .A(\A<0> ), .Y(n62) );
  INVX1 U70 ( .A(n68), .Y(n82) );
  INVX1 U71 ( .A(n39), .Y(n64) );
  INVX1 U72 ( .A(n64), .Y(n65) );
  INVX1 U73 ( .A(n39), .Y(n80) );
  BUFX4 U74 ( .A(\A<0> ), .Y(n66) );
  NAND3X1 U75 ( .A(n22), .B(n16), .C(n87), .Y(n69) );
  NAND3X1 U76 ( .A(n60), .B(n13), .C(n88), .Y(n72) );
  OAI21X1 U77 ( .A(n42), .B(n59), .C(n56), .Y(n68) );
  NAND3X1 U78 ( .A(n62), .B(n8), .C(n86), .Y(n71) );
  AOI21X1 U79 ( .A(n64), .B(n45), .C(n73), .Y(n70) );
  NAND3X1 U80 ( .A(\A<3> ), .B(\B<3> ), .C(n89), .Y(n83) );
  NAND3X1 U81 ( .A(n12), .B(n10), .C(n80), .Y(n75) );
  AOI22X1 U82 ( .A(n47), .B(n77), .C(n30), .D(n76), .Y(GG) );
  NAND3X1 U83 ( .A(n14), .B(n15), .C(n27), .Y(n79) );
  NAND3X1 U84 ( .A(n93), .B(n90), .C(n41), .Y(n78) );
  OAI21X1 U85 ( .A(n64), .B(n5), .C(n57), .Y(n81) );
  NAND2X1 U86 ( .A(n47), .B(n53), .Y(Cout) );
endmodule


module cla4_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80;

  fulladder1_3 \fa[0]  ( .A(\A<0> ), .B(n47), .Cin(Cin), .S(\S<0> ), .P(n77), 
        .G(n73) );
  fulladder1_2 \fa[1]  ( .A(\A<1> ), .B(n48), .Cin(n72), .S(\S<1> ), .P(n78), 
        .G(n74) );
  fulladder1_1 \fa[2]  ( .A(\A<2> ), .B(n46), .Cin(n1), .S(\S<2> ), .P(n79), 
        .G(n75) );
  fulladder1_0 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n3), .S(\S<3> ), .P(n80), 
        .G(n76) );
  AND2X2 U1 ( .A(n21), .B(n2), .Y(n1) );
  INVX8 U2 ( .A(n51), .Y(n2) );
  AND2X2 U3 ( .A(n22), .B(n4), .Y(n3) );
  INVX8 U4 ( .A(n11), .Y(n4) );
  INVX1 U5 ( .A(\A<0> ), .Y(n7) );
  INVX1 U6 ( .A(\A<2> ), .Y(n9) );
  INVX1 U7 ( .A(n44), .Y(n67) );
  BUFX2 U8 ( .A(n42), .Y(n5) );
  XNOR2X1 U9 ( .A(n7), .B(n47), .Y(n6) );
  INVX1 U10 ( .A(n40), .Y(n8) );
  XNOR2X1 U11 ( .A(n46), .B(n9), .Y(n52) );
  BUFX2 U12 ( .A(n77), .Y(n10) );
  AND2X2 U13 ( .A(n68), .B(n24), .Y(n11) );
  OR2X2 U14 ( .A(n18), .B(n37), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(PG) );
  AND2X2 U16 ( .A(n80), .B(n62), .Y(n14) );
  AND2X2 U17 ( .A(n77), .B(n6), .Y(n15) );
  INVX1 U18 ( .A(n15), .Y(n16) );
  AND2X2 U19 ( .A(n6), .B(n14), .Y(n17) );
  INVX1 U20 ( .A(n17), .Y(n18) );
  AND2X2 U21 ( .A(n68), .B(n44), .Y(n19) );
  INVX1 U22 ( .A(n19), .Y(n20) );
  OR2X2 U23 ( .A(Cin), .B(n36), .Y(n21) );
  OR2X2 U24 ( .A(Cin), .B(n20), .Y(n22) );
  AND2X2 U25 ( .A(n30), .B(n26), .Y(n23) );
  INVX1 U26 ( .A(n23), .Y(n24) );
  BUFX2 U27 ( .A(n63), .Y(n25) );
  AND2X2 U28 ( .A(n50), .B(n29), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  AND2X2 U30 ( .A(n43), .B(n16), .Y(n28) );
  INVX1 U31 ( .A(n28), .Y(n29) );
  AND2X2 U32 ( .A(n79), .B(n52), .Y(n30) );
  INVX1 U33 ( .A(n30), .Y(n31) );
  INVX1 U34 ( .A(n27), .Y(n66) );
  INVX1 U35 ( .A(n14), .Y(n32) );
  AND2X2 U36 ( .A(n14), .B(n70), .Y(n33) );
  INVX1 U37 ( .A(n33), .Y(n34) );
  AND2X2 U38 ( .A(n41), .B(n44), .Y(n35) );
  INVX1 U39 ( .A(n35), .Y(n36) );
  BUFX2 U40 ( .A(n64), .Y(n37) );
  BUFX2 U41 ( .A(n71), .Y(n38) );
  INVX1 U42 ( .A(n60), .Y(n39) );
  INVX1 U43 ( .A(n59), .Y(n60) );
  INVX1 U44 ( .A(n57), .Y(n40) );
  INVX1 U45 ( .A(n40), .Y(n41) );
  INVX1 U46 ( .A(n65), .Y(n42) );
  INVX1 U47 ( .A(n42), .Y(n43) );
  INVX1 U48 ( .A(n5), .Y(n44) );
  INVX1 U49 ( .A(n30), .Y(n45) );
  BUFX4 U50 ( .A(\B<2> ), .Y(n46) );
  BUFX4 U51 ( .A(\B<0> ), .Y(n47) );
  BUFX4 U52 ( .A(\B<1> ), .Y(n48) );
  INVX1 U53 ( .A(n56), .Y(n49) );
  INVX1 U54 ( .A(n29), .Y(n55) );
  AND2X2 U55 ( .A(n78), .B(n54), .Y(n50) );
  INVX1 U56 ( .A(n50), .Y(n58) );
  AND2X2 U57 ( .A(n41), .B(n27), .Y(n51) );
  INVX1 U58 ( .A(Cin), .Y(n56) );
  NAND3X1 U59 ( .A(\A<1> ), .B(n48), .C(n74), .Y(n57) );
  NAND3X1 U60 ( .A(\A<2> ), .B(n46), .C(n75), .Y(n59) );
  OAI21X1 U61 ( .A(n8), .B(n31), .C(n39), .Y(n53) );
  INVX2 U62 ( .A(n53), .Y(n68) );
  XOR2X1 U63 ( .A(n48), .B(\A<1> ), .Y(n54) );
  NAND3X1 U64 ( .A(\A<0> ), .B(n47), .C(n73), .Y(n65) );
  AOI21X1 U65 ( .A(n43), .B(n56), .C(n55), .Y(n72) );
  OAI21X1 U66 ( .A(n44), .B(n58), .C(n41), .Y(n61) );
  AOI21X1 U67 ( .A(n30), .B(n61), .C(n60), .Y(n63) );
  XOR2X1 U68 ( .A(\B<3> ), .B(\A<3> ), .Y(n62) );
  NAND3X1 U69 ( .A(\A<3> ), .B(\B<3> ), .C(n76), .Y(n71) );
  OAI21X1 U70 ( .A(n32), .B(n25), .C(n38), .Y(GG) );
  NAND3X1 U71 ( .A(n10), .B(n50), .C(n30), .Y(n64) );
  OAI21X1 U72 ( .A(n67), .B(n49), .C(n66), .Y(n69) );
  OAI21X1 U73 ( .A(n69), .B(n45), .C(n68), .Y(n70) );
  NAND2X1 U74 ( .A(n38), .B(n34), .Y(Cout) );
endmodule


module fulladder1_44 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(P) );
  XNOR2X1 U5 ( .A(P), .B(n2), .Y(S) );
endmodule


module fulladder1_45 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_46 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_47 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_43 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_42 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_41 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_40 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_39 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_38 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_37 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_36 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_35 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_34 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_33 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_32 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n2) );
  AND2X1 U4 ( .A(n1), .B(n2), .Y(N3) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX8 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module mux4to1_16_4 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n4, n5, n6, n8, n9, n10, n11, n13, n15, n17, n19, n21, n23,
         n25, n27, n29, n31, n33, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n76, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137;

  INVX2 U1 ( .A(n47), .Y(n48) );
  INVX1 U2 ( .A(\InD<5> ), .Y(n103) );
  INVX1 U3 ( .A(\InD<12> ), .Y(n124) );
  INVX1 U4 ( .A(\InD<2> ), .Y(n93) );
  INVX1 U5 ( .A(\InD<9> ), .Y(n115) );
  INVX1 U6 ( .A(\InD<3> ), .Y(n96) );
  INVX1 U7 ( .A(\InD<13> ), .Y(n127) );
  INVX1 U8 ( .A(\InD<6> ), .Y(n106) );
  INVX1 U9 ( .A(\InD<10> ), .Y(n118) );
  INVX1 U10 ( .A(\InD<8> ), .Y(n112) );
  INVX1 U11 ( .A(\InD<11> ), .Y(n121) );
  INVX1 U12 ( .A(\InD<14> ), .Y(n130) );
  INVX1 U13 ( .A(\InD<15> ), .Y(n134) );
  INVX1 U14 ( .A(\InD<4> ), .Y(n100) );
  INVX1 U15 ( .A(\InD<7> ), .Y(n109) );
  AND2X2 U16 ( .A(\InC<0> ), .B(n135), .Y(n1) );
  AND2X2 U17 ( .A(\InC<1> ), .B(n135), .Y(n2) );
  OR2X2 U18 ( .A(n1), .B(n4), .Y(\Out<0> ) );
  OR2X2 U19 ( .A(n5), .B(n6), .Y(n4) );
  INVX1 U20 ( .A(n89), .Y(n5) );
  INVX1 U21 ( .A(n88), .Y(n6) );
  OR2X2 U22 ( .A(n2), .B(n8), .Y(\Out<1> ) );
  OR2X2 U23 ( .A(n9), .B(n10), .Y(n8) );
  INVX1 U24 ( .A(n92), .Y(n9) );
  INVX1 U25 ( .A(n91), .Y(n10) );
  INVX4 U26 ( .A(n46), .Y(n81) );
  AND2X2 U27 ( .A(n95), .B(n94), .Y(n11) );
  INVX1 U28 ( .A(n11), .Y(\Out<2> ) );
  AND2X2 U29 ( .A(n99), .B(n98), .Y(n13) );
  INVX1 U30 ( .A(n13), .Y(\Out<3> ) );
  AND2X2 U31 ( .A(n102), .B(n101), .Y(n15) );
  INVX1 U32 ( .A(n15), .Y(\Out<4> ) );
  AND2X2 U33 ( .A(n105), .B(n104), .Y(n17) );
  INVX1 U34 ( .A(n17), .Y(\Out<5> ) );
  AND2X2 U35 ( .A(n108), .B(n107), .Y(n19) );
  INVX1 U36 ( .A(n19), .Y(\Out<6> ) );
  AND2X2 U37 ( .A(n111), .B(n110), .Y(n21) );
  INVX1 U38 ( .A(n21), .Y(\Out<7> ) );
  AND2X2 U39 ( .A(n114), .B(n113), .Y(n23) );
  INVX1 U40 ( .A(n23), .Y(\Out<8> ) );
  AND2X2 U41 ( .A(n117), .B(n116), .Y(n25) );
  INVX1 U42 ( .A(n25), .Y(\Out<9> ) );
  AND2X2 U43 ( .A(n120), .B(n119), .Y(n27) );
  INVX1 U44 ( .A(n27), .Y(\Out<10> ) );
  AND2X2 U45 ( .A(n123), .B(n122), .Y(n29) );
  INVX1 U46 ( .A(n29), .Y(\Out<11> ) );
  AND2X2 U47 ( .A(n132), .B(n131), .Y(n31) );
  INVX1 U48 ( .A(n31), .Y(\Out<14> ) );
  AND2X2 U49 ( .A(n137), .B(n136), .Y(n33) );
  INVX1 U50 ( .A(n33), .Y(\Out<15> ) );
  OR2X2 U51 ( .A(n48), .B(n106), .Y(n35) );
  INVX1 U52 ( .A(n35), .Y(n36) );
  OR2X2 U53 ( .A(n118), .B(n83), .Y(n37) );
  INVX1 U54 ( .A(n37), .Y(n38) );
  OR2X2 U55 ( .A(n48), .B(n130), .Y(n39) );
  INVX1 U56 ( .A(n39), .Y(n40) );
  AND2X2 U57 ( .A(n84), .B(\S<1> ), .Y(n41) );
  INVX1 U58 ( .A(n41), .Y(n42) );
  INVX1 U59 ( .A(n41), .Y(n43) );
  AND2X2 U60 ( .A(\S<0> ), .B(n86), .Y(n44) );
  INVX1 U61 ( .A(n44), .Y(n45) );
  INVX1 U62 ( .A(n44), .Y(n46) );
  AND2X2 U63 ( .A(\S<1> ), .B(\S<0> ), .Y(n47) );
  INVX1 U64 ( .A(n47), .Y(n49) );
  INVX2 U65 ( .A(n45), .Y(n50) );
  INVX1 U66 ( .A(n45), .Y(n51) );
  OR2X2 U67 ( .A(n48), .B(n109), .Y(n60) );
  INVX1 U68 ( .A(n87), .Y(n52) );
  INVX1 U69 ( .A(n87), .Y(n53) );
  OR2X2 U70 ( .A(n48), .B(n93), .Y(n54) );
  INVX1 U71 ( .A(n54), .Y(n55) );
  OR2X2 U72 ( .A(n83), .B(n100), .Y(n56) );
  INVX1 U73 ( .A(n56), .Y(n57) );
  OR2X2 U74 ( .A(n48), .B(n103), .Y(n58) );
  INVX1 U75 ( .A(n58), .Y(n59) );
  INVX1 U76 ( .A(n60), .Y(n61) );
  OR2X2 U77 ( .A(n83), .B(n112), .Y(n62) );
  INVX1 U78 ( .A(n62), .Y(n63) );
  OR2X2 U79 ( .A(n48), .B(n115), .Y(n64) );
  INVX1 U80 ( .A(n64), .Y(n65) );
  OR2X2 U81 ( .A(n83), .B(n121), .Y(n66) );
  INVX1 U82 ( .A(n66), .Y(n67) );
  OR2X2 U83 ( .A(n83), .B(n124), .Y(n68) );
  INVX1 U84 ( .A(n68), .Y(n69) );
  OR2X2 U85 ( .A(n82), .B(n127), .Y(n70) );
  INVX1 U86 ( .A(n70), .Y(n71) );
  OR2X2 U87 ( .A(n82), .B(n134), .Y(n72) );
  INVX1 U88 ( .A(n72), .Y(n73) );
  AND2X2 U89 ( .A(n126), .B(n125), .Y(n74) );
  INVX1 U90 ( .A(n74), .Y(\Out<12> ) );
  AND2X2 U91 ( .A(n129), .B(n128), .Y(n76) );
  INVX1 U92 ( .A(n76), .Y(\Out<13> ) );
  NAND2X1 U93 ( .A(n85), .B(\InD<0> ), .Y(n89) );
  INVX1 U94 ( .A(n87), .Y(n78) );
  INVX1 U95 ( .A(n87), .Y(n133) );
  INVX1 U96 ( .A(n87), .Y(n79) );
  INVX4 U97 ( .A(n42), .Y(n80) );
  INVX1 U98 ( .A(n43), .Y(n135) );
  BUFX2 U99 ( .A(n49), .Y(n82) );
  BUFX2 U100 ( .A(n49), .Y(n83) );
  INVX1 U101 ( .A(n83), .Y(n85) );
  INVX1 U102 ( .A(\S<0> ), .Y(n84) );
  INVX1 U103 ( .A(\S<1> ), .Y(n86) );
  INVX1 U104 ( .A(n48), .Y(n90) );
  OR2X2 U105 ( .A(\S<1> ), .B(\S<0> ), .Y(n87) );
  AOI22X1 U106 ( .A(\InB<0> ), .B(n81), .C(\InA<0> ), .D(n78), .Y(n88) );
  NAND2X1 U107 ( .A(\InD<1> ), .B(n90), .Y(n92) );
  AOI22X1 U108 ( .A(\InB<1> ), .B(n44), .C(\InA<1> ), .D(n53), .Y(n91) );
  AOI22X1 U109 ( .A(\InA<2> ), .B(n133), .C(\InB<2> ), .D(n81), .Y(n95) );
  AOI21X1 U110 ( .A(\InC<2> ), .B(n135), .C(n55), .Y(n94) );
  AOI22X1 U111 ( .A(\InA<3> ), .B(n53), .C(\InB<3> ), .D(n81), .Y(n99) );
  NOR2X1 U112 ( .A(n96), .B(n48), .Y(n97) );
  AOI21X1 U113 ( .A(n80), .B(\InC<3> ), .C(n97), .Y(n98) );
  AOI22X1 U114 ( .A(\InA<4> ), .B(n52), .C(\InB<4> ), .D(n81), .Y(n102) );
  AOI21X1 U115 ( .A(\InC<4> ), .B(n80), .C(n57), .Y(n101) );
  AOI22X1 U116 ( .A(\InA<5> ), .B(n52), .C(\InB<5> ), .D(n81), .Y(n105) );
  AOI21X1 U117 ( .A(n80), .B(\InC<5> ), .C(n59), .Y(n104) );
  AOI22X1 U118 ( .A(\InA<6> ), .B(n78), .C(\InB<6> ), .D(n50), .Y(n108) );
  AOI21X1 U119 ( .A(\InC<6> ), .B(n80), .C(n36), .Y(n107) );
  AOI22X1 U120 ( .A(\InA<7> ), .B(n53), .C(\InB<7> ), .D(n50), .Y(n111) );
  AOI21X1 U121 ( .A(\InC<7> ), .B(n80), .C(n61), .Y(n110) );
  AOI22X1 U122 ( .A(\InA<8> ), .B(n52), .C(\InB<8> ), .D(n50), .Y(n114) );
  AOI21X1 U123 ( .A(\InC<8> ), .B(n80), .C(n63), .Y(n113) );
  AOI22X1 U124 ( .A(\InA<9> ), .B(n133), .C(\InB<9> ), .D(n50), .Y(n117) );
  AOI21X1 U125 ( .A(\InC<9> ), .B(n80), .C(n65), .Y(n116) );
  AOI22X1 U126 ( .A(\InA<10> ), .B(n52), .C(\InB<10> ), .D(n50), .Y(n120) );
  AOI21X1 U127 ( .A(\InC<10> ), .B(n80), .C(n38), .Y(n119) );
  AOI22X1 U128 ( .A(\InA<11> ), .B(n78), .C(\InB<11> ), .D(n50), .Y(n123) );
  AOI21X1 U129 ( .A(\InC<11> ), .B(n135), .C(n67), .Y(n122) );
  AOI22X1 U130 ( .A(\InA<12> ), .B(n79), .C(\InB<12> ), .D(n51), .Y(n126) );
  AOI21X1 U131 ( .A(\InC<12> ), .B(n80), .C(n69), .Y(n125) );
  AOI22X1 U132 ( .A(\InA<13> ), .B(n79), .C(\InB<13> ), .D(n51), .Y(n129) );
  AOI21X1 U133 ( .A(\InC<13> ), .B(n80), .C(n71), .Y(n128) );
  AOI22X1 U134 ( .A(\InA<14> ), .B(n79), .C(\InB<14> ), .D(n50), .Y(n132) );
  AOI21X1 U135 ( .A(\InC<14> ), .B(n80), .C(n40), .Y(n131) );
  AOI22X1 U136 ( .A(\InA<15> ), .B(n133), .C(\InB<15> ), .D(n51), .Y(n137) );
  AOI21X1 U137 ( .A(\InC<15> ), .B(n80), .C(n73), .Y(n136) );
endmodule


module mux4to1_16_3 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n3, n4, n6, n7, n8, n10, n11, n12, n13, n15, n17, n19, n21,
         n23, n25, n27, n29, n31, n33, n35, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n80, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140;

  INVX1 U1 ( .A(\InD<4> ), .Y(n103) );
  INVX1 U2 ( .A(\InD<5> ), .Y(n106) );
  INVX1 U3 ( .A(\InD<12> ), .Y(n127) );
  INVX1 U4 ( .A(\InD<10> ), .Y(n122) );
  INVX1 U5 ( .A(\InD<2> ), .Y(n96) );
  INVX1 U6 ( .A(\InD<9> ), .Y(n118) );
  INVX1 U7 ( .A(\InD<3> ), .Y(n100) );
  INVX1 U8 ( .A(\InD<13> ), .Y(n130) );
  INVX1 U9 ( .A(\InD<8> ), .Y(n115) );
  INVX1 U10 ( .A(\InD<11> ), .Y(n124) );
  INVX1 U11 ( .A(\InD<15> ), .Y(n138) );
  INVX1 U12 ( .A(\InD<6> ), .Y(n109) );
  INVX1 U13 ( .A(\InD<14> ), .Y(n133) );
  INVX1 U14 ( .A(\InD<7> ), .Y(n112) );
  INVX4 U15 ( .A(n90), .Y(n137) );
  AND2X2 U16 ( .A(n82), .B(\InC<1> ), .Y(n1) );
  AND2X2 U17 ( .A(\InC<0> ), .B(n82), .Y(n2) );
  OR2X2 U18 ( .A(n45), .B(n133), .Y(n3) );
  INVX1 U19 ( .A(n3), .Y(n4) );
  OR2X2 U20 ( .A(n2), .B(n6), .Y(\Out<0> ) );
  OR2X2 U21 ( .A(n7), .B(n8), .Y(n6) );
  INVX1 U22 ( .A(n91), .Y(n7) );
  INVX1 U23 ( .A(n92), .Y(n8) );
  OR2X2 U24 ( .A(n1), .B(n10), .Y(\Out<1> ) );
  OR2X2 U25 ( .A(n11), .B(n12), .Y(n10) );
  INVX1 U26 ( .A(n94), .Y(n11) );
  INVX1 U27 ( .A(n95), .Y(n12) );
  AND2X2 U28 ( .A(n99), .B(n98), .Y(n13) );
  INVX1 U29 ( .A(n13), .Y(\Out<2> ) );
  AND2X2 U30 ( .A(n102), .B(n101), .Y(n15) );
  INVX1 U31 ( .A(n15), .Y(\Out<3> ) );
  AND2X2 U32 ( .A(n105), .B(n104), .Y(n17) );
  INVX1 U33 ( .A(n17), .Y(\Out<4> ) );
  AND2X2 U34 ( .A(n108), .B(n107), .Y(n19) );
  INVX1 U35 ( .A(n19), .Y(\Out<5> ) );
  AND2X2 U36 ( .A(n111), .B(n110), .Y(n21) );
  INVX1 U37 ( .A(n21), .Y(\Out<6> ) );
  AND2X2 U38 ( .A(n114), .B(n113), .Y(n23) );
  INVX1 U39 ( .A(n23), .Y(\Out<7> ) );
  AND2X2 U40 ( .A(n117), .B(n116), .Y(n25) );
  INVX1 U41 ( .A(n25), .Y(\Out<8> ) );
  AND2X2 U42 ( .A(n121), .B(n120), .Y(n27) );
  INVX1 U43 ( .A(n27), .Y(\Out<9> ) );
  AND2X2 U44 ( .A(n123), .B(n38), .Y(n29) );
  INVX1 U45 ( .A(n29), .Y(\Out<10> ) );
  AND2X2 U46 ( .A(n126), .B(n125), .Y(n31) );
  INVX1 U47 ( .A(n31), .Y(\Out<11> ) );
  AND2X2 U48 ( .A(n135), .B(n134), .Y(n33) );
  INVX1 U49 ( .A(n33), .Y(\Out<14> ) );
  AND2X2 U50 ( .A(n140), .B(n139), .Y(n35) );
  INVX1 U51 ( .A(n35), .Y(\Out<15> ) );
  OR2X2 U52 ( .A(n56), .B(n71), .Y(n37) );
  INVX1 U53 ( .A(n37), .Y(n38) );
  OR2X2 U54 ( .A(n85), .B(n138), .Y(n39) );
  INVX1 U55 ( .A(n39), .Y(n40) );
  AND2X2 U56 ( .A(n54), .B(n87), .Y(n41) );
  INVX1 U57 ( .A(n41), .Y(n42) );
  INVX1 U58 ( .A(n41), .Y(n43) );
  AND2X2 U59 ( .A(\S<1> ), .B(\S<0> ), .Y(n44) );
  INVX1 U60 ( .A(n44), .Y(n45) );
  INVX1 U61 ( .A(n44), .Y(n46) );
  AND2X2 U62 ( .A(n54), .B(n87), .Y(n47) );
  INVX1 U63 ( .A(n47), .Y(n48) );
  AND2X2 U64 ( .A(\S<0> ), .B(n89), .Y(n49) );
  INVX1 U65 ( .A(n49), .Y(n50) );
  INVX1 U66 ( .A(n49), .Y(n51) );
  INVX1 U67 ( .A(n51), .Y(n136) );
  BUFX2 U68 ( .A(\S<0> ), .Y(n52) );
  INVX1 U69 ( .A(n43), .Y(n53) );
  INVX1 U70 ( .A(n89), .Y(n54) );
  INVX4 U71 ( .A(n48), .Y(n55) );
  INVX1 U72 ( .A(n42), .Y(n82) );
  AND2X2 U73 ( .A(\InC<10> ), .B(n82), .Y(n56) );
  INVX1 U74 ( .A(n90), .Y(n57) );
  OR2X2 U75 ( .A(n45), .B(n100), .Y(n58) );
  INVX1 U76 ( .A(n58), .Y(n59) );
  OR2X2 U77 ( .A(n86), .B(n103), .Y(n60) );
  INVX1 U78 ( .A(n60), .Y(n61) );
  OR2X2 U79 ( .A(n45), .B(n106), .Y(n62) );
  INVX1 U80 ( .A(n62), .Y(n63) );
  OR2X2 U81 ( .A(n86), .B(n109), .Y(n64) );
  INVX1 U82 ( .A(n64), .Y(n65) );
  OR2X2 U83 ( .A(n86), .B(n112), .Y(n66) );
  INVX1 U84 ( .A(n66), .Y(n67) );
  OR2X2 U85 ( .A(n45), .B(n115), .Y(n68) );
  INVX1 U86 ( .A(n68), .Y(n69) );
  OR2X2 U87 ( .A(n85), .B(n122), .Y(n70) );
  INVX1 U88 ( .A(n70), .Y(n71) );
  OR2X2 U89 ( .A(n85), .B(n124), .Y(n72) );
  INVX1 U90 ( .A(n72), .Y(n73) );
  OR2X2 U91 ( .A(n85), .B(n127), .Y(n74) );
  INVX1 U92 ( .A(n74), .Y(n75) );
  OR2X2 U93 ( .A(n86), .B(n130), .Y(n76) );
  INVX1 U94 ( .A(n76), .Y(n77) );
  AND2X2 U95 ( .A(n129), .B(n128), .Y(n78) );
  INVX1 U96 ( .A(n78), .Y(\Out<12> ) );
  AND2X2 U97 ( .A(n132), .B(n131), .Y(n80) );
  INVX1 U98 ( .A(n80), .Y(\Out<13> ) );
  INVX4 U99 ( .A(n50), .Y(n84) );
  INVX1 U100 ( .A(n90), .Y(n83) );
  BUFX2 U101 ( .A(n46), .Y(n85) );
  BUFX2 U102 ( .A(n46), .Y(n86) );
  INVX1 U103 ( .A(n85), .Y(n88) );
  INVX1 U104 ( .A(n45), .Y(n93) );
  INVX1 U105 ( .A(\S<1> ), .Y(n89) );
  INVX1 U106 ( .A(n52), .Y(n87) );
  NAND2X1 U107 ( .A(\InD<0> ), .B(n88), .Y(n92) );
  OR2X2 U108 ( .A(\S<1> ), .B(\S<0> ), .Y(n90) );
  AOI22X1 U109 ( .A(\InB<0> ), .B(n136), .C(n137), .D(\InA<0> ), .Y(n91) );
  NAND2X1 U110 ( .A(\InD<1> ), .B(n93), .Y(n95) );
  AOI22X1 U111 ( .A(\InB<1> ), .B(n136), .C(\InA<1> ), .D(n137), .Y(n94) );
  AOI22X1 U112 ( .A(\InA<2> ), .B(n137), .C(\InB<2> ), .D(n84), .Y(n99) );
  NOR2X1 U113 ( .A(n85), .B(n96), .Y(n97) );
  AOI21X1 U114 ( .A(\InC<2> ), .B(n55), .C(n97), .Y(n98) );
  AOI22X1 U115 ( .A(\InA<3> ), .B(n137), .C(\InB<3> ), .D(n84), .Y(n102) );
  AOI21X1 U116 ( .A(\InC<3> ), .B(n55), .C(n59), .Y(n101) );
  AOI22X1 U117 ( .A(\InA<4> ), .B(n137), .C(\InB<4> ), .D(n136), .Y(n105) );
  AOI21X1 U118 ( .A(\InC<4> ), .B(n55), .C(n61), .Y(n104) );
  AOI22X1 U119 ( .A(\InA<5> ), .B(n137), .C(\InB<5> ), .D(n84), .Y(n108) );
  AOI21X1 U120 ( .A(\InC<5> ), .B(n55), .C(n63), .Y(n107) );
  AOI22X1 U121 ( .A(\InA<6> ), .B(n137), .C(\InB<6> ), .D(n84), .Y(n111) );
  AOI21X1 U122 ( .A(\InC<6> ), .B(n55), .C(n65), .Y(n110) );
  AOI22X1 U123 ( .A(\InA<7> ), .B(n137), .C(\InB<7> ), .D(n84), .Y(n114) );
  AOI21X1 U124 ( .A(\InC<7> ), .B(n55), .C(n67), .Y(n113) );
  AOI22X1 U125 ( .A(\InA<8> ), .B(n57), .C(\InB<8> ), .D(n84), .Y(n117) );
  AOI21X1 U126 ( .A(\InC<8> ), .B(n55), .C(n69), .Y(n116) );
  AOI22X1 U127 ( .A(\InA<9> ), .B(n57), .C(\InB<9> ), .D(n84), .Y(n121) );
  NOR2X1 U128 ( .A(n86), .B(n118), .Y(n119) );
  AOI21X1 U129 ( .A(\InC<9> ), .B(n55), .C(n119), .Y(n120) );
  AOI22X1 U130 ( .A(\InA<10> ), .B(n137), .C(\InB<10> ), .D(n84), .Y(n123) );
  AOI22X1 U131 ( .A(\InA<11> ), .B(n57), .C(\InB<11> ), .D(n84), .Y(n126) );
  AOI21X1 U132 ( .A(\InC<11> ), .B(n55), .C(n73), .Y(n125) );
  AOI22X1 U133 ( .A(\InA<12> ), .B(n83), .C(\InB<12> ), .D(n84), .Y(n129) );
  AOI21X1 U134 ( .A(\InC<12> ), .B(n53), .C(n75), .Y(n128) );
  AOI22X1 U135 ( .A(\InA<13> ), .B(n83), .C(\InB<13> ), .D(n84), .Y(n132) );
  AOI21X1 U136 ( .A(\InC<13> ), .B(n55), .C(n77), .Y(n131) );
  AOI22X1 U137 ( .A(\InA<14> ), .B(n83), .C(\InB<14> ), .D(n84), .Y(n135) );
  AOI21X1 U138 ( .A(\InC<14> ), .B(n53), .C(n4), .Y(n134) );
  AOI22X1 U139 ( .A(\InA<15> ), .B(n57), .C(\InB<15> ), .D(n84), .Y(n140) );
  AOI21X1 U140 ( .A(\InC<15> ), .B(n53), .C(n40), .Y(n139) );
endmodule


module mux4to1_16_2 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n33, n34, n35, n37, n38, n40, n41, n42, n44, n46, n48, n50, n52, n54,
         n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  INVX1 U1 ( .A(n22), .Y(n1) );
  AND2X2 U2 ( .A(n17), .B(n11), .Y(n2) );
  AND2X2 U3 ( .A(\InB<5> ), .B(n26), .Y(n3) );
  AND2X2 U4 ( .A(\InB<4> ), .B(n90), .Y(n4) );
  AND2X2 U5 ( .A(\InB<15> ), .B(n90), .Y(n5) );
  AND2X2 U6 ( .A(\InB<10> ), .B(n14), .Y(n6) );
  INVX1 U7 ( .A(\InA<1> ), .Y(n127) );
  INVX1 U8 ( .A(\InA<3> ), .Y(n117) );
  INVX1 U9 ( .A(\InA<2> ), .Y(n133) );
  INVX1 U10 ( .A(n94), .Y(n104) );
  AND2X2 U11 ( .A(\InB<11> ), .B(n90), .Y(n7) );
  AND2X2 U12 ( .A(\InA<15> ), .B(n16), .Y(n8) );
  INVX1 U13 ( .A(n99), .Y(n9) );
  INVX1 U14 ( .A(n99), .Y(n100) );
  INVX1 U15 ( .A(n118), .Y(n10) );
  AND2X2 U16 ( .A(\InB<1> ), .B(n1), .Y(n11) );
  INVX1 U17 ( .A(n123), .Y(n12) );
  INVX1 U18 ( .A(n113), .Y(n13) );
  INVX1 U19 ( .A(n15), .Y(n14) );
  INVX1 U20 ( .A(n25), .Y(n15) );
  INVX1 U21 ( .A(n95), .Y(n16) );
  INVX1 U22 ( .A(n118), .Y(n17) );
  AND2X2 U23 ( .A(n25), .B(\InB<0> ), .Y(n18) );
  INVX1 U24 ( .A(n18), .Y(n19) );
  AND2X2 U25 ( .A(\InB<14> ), .B(n102), .Y(n20) );
  INVX1 U26 ( .A(n20), .Y(n21) );
  INVX1 U27 ( .A(\S<0> ), .Y(n22) );
  INVX1 U28 ( .A(n22), .Y(n23) );
  INVX2 U29 ( .A(n98), .Y(n106) );
  INVX1 U30 ( .A(n113), .Y(n105) );
  INVX1 U31 ( .A(n10), .Y(n24) );
  AND2X2 U32 ( .A(n115), .B(n23), .Y(n25) );
  INVX1 U33 ( .A(n25), .Y(n28) );
  AND2X2 U34 ( .A(\InC<3> ), .B(n96), .Y(n121) );
  INVX1 U35 ( .A(\S<1> ), .Y(n115) );
  INVX1 U36 ( .A(n28), .Y(n26) );
  INVX1 U37 ( .A(n97), .Y(n27) );
  INVX2 U38 ( .A(\S<0> ), .Y(n113) );
  INVX1 U39 ( .A(n15), .Y(n90) );
  BUFX4 U40 ( .A(\S<1> ), .Y(n123) );
  OR2X2 U41 ( .A(n83), .B(n30), .Y(\Out<4> ) );
  OR2X2 U42 ( .A(n31), .B(n4), .Y(n30) );
  INVX1 U43 ( .A(n140), .Y(n31) );
  OR2X2 U44 ( .A(n85), .B(n33), .Y(\Out<6> ) );
  OR2X2 U45 ( .A(n34), .B(n35), .Y(n33) );
  INVX1 U46 ( .A(n142), .Y(n34) );
  INVX1 U47 ( .A(n143), .Y(n35) );
  OR2X2 U48 ( .A(n38), .B(n37), .Y(\Out<10> ) );
  OR2X2 U49 ( .A(n101), .B(n6), .Y(n37) );
  INVX1 U50 ( .A(n153), .Y(n38) );
  OR2X2 U51 ( .A(n7), .B(n40), .Y(\Out<11> ) );
  OR2X2 U52 ( .A(n41), .B(n107), .Y(n40) );
  INVX1 U53 ( .A(n154), .Y(n41) );
  AND2X2 U54 ( .A(n144), .B(n59), .Y(n42) );
  INVX1 U55 ( .A(n42), .Y(\Out<7> ) );
  AND2X2 U56 ( .A(n125), .B(n60), .Y(n44) );
  INVX1 U57 ( .A(n44), .Y(\Out<0> ) );
  AND2X2 U58 ( .A(n147), .B(n63), .Y(n46) );
  INVX1 U59 ( .A(n46), .Y(\Out<8> ) );
  AND2X2 U60 ( .A(n150), .B(n64), .Y(n48) );
  INVX1 U61 ( .A(n48), .Y(\Out<9> ) );
  AND2X2 U62 ( .A(n155), .B(n65), .Y(n50) );
  INVX1 U63 ( .A(n50), .Y(\Out<12> ) );
  AND2X2 U64 ( .A(n159), .B(n66), .Y(n52) );
  INVX1 U65 ( .A(n52), .Y(\Out<14> ) );
  AND2X2 U66 ( .A(n131), .B(n73), .Y(n54) );
  INVX1 U67 ( .A(n54), .Y(\Out<1> ) );
  OR2X2 U68 ( .A(n84), .B(n57), .Y(\Out<5> ) );
  OR2X2 U69 ( .A(n58), .B(n3), .Y(n57) );
  INVX1 U70 ( .A(n141), .Y(n58) );
  AND2X2 U71 ( .A(n145), .B(n146), .Y(n59) );
  AND2X2 U72 ( .A(n19), .B(n126), .Y(n60) );
  OR2X2 U73 ( .A(n8), .B(n62), .Y(\Out<15> ) );
  OR2X2 U74 ( .A(n110), .B(n5), .Y(n62) );
  AND2X2 U75 ( .A(n149), .B(n148), .Y(n63) );
  AND2X2 U76 ( .A(n152), .B(n151), .Y(n64) );
  AND2X2 U77 ( .A(n157), .B(n156), .Y(n65) );
  AND2X2 U78 ( .A(n76), .B(n21), .Y(n66) );
  AND2X2 U79 ( .A(n113), .B(n116), .Y(n67) );
  OR2X2 U80 ( .A(n113), .B(n17), .Y(n68) );
  OR2X2 U81 ( .A(n129), .B(n105), .Y(n69) );
  INVX1 U82 ( .A(n69), .Y(n70) );
  AND2X2 U83 ( .A(n137), .B(n74), .Y(n71) );
  INVX1 U84 ( .A(n71), .Y(\Out<2> ) );
  BUFX2 U85 ( .A(n132), .Y(n73) );
  BUFX2 U86 ( .A(n138), .Y(n74) );
  AND2X2 U87 ( .A(\InA<14> ), .B(n160), .Y(n75) );
  INVX1 U88 ( .A(n75), .Y(n76) );
  OR2X2 U89 ( .A(n134), .B(n123), .Y(n77) );
  INVX1 U90 ( .A(n77), .Y(n78) );
  OR2X2 U91 ( .A(n136), .B(n105), .Y(n79) );
  INVX1 U92 ( .A(n79), .Y(n80) );
  AND2X2 U93 ( .A(\InB<3> ), .B(n14), .Y(n81) );
  INVX1 U94 ( .A(n81), .Y(n82) );
  AND2X2 U95 ( .A(\InA<4> ), .B(n160), .Y(n83) );
  AND2X2 U96 ( .A(\InA<5> ), .B(n160), .Y(n84) );
  AND2X2 U97 ( .A(\InA<6> ), .B(n104), .Y(n85) );
  AND2X2 U98 ( .A(\InB<13> ), .B(n26), .Y(n86) );
  INVX1 U99 ( .A(n86), .Y(n87) );
  OR2X2 U100 ( .A(n121), .B(n120), .Y(n88) );
  INVX1 U101 ( .A(n88), .Y(n89) );
  AND2X2 U102 ( .A(n10), .B(n113), .Y(n91) );
  INVX1 U103 ( .A(n91), .Y(n92) );
  AND2X2 U104 ( .A(n113), .B(n12), .Y(n93) );
  INVX1 U105 ( .A(n93), .Y(n94) );
  INVX1 U106 ( .A(n93), .Y(n95) );
  AND2X2 U107 ( .A(n123), .B(n113), .Y(n96) );
  INVX1 U108 ( .A(n96), .Y(n97) );
  INVX1 U109 ( .A(n96), .Y(n98) );
  INVX1 U110 ( .A(n130), .Y(n99) );
  AND2X2 U111 ( .A(n16), .B(\InA<10> ), .Y(n101) );
  INVX1 U112 ( .A(n28), .Y(n102) );
  INVX1 U113 ( .A(n95), .Y(n103) );
  INVX1 U114 ( .A(n94), .Y(n160) );
  INVX1 U115 ( .A(n22), .Y(n124) );
  AND2X2 U116 ( .A(\InA<11> ), .B(n91), .Y(n107) );
  AND2X2 U117 ( .A(\InA<13> ), .B(n91), .Y(n108) );
  INVX1 U118 ( .A(n108), .Y(n109) );
  INVX1 U119 ( .A(n161), .Y(n110) );
  INVX1 U120 ( .A(n68), .Y(n111) );
  INVX1 U121 ( .A(n68), .Y(n112) );
  AND2X2 U122 ( .A(n116), .B(n13), .Y(n114) );
  INVX1 U123 ( .A(n115), .Y(n116) );
  OR2X2 U124 ( .A(n92), .B(n117), .Y(n139) );
  AND2X2 U125 ( .A(\S<0> ), .B(n123), .Y(n130) );
  INVX1 U126 ( .A(n115), .Y(n118) );
  INVX1 U127 ( .A(n118), .Y(n122) );
  AND2X2 U128 ( .A(n116), .B(n13), .Y(n119) );
  AND2X2 U129 ( .A(\InD<3> ), .B(n130), .Y(n120) );
  NAND2X1 U130 ( .A(\InA<0> ), .B(n103), .Y(n126) );
  AOI22X1 U131 ( .A(\InD<0> ), .B(n100), .C(\InC<0> ), .D(n67), .Y(n125) );
  NOR2X1 U132 ( .A(n13), .B(n127), .Y(n128) );
  AOI21X1 U133 ( .A(n128), .B(n122), .C(n2), .Y(n132) );
  NAND2X1 U134 ( .A(\InC<1> ), .B(n24), .Y(n129) );
  AOI21X1 U135 ( .A(\InD<1> ), .B(n9), .C(n70), .Y(n131) );
  NOR2X1 U136 ( .A(n105), .B(n133), .Y(n135) );
  NAND2X1 U137 ( .A(\InB<2> ), .B(n124), .Y(n134) );
  AOI21X1 U138 ( .A(n135), .B(n122), .C(n78), .Y(n138) );
  NAND2X1 U139 ( .A(\InC<2> ), .B(n116), .Y(n136) );
  AOI21X1 U140 ( .A(\InD<2> ), .B(n9), .C(n80), .Y(n137) );
  NAND3X1 U141 ( .A(n139), .B(n82), .C(n89), .Y(\Out<3> ) );
  AOI22X1 U142 ( .A(\InD<4> ), .B(n112), .C(\InC<4> ), .D(n27), .Y(n140) );
  AOI22X1 U143 ( .A(\InD<5> ), .B(n111), .C(\InC<5> ), .D(n27), .Y(n141) );
  NAND2X1 U144 ( .A(\InB<6> ), .B(n102), .Y(n143) );
  AOI22X1 U145 ( .A(\InD<6> ), .B(n119), .C(\InC<6> ), .D(n106), .Y(n142) );
  NAND2X1 U146 ( .A(\InA<7> ), .B(n104), .Y(n146) );
  NAND2X1 U147 ( .A(\InB<7> ), .B(n102), .Y(n145) );
  AOI22X1 U148 ( .A(\InD<7> ), .B(n100), .C(\InC<7> ), .D(n67), .Y(n144) );
  NAND2X1 U149 ( .A(\InA<8> ), .B(n104), .Y(n149) );
  NAND2X1 U150 ( .A(\InB<8> ), .B(n26), .Y(n148) );
  AOI22X1 U151 ( .A(\InD<8> ), .B(n119), .C(\InC<8> ), .D(n106), .Y(n147) );
  NAND2X1 U152 ( .A(\InA<9> ), .B(n91), .Y(n152) );
  NAND2X1 U153 ( .A(\InB<9> ), .B(n90), .Y(n151) );
  AOI22X1 U154 ( .A(\InD<9> ), .B(n114), .C(\InC<9> ), .D(n106), .Y(n150) );
  AOI22X1 U155 ( .A(\InD<10> ), .B(n9), .C(\InC<10> ), .D(n67), .Y(n153) );
  AOI22X1 U156 ( .A(\InD<11> ), .B(n119), .C(\InC<11> ), .D(n67), .Y(n154) );
  NAND2X1 U157 ( .A(\InA<12> ), .B(n104), .Y(n157) );
  NAND2X1 U158 ( .A(\InB<12> ), .B(n102), .Y(n156) );
  AOI22X1 U159 ( .A(\InD<12> ), .B(n119), .C(\InC<12> ), .D(n67), .Y(n155) );
  AOI22X1 U160 ( .A(\InD<13> ), .B(n114), .C(\InC<13> ), .D(n106), .Y(n158) );
  NAND3X1 U161 ( .A(n158), .B(n109), .C(n87), .Y(\Out<13> ) );
  AOI22X1 U162 ( .A(\InD<14> ), .B(n112), .C(\InC<14> ), .D(n67), .Y(n159) );
  AOI22X1 U163 ( .A(\InD<15> ), .B(n114), .C(\InC<15> ), .D(n106), .Y(n161) );
endmodule


module mux4to1_16_1 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n38, n39, n40, n42, n43, n45, n46, n48,
         n49, n50, n52, n53, n55, n56, n58, n59, n60, n63, n64, n66, n67, n69,
         n70, n72, n73, n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87,
         n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156;

  INVX1 U1 ( .A(n117), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(\S<0> ), .Y(n3) );
  NAND2X1 U4 ( .A(n4), .B(n8), .Y(n95) );
  AND2X2 U5 ( .A(n123), .B(\InB<1> ), .Y(n4) );
  INVX1 U6 ( .A(n126), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  INVX1 U8 ( .A(n5), .Y(n7) );
  INVX1 U9 ( .A(n126), .Y(n8) );
  AND2X2 U10 ( .A(\InB<14> ), .B(n120), .Y(n9) );
  AND2X2 U11 ( .A(\InA<3> ), .B(n109), .Y(n10) );
  AND2X2 U12 ( .A(\InB<8> ), .B(n31), .Y(n11) );
  INVX1 U13 ( .A(\InA<2> ), .Y(n134) );
  INVX1 U14 ( .A(n128), .Y(n118) );
  AND2X2 U15 ( .A(\InB<13> ), .B(n120), .Y(n12) );
  AND2X2 U16 ( .A(\InB<15> ), .B(n120), .Y(n13) );
  AND2X2 U17 ( .A(\InB<6> ), .B(n31), .Y(n14) );
  AND2X2 U18 ( .A(\InB<5> ), .B(n118), .Y(n15) );
  AND2X2 U19 ( .A(\InB<11> ), .B(n155), .Y(n16) );
  AND2X2 U20 ( .A(\InB<10> ), .B(n155), .Y(n17) );
  AND2X2 U21 ( .A(\InB<9> ), .B(n118), .Y(n18) );
  AND2X2 U22 ( .A(\InA<0> ), .B(n119), .Y(n19) );
  AND2X2 U23 ( .A(\InA<4> ), .B(n119), .Y(n20) );
  AND2X2 U24 ( .A(\InA<6> ), .B(n119), .Y(n21) );
  AND2X2 U25 ( .A(\InA<7> ), .B(n119), .Y(n22) );
  AND2X2 U26 ( .A(\InA<5> ), .B(n119), .Y(n23) );
  INVX1 U27 ( .A(n27), .Y(n24) );
  INVX1 U28 ( .A(n111), .Y(n25) );
  INVX1 U29 ( .A(n25), .Y(n26) );
  INVX1 U30 ( .A(n111), .Y(n27) );
  INVX1 U31 ( .A(n27), .Y(n28) );
  INVX1 U32 ( .A(n123), .Y(n29) );
  INVX1 U33 ( .A(n29), .Y(n30) );
  INVX1 U34 ( .A(n128), .Y(n31) );
  INVX1 U35 ( .A(n128), .Y(n155) );
  INVX1 U36 ( .A(n3), .Y(n32) );
  BUFX2 U37 ( .A(\S<1> ), .Y(n126) );
  AND2X2 U38 ( .A(\InB<4> ), .B(n155), .Y(n33) );
  INVX1 U39 ( .A(n113), .Y(n34) );
  INVX1 U40 ( .A(n124), .Y(n122) );
  INVX1 U41 ( .A(\S<0> ), .Y(n127) );
  OR2X2 U42 ( .A(n101), .B(n55), .Y(\Out<10> ) );
  INVX2 U43 ( .A(n110), .Y(n119) );
  AND2X2 U44 ( .A(n107), .B(\InB<3> ), .Y(n36) );
  INVX1 U45 ( .A(\S<0> ), .Y(n114) );
  AND2X2 U46 ( .A(n126), .B(n114), .Y(n35) );
  INVX1 U47 ( .A(\S<0> ), .Y(n124) );
  OR2X2 U48 ( .A(n19), .B(n38), .Y(\Out<0> ) );
  OR2X2 U49 ( .A(n39), .B(n40), .Y(n38) );
  INVX1 U50 ( .A(n129), .Y(n39) );
  INVX1 U51 ( .A(n130), .Y(n40) );
  OR2X2 U52 ( .A(n20), .B(n42), .Y(\Out<4> ) );
  OR2X2 U53 ( .A(n43), .B(n33), .Y(n42) );
  INVX1 U54 ( .A(n142), .Y(n43) );
  OR2X2 U55 ( .A(n21), .B(n45), .Y(\Out<6> ) );
  OR2X2 U56 ( .A(n46), .B(n14), .Y(n45) );
  INVX1 U57 ( .A(n144), .Y(n46) );
  OR2X2 U58 ( .A(n22), .B(n48), .Y(\Out<7> ) );
  OR2X2 U59 ( .A(n49), .B(n50), .Y(n48) );
  INVX1 U60 ( .A(n145), .Y(n49) );
  INVX1 U61 ( .A(n146), .Y(n50) );
  OR2X2 U62 ( .A(n100), .B(n52), .Y(\Out<9> ) );
  OR2X2 U63 ( .A(n53), .B(n18), .Y(n52) );
  INVX1 U64 ( .A(n148), .Y(n53) );
  OR2X2 U65 ( .A(n56), .B(n17), .Y(n55) );
  INVX1 U66 ( .A(n149), .Y(n56) );
  OR2X2 U67 ( .A(n104), .B(n58), .Y(\Out<13> ) );
  OR2X2 U68 ( .A(n59), .B(n12), .Y(n58) );
  INVX1 U69 ( .A(n153), .Y(n59) );
  AND2X2 U70 ( .A(n133), .B(n92), .Y(n60) );
  INVX1 U71 ( .A(n60), .Y(\Out<1> ) );
  OR2X2 U72 ( .A(n64), .B(n63), .Y(\Out<3> ) );
  OR2X2 U73 ( .A(n10), .B(n36), .Y(n63) );
  INVX1 U74 ( .A(n141), .Y(n64) );
  OR2X2 U75 ( .A(n23), .B(n66), .Y(\Out<5> ) );
  OR2X2 U76 ( .A(n67), .B(n15), .Y(n66) );
  INVX1 U77 ( .A(n143), .Y(n67) );
  OR2X2 U78 ( .A(n99), .B(n69), .Y(\Out<8> ) );
  OR2X2 U79 ( .A(n70), .B(n11), .Y(n69) );
  INVX1 U80 ( .A(n147), .Y(n70) );
  OR2X2 U81 ( .A(n102), .B(n72), .Y(\Out<11> ) );
  OR2X2 U82 ( .A(n73), .B(n16), .Y(n72) );
  INVX1 U83 ( .A(n150), .Y(n73) );
  OR2X2 U84 ( .A(n103), .B(n75), .Y(\Out<12> ) );
  OR2X2 U85 ( .A(n76), .B(n77), .Y(n75) );
  INVX1 U86 ( .A(n151), .Y(n76) );
  INVX1 U87 ( .A(n152), .Y(n77) );
  OR2X2 U88 ( .A(n105), .B(n79), .Y(\Out<14> ) );
  OR2X2 U89 ( .A(n80), .B(n9), .Y(n79) );
  INVX1 U90 ( .A(n154), .Y(n80) );
  OR2X2 U91 ( .A(n106), .B(n82), .Y(\Out<15> ) );
  OR2X2 U92 ( .A(n83), .B(n13), .Y(n82) );
  INVX1 U93 ( .A(n156), .Y(n83) );
  OR2X2 U94 ( .A(n132), .B(n30), .Y(n84) );
  INVX1 U95 ( .A(n84), .Y(n85) );
  OR2X2 U96 ( .A(n94), .B(n32), .Y(n86) );
  INVX1 U97 ( .A(n86), .Y(n87) );
  AND2X2 U98 ( .A(n139), .B(n90), .Y(n88) );
  INVX1 U99 ( .A(n88), .Y(\Out<2> ) );
  BUFX2 U100 ( .A(n140), .Y(n90) );
  OR2X2 U101 ( .A(n96), .B(n112), .Y(n91) );
  INVX1 U102 ( .A(n91), .Y(n92) );
  AND2X2 U103 ( .A(n115), .B(\InC<2> ), .Y(n93) );
  INVX1 U104 ( .A(n93), .Y(n94) );
  INVX1 U105 ( .A(n95), .Y(n96) );
  OR2X2 U106 ( .A(n113), .B(n135), .Y(n97) );
  INVX1 U107 ( .A(n97), .Y(n98) );
  AND2X2 U108 ( .A(\InA<8> ), .B(n119), .Y(n99) );
  AND2X2 U109 ( .A(\InA<9> ), .B(n119), .Y(n100) );
  AND2X2 U110 ( .A(\InA<10> ), .B(n119), .Y(n101) );
  AND2X2 U111 ( .A(\InA<11> ), .B(n119), .Y(n102) );
  AND2X2 U112 ( .A(\InA<12> ), .B(n119), .Y(n103) );
  AND2X2 U113 ( .A(\InA<13> ), .B(n119), .Y(n104) );
  AND2X2 U114 ( .A(\InA<14> ), .B(n119), .Y(n105) );
  AND2X2 U115 ( .A(n109), .B(\InA<15> ), .Y(n106) );
  AND2X2 U116 ( .A(n137), .B(n121), .Y(n107) );
  INVX1 U117 ( .A(n107), .Y(n108) );
  AND2X2 U118 ( .A(n137), .B(n127), .Y(n109) );
  INVX1 U119 ( .A(n109), .Y(n110) );
  AND2X2 U120 ( .A(\S<1> ), .B(\S<0> ), .Y(n111) );
  AND2X2 U121 ( .A(n131), .B(n34), .Y(n112) );
  INVX1 U122 ( .A(n137), .Y(n113) );
  INVX1 U123 ( .A(n137), .Y(n115) );
  AND2X2 U124 ( .A(n126), .B(n3), .Y(n116) );
  AND2X2 U125 ( .A(n127), .B(n115), .Y(n117) );
  INVX1 U126 ( .A(n108), .Y(n120) );
  OR2X2 U127 ( .A(\S<1> ), .B(n124), .Y(n128) );
  INVX1 U128 ( .A(\S<1> ), .Y(n137) );
  INVX1 U129 ( .A(n3), .Y(n121) );
  INVX1 U130 ( .A(n127), .Y(n123) );
  AND2X2 U131 ( .A(n114), .B(\InA<1> ), .Y(n131) );
  AND2X2 U132 ( .A(n115), .B(n122), .Y(n125) );
  NAND2X1 U133 ( .A(\InB<0> ), .B(n31), .Y(n130) );
  AOI22X1 U134 ( .A(\InD<0> ), .B(n111), .C(\InC<0> ), .D(n116), .Y(n129) );
  NAND2X1 U135 ( .A(\InC<1> ), .B(n6), .Y(n132) );
  AOI21X1 U136 ( .A(\InD<1> ), .B(n26), .C(n85), .Y(n133) );
  NOR2X1 U137 ( .A(n32), .B(n134), .Y(n136) );
  NAND2X1 U138 ( .A(\InB<2> ), .B(n122), .Y(n135) );
  AOI21X1 U139 ( .A(n8), .B(n136), .C(n98), .Y(n140) );
  AND2X2 U140 ( .A(n7), .B(n32), .Y(n138) );
  AOI21X1 U141 ( .A(\InD<2> ), .B(n138), .C(n87), .Y(n139) );
  AOI22X1 U142 ( .A(\InD<3> ), .B(n28), .C(\InC<3> ), .D(n117), .Y(n141) );
  AOI22X1 U143 ( .A(\InD<4> ), .B(n26), .C(\InC<4> ), .D(n117), .Y(n142) );
  AOI22X1 U144 ( .A(\InD<5> ), .B(n111), .C(\InC<5> ), .D(n117), .Y(n143) );
  AOI22X1 U145 ( .A(\InD<6> ), .B(n24), .C(\InC<6> ), .D(n117), .Y(n144) );
  NAND2X1 U146 ( .A(\InB<7> ), .B(n118), .Y(n146) );
  AOI22X1 U147 ( .A(\InD<7> ), .B(n111), .C(n116), .D(\InC<7> ), .Y(n145) );
  AOI22X1 U148 ( .A(\InD<8> ), .B(n111), .C(\InC<8> ), .D(n35), .Y(n147) );
  AOI22X1 U149 ( .A(\InD<9> ), .B(n125), .C(\InC<9> ), .D(n116), .Y(n148) );
  AOI22X1 U150 ( .A(\InD<10> ), .B(n111), .C(\InC<10> ), .D(n35), .Y(n149) );
  AOI22X1 U151 ( .A(\InD<11> ), .B(n138), .C(\InC<11> ), .D(n35), .Y(n150) );
  NAND2X1 U152 ( .A(\InB<12> ), .B(n120), .Y(n152) );
  AOI22X1 U153 ( .A(\InD<12> ), .B(n111), .C(\InC<12> ), .D(n117), .Y(n151) );
  AOI22X1 U154 ( .A(\InD<13> ), .B(n138), .C(\InC<13> ), .D(n2), .Y(n153) );
  AOI22X1 U155 ( .A(\InD<14> ), .B(n111), .C(\InC<14> ), .D(n35), .Y(n154) );
  AOI22X1 U156 ( .A(\InD<15> ), .B(n138), .C(\InC<15> ), .D(n35), .Y(n156) );
endmodule


module demux1to8_0 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n3, n4, n5, n6, n7, n8, n10, n12, n14, n16, n18, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41;

  AND2X1 U1 ( .A(n7), .B(n40), .Y(Out1) );
  INVX1 U2 ( .A(\S<2> ), .Y(n38) );
  AND2X2 U3 ( .A(n5), .B(n23), .Y(Out5) );
  INVX1 U4 ( .A(In), .Y(n3) );
  INVX1 U5 ( .A(In), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(n5) );
  INVX1 U7 ( .A(n4), .Y(n6) );
  INVX1 U8 ( .A(n3), .Y(n7) );
  OR2X2 U9 ( .A(n32), .B(n20), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(Out7) );
  OR2X2 U11 ( .A(n3), .B(n33), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(Out4) );
  OR2X2 U13 ( .A(n3), .B(n24), .Y(n12) );
  INVX1 U14 ( .A(n12), .Y(Out3) );
  OR2X2 U15 ( .A(n34), .B(n35), .Y(n14) );
  INVX1 U16 ( .A(n14), .Y(Out0) );
  OR2X2 U17 ( .A(n36), .B(n25), .Y(n16) );
  INVX1 U18 ( .A(n16), .Y(Out2) );
  OR2X2 U19 ( .A(n36), .B(n21), .Y(n18) );
  INVX1 U20 ( .A(n18), .Y(Out6) );
  OR2X1 U21 ( .A(n29), .B(n37), .Y(n20) );
  OR2X1 U22 ( .A(n29), .B(\S<0> ), .Y(n21) );
  OR2X1 U23 ( .A(n27), .B(\S<1> ), .Y(n22) );
  INVX1 U24 ( .A(n22), .Y(n23) );
  OR2X1 U25 ( .A(n31), .B(n37), .Y(n24) );
  INVX1 U26 ( .A(\S<0> ), .Y(n37) );
  OR2X1 U27 ( .A(n31), .B(\S<0> ), .Y(n25) );
  AND2X1 U28 ( .A(\S<0> ), .B(\S<2> ), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  AND2X1 U30 ( .A(\S<2> ), .B(\S<1> ), .Y(n28) );
  INVX1 U31 ( .A(n28), .Y(n29) );
  AND2X1 U32 ( .A(n38), .B(\S<1> ), .Y(n30) );
  INVX1 U33 ( .A(n30), .Y(n31) );
  INVX1 U34 ( .A(n5), .Y(n32) );
  INVX1 U35 ( .A(n39), .Y(n33) );
  INVX1 U36 ( .A(n6), .Y(n34) );
  INVX1 U37 ( .A(n41), .Y(n35) );
  INVX1 U38 ( .A(n6), .Y(n36) );
  NOR3X1 U39 ( .A(\S<1> ), .B(n38), .C(\S<0> ), .Y(n39) );
  NOR3X1 U40 ( .A(\S<1> ), .B(\S<2> ), .C(n37), .Y(n40) );
  NOR3X1 U41 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n41) );
endmodule


module demux1to8_1 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;

  AND2X1 U1 ( .A(n2), .B(n25), .Y(Out4) );
  AND2X1 U2 ( .A(n22), .B(n26), .Y(Out1) );
  AND2X1 U3 ( .A(In), .B(n27), .Y(Out0) );
  INVX1 U4 ( .A(\S<0> ), .Y(n23) );
  INVX1 U5 ( .A(\S<2> ), .Y(n24) );
  INVX1 U6 ( .A(n3), .Y(n2) );
  INVX1 U7 ( .A(In), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(n4) );
  OR2X2 U9 ( .A(n3), .B(n7), .Y(n5) );
  INVX1 U10 ( .A(n5), .Y(Out2) );
  OR2X1 U11 ( .A(n21), .B(\S<0> ), .Y(n7) );
  OR2X1 U12 ( .A(n19), .B(n23), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  OR2X1 U14 ( .A(n19), .B(\S<0> ), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  OR2X1 U16 ( .A(n17), .B(\S<1> ), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  OR2X1 U18 ( .A(n21), .B(n23), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  AND2X1 U20 ( .A(\S<0> ), .B(\S<2> ), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  AND2X1 U22 ( .A(\S<2> ), .B(\S<1> ), .Y(n18) );
  INVX1 U23 ( .A(n18), .Y(n19) );
  AND2X1 U24 ( .A(n24), .B(\S<1> ), .Y(n20) );
  INVX1 U25 ( .A(n20), .Y(n21) );
  INVX1 U26 ( .A(n3), .Y(n22) );
  AND2X2 U27 ( .A(n4), .B(n9), .Y(Out7) );
  AND2X2 U28 ( .A(n2), .B(n11), .Y(Out6) );
  AND2X2 U29 ( .A(n4), .B(n13), .Y(Out5) );
  NOR3X1 U30 ( .A(\S<1> ), .B(n24), .C(\S<0> ), .Y(n25) );
  AND2X2 U31 ( .A(n22), .B(n15), .Y(Out3) );
  NOR3X1 U32 ( .A(\S<1> ), .B(\S<2> ), .C(n23), .Y(n26) );
  NOR3X1 U33 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n27) );
endmodule


module demux1to8_2 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n3, n5, n7, n9, n11, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39;

  INVX1 U1 ( .A(\S<2> ), .Y(n36) );
  OR2X2 U2 ( .A(n29), .B(n18), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out6) );
  OR2X2 U4 ( .A(n31), .B(n21), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out2) );
  OR2X2 U6 ( .A(n34), .B(n28), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out0) );
  OR2X2 U8 ( .A(n29), .B(n30), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out4) );
  OR2X2 U10 ( .A(n31), .B(n32), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out1) );
  OR2X2 U12 ( .A(n33), .B(n17), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(Out7) );
  OR2X2 U14 ( .A(n33), .B(n19), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(Out5) );
  OR2X2 U16 ( .A(n34), .B(n20), .Y(n15) );
  INVX1 U17 ( .A(n15), .Y(Out3) );
  OR2X1 U18 ( .A(n25), .B(n35), .Y(n17) );
  OR2X1 U19 ( .A(n25), .B(\S<0> ), .Y(n18) );
  OR2X1 U20 ( .A(n23), .B(\S<1> ), .Y(n19) );
  OR2X1 U21 ( .A(n27), .B(n35), .Y(n20) );
  INVX1 U22 ( .A(\S<0> ), .Y(n35) );
  OR2X1 U23 ( .A(n27), .B(\S<0> ), .Y(n21) );
  AND2X1 U24 ( .A(\S<0> ), .B(\S<2> ), .Y(n22) );
  INVX1 U25 ( .A(n22), .Y(n23) );
  AND2X1 U26 ( .A(\S<2> ), .B(\S<1> ), .Y(n24) );
  INVX1 U27 ( .A(n24), .Y(n25) );
  AND2X1 U28 ( .A(n36), .B(\S<1> ), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  INVX1 U30 ( .A(n39), .Y(n28) );
  INVX1 U31 ( .A(In), .Y(n29) );
  INVX1 U32 ( .A(n37), .Y(n30) );
  INVX1 U33 ( .A(In), .Y(n31) );
  INVX1 U34 ( .A(n38), .Y(n32) );
  INVX1 U35 ( .A(In), .Y(n33) );
  INVX1 U36 ( .A(In), .Y(n34) );
  NOR3X1 U37 ( .A(\S<1> ), .B(n36), .C(\S<0> ), .Y(n37) );
  NOR3X1 U38 ( .A(\S<1> ), .B(\S<2> ), .C(n35), .Y(n38) );
  NOR3X1 U39 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n39) );
endmodule


module demux1to8_3 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n3, n5, n7, n9, n11, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43;

  INVX1 U1 ( .A(\S<2> ), .Y(n40) );
  OR2X2 U2 ( .A(n28), .B(n18), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out6) );
  OR2X2 U4 ( .A(n29), .B(n21), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out2) );
  OR2X2 U6 ( .A(n30), .B(n31), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out0) );
  OR2X2 U8 ( .A(n32), .B(n33), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out4) );
  OR2X2 U10 ( .A(n34), .B(n35), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out1) );
  OR2X2 U12 ( .A(n36), .B(n17), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(Out7) );
  OR2X2 U14 ( .A(n37), .B(n19), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(Out5) );
  OR2X2 U16 ( .A(n38), .B(n20), .Y(n15) );
  INVX1 U17 ( .A(n15), .Y(Out3) );
  OR2X1 U18 ( .A(n25), .B(n39), .Y(n17) );
  OR2X1 U19 ( .A(n25), .B(\S<0> ), .Y(n18) );
  OR2X1 U20 ( .A(n23), .B(\S<1> ), .Y(n19) );
  OR2X1 U21 ( .A(n27), .B(n39), .Y(n20) );
  INVX1 U22 ( .A(\S<0> ), .Y(n39) );
  OR2X1 U23 ( .A(n27), .B(\S<0> ), .Y(n21) );
  AND2X1 U24 ( .A(\S<0> ), .B(\S<2> ), .Y(n22) );
  INVX1 U25 ( .A(n22), .Y(n23) );
  AND2X1 U26 ( .A(\S<2> ), .B(\S<1> ), .Y(n24) );
  INVX1 U27 ( .A(n24), .Y(n25) );
  AND2X1 U28 ( .A(n40), .B(\S<1> ), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  INVX1 U30 ( .A(In), .Y(n28) );
  INVX1 U31 ( .A(In), .Y(n29) );
  INVX1 U32 ( .A(In), .Y(n30) );
  INVX1 U33 ( .A(n43), .Y(n31) );
  INVX1 U34 ( .A(In), .Y(n32) );
  INVX1 U35 ( .A(n41), .Y(n33) );
  INVX1 U36 ( .A(In), .Y(n34) );
  INVX1 U37 ( .A(n42), .Y(n35) );
  INVX1 U38 ( .A(In), .Y(n36) );
  INVX1 U39 ( .A(In), .Y(n37) );
  INVX1 U40 ( .A(In), .Y(n38) );
  NOR3X1 U41 ( .A(\S<1> ), .B(n40), .C(\S<0> ), .Y(n41) );
  NOR3X1 U42 ( .A(\S<1> ), .B(\S<2> ), .C(n39), .Y(n42) );
  NOR3X1 U43 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n43) );
endmodule


module demux1to8_4 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;

  AND2X1 U1 ( .A(n1), .B(n21), .Y(Out4) );
  AND2X1 U2 ( .A(n1), .B(n23), .Y(Out0) );
  INVX1 U3 ( .A(\S<2> ), .Y(n20) );
  INVX1 U4 ( .A(\S<0> ), .Y(n19) );
  INVX1 U5 ( .A(n18), .Y(n1) );
  OR2X1 U6 ( .A(n15), .B(n19), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  OR2X1 U8 ( .A(n15), .B(\S<0> ), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(n5) );
  OR2X1 U10 ( .A(n13), .B(\S<1> ), .Y(n6) );
  INVX1 U11 ( .A(n6), .Y(n7) );
  OR2X1 U12 ( .A(n17), .B(n19), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  OR2X1 U14 ( .A(n17), .B(\S<0> ), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  AND2X1 U16 ( .A(\S<0> ), .B(\S<2> ), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  AND2X1 U18 ( .A(\S<2> ), .B(\S<1> ), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  AND2X1 U20 ( .A(n20), .B(\S<1> ), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  INVX1 U22 ( .A(In), .Y(n18) );
  AND2X2 U23 ( .A(In), .B(n3), .Y(Out7) );
  AND2X2 U24 ( .A(In), .B(n5), .Y(Out6) );
  AND2X2 U25 ( .A(n1), .B(n7), .Y(Out5) );
  NOR3X1 U26 ( .A(\S<1> ), .B(n20), .C(\S<0> ), .Y(n21) );
  AND2X2 U27 ( .A(In), .B(n9), .Y(Out3) );
  AND2X2 U28 ( .A(In), .B(n11), .Y(Out2) );
  NOR3X1 U29 ( .A(\S<1> ), .B(\S<2> ), .C(n19), .Y(n22) );
  AND2X2 U30 ( .A(In), .B(n22), .Y(Out1) );
  NOR3X1 U31 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n23) );
endmodule


module demux1to8_5 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  INVX1 U1 ( .A(n20), .Y(n1) );
  AND2X1 U2 ( .A(n21), .B(n26), .Y(Out0) );
  AND2X1 U3 ( .A(n19), .B(n25), .Y(Out1) );
  INVX1 U4 ( .A(\S<0> ), .Y(n22) );
  INVX1 U5 ( .A(\S<2> ), .Y(n23) );
  OR2X1 U6 ( .A(n15), .B(n22), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  OR2X1 U8 ( .A(n15), .B(\S<0> ), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(n5) );
  OR2X1 U10 ( .A(n13), .B(\S<1> ), .Y(n6) );
  INVX1 U11 ( .A(n6), .Y(n7) );
  OR2X1 U12 ( .A(n17), .B(n22), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  OR2X1 U14 ( .A(n17), .B(\S<0> ), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  AND2X1 U16 ( .A(\S<0> ), .B(\S<2> ), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  AND2X1 U18 ( .A(\S<2> ), .B(\S<1> ), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  AND2X1 U20 ( .A(n23), .B(\S<1> ), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  INVX1 U22 ( .A(In), .Y(n18) );
  INVX1 U23 ( .A(n18), .Y(n19) );
  INVX1 U24 ( .A(In), .Y(n20) );
  INVX1 U25 ( .A(n20), .Y(n21) );
  AND2X2 U26 ( .A(n1), .B(n3), .Y(Out7) );
  AND2X2 U27 ( .A(n21), .B(n5), .Y(Out6) );
  AND2X2 U28 ( .A(n1), .B(n7), .Y(Out5) );
  NOR3X1 U29 ( .A(\S<1> ), .B(n23), .C(\S<0> ), .Y(n24) );
  AND2X2 U30 ( .A(In), .B(n24), .Y(Out4) );
  AND2X2 U31 ( .A(n1), .B(n9), .Y(Out3) );
  AND2X2 U32 ( .A(n19), .B(n11), .Y(Out2) );
  NOR3X1 U33 ( .A(\S<1> ), .B(\S<2> ), .C(n22), .Y(n25) );
  NOR3X1 U34 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n26) );
endmodule


module demux1to8_6 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;

  INVX1 U1 ( .A(\S<2> ), .Y(n24) );
  INVX1 U2 ( .A(\S<0> ), .Y(n23) );
  AND2X1 U3 ( .A(n2), .B(n26), .Y(Out1) );
  INVX1 U4 ( .A(n5), .Y(n2) );
  OR2X2 U5 ( .A(n22), .B(n10), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(Out5) );
  INVX1 U7 ( .A(In), .Y(n5) );
  OR2X1 U8 ( .A(n18), .B(n23), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(n7) );
  OR2X1 U10 ( .A(n18), .B(\S<0> ), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  OR2X1 U12 ( .A(n16), .B(\S<1> ), .Y(n10) );
  OR2X1 U13 ( .A(n20), .B(n23), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(n12) );
  OR2X1 U15 ( .A(n20), .B(\S<0> ), .Y(n13) );
  INVX1 U16 ( .A(n13), .Y(n14) );
  AND2X1 U17 ( .A(\S<0> ), .B(\S<2> ), .Y(n15) );
  INVX1 U18 ( .A(n15), .Y(n16) );
  AND2X1 U19 ( .A(\S<2> ), .B(\S<1> ), .Y(n17) );
  INVX1 U20 ( .A(n17), .Y(n18) );
  AND2X1 U21 ( .A(n24), .B(\S<1> ), .Y(n19) );
  INVX1 U22 ( .A(n19), .Y(n20) );
  INVX1 U23 ( .A(n22), .Y(n21) );
  INVX1 U24 ( .A(In), .Y(n22) );
  AND2X2 U25 ( .A(n21), .B(n7), .Y(Out7) );
  AND2X2 U26 ( .A(n21), .B(n9), .Y(Out6) );
  NOR3X1 U27 ( .A(\S<1> ), .B(n24), .C(\S<0> ), .Y(n25) );
  AND2X2 U28 ( .A(n21), .B(n25), .Y(Out4) );
  AND2X2 U29 ( .A(n2), .B(n12), .Y(Out3) );
  AND2X2 U30 ( .A(n2), .B(n14), .Y(Out2) );
  NOR3X1 U31 ( .A(\S<1> ), .B(\S<2> ), .C(n23), .Y(n26) );
  NOR3X1 U32 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n27) );
  AND2X2 U33 ( .A(n21), .B(n27), .Y(Out0) );
endmodule


module demux1to8_7 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  AND2X1 U1 ( .A(n3), .B(n24), .Y(Out4) );
  AND2X1 U2 ( .A(n3), .B(n26), .Y(Out0) );
  INVX1 U3 ( .A(\S<2> ), .Y(n23) );
  INVX1 U4 ( .A(\S<0> ), .Y(n22) );
  INVX1 U5 ( .A(In), .Y(n1) );
  INVX1 U6 ( .A(In), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  INVX1 U8 ( .A(n2), .Y(n4) );
  INVX1 U9 ( .A(n1), .Y(n5) );
  OR2X1 U10 ( .A(n19), .B(n22), .Y(n6) );
  INVX1 U11 ( .A(n6), .Y(n7) );
  OR2X1 U12 ( .A(n19), .B(\S<0> ), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  OR2X1 U14 ( .A(n17), .B(\S<1> ), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  OR2X1 U16 ( .A(n21), .B(n22), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  OR2X1 U18 ( .A(n21), .B(\S<0> ), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  AND2X1 U20 ( .A(\S<0> ), .B(\S<2> ), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  AND2X1 U22 ( .A(\S<2> ), .B(\S<1> ), .Y(n18) );
  INVX1 U23 ( .A(n18), .Y(n19) );
  AND2X1 U24 ( .A(n23), .B(\S<1> ), .Y(n20) );
  INVX1 U25 ( .A(n20), .Y(n21) );
  AND2X2 U26 ( .A(n5), .B(n7), .Y(Out7) );
  AND2X2 U27 ( .A(n5), .B(n9), .Y(Out6) );
  AND2X2 U28 ( .A(n4), .B(n11), .Y(Out5) );
  NOR3X1 U29 ( .A(\S<1> ), .B(n23), .C(\S<0> ), .Y(n24) );
  AND2X2 U30 ( .A(n4), .B(n13), .Y(Out3) );
  AND2X2 U31 ( .A(n4), .B(n15), .Y(Out2) );
  NOR3X1 U32 ( .A(\S<1> ), .B(\S<2> ), .C(n22), .Y(n25) );
  AND2X2 U33 ( .A(n5), .B(n25), .Y(Out1) );
  NOR3X1 U34 ( .A(\S<1> ), .B(\S<2> ), .C(\S<0> ), .Y(n26) );
endmodule


module demux1to8_8 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n2, n3, n4, n5, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20;

  AND2X1 U1 ( .A(n17), .B(n2), .Y(Out2) );
  INVX8 U2 ( .A(\S<0> ), .Y(n2) );
  OR2X1 U3 ( .A(\S<2> ), .B(n13), .Y(n3) );
  OR2X1 U4 ( .A(n4), .B(\S<0> ), .Y(n7) );
  INVX1 U5 ( .A(\S<0> ), .Y(n18) );
  OR2X2 U6 ( .A(n16), .B(n11), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n18), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out7) );
  INVX1 U9 ( .A(n7), .Y(Out6) );
  OR2X2 U10 ( .A(n20), .B(n18), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out3) );
  OR2X2 U12 ( .A(n15), .B(n14), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  NOR3X1 U14 ( .A(n16), .B(n13), .C(\S<2> ), .Y(n17) );
  INVX1 U15 ( .A(In), .Y(n13) );
  INVX1 U16 ( .A(\S<2> ), .Y(n14) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(\S<1> ), .Y(n16) );
  INVX1 U19 ( .A(n17), .Y(n20) );
  INVX1 U20 ( .A(n12), .Y(n19) );
  NOR3X1 U21 ( .A(\S<1> ), .B(n19), .C(n18), .Y(Out5) );
  NOR3X1 U22 ( .A(\S<1> ), .B(n19), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U23 ( .A(\S<1> ), .B(n3), .C(n18), .Y(Out1) );
  NOR3X1 U24 ( .A(\S<1> ), .B(n3), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_9 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n7, n9, n11, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22;

  INVX1 U1 ( .A(n14), .Y(n1) );
  OR2X1 U2 ( .A(n2), .B(\S<0> ), .Y(n11) );
  OR2X1 U3 ( .A(n15), .B(\S<2> ), .Y(n3) );
  OR2X1 U4 ( .A(n4), .B(\S<0> ), .Y(n7) );
  INVX1 U5 ( .A(\S<0> ), .Y(n20) );
  INVX1 U6 ( .A(n19), .Y(n2) );
  OR2X2 U7 ( .A(n18), .B(n13), .Y(n4) );
  OR2X2 U8 ( .A(n4), .B(n20), .Y(n5) );
  INVX1 U9 ( .A(n5), .Y(Out7) );
  INVX1 U10 ( .A(n7), .Y(Out6) );
  OR2X2 U11 ( .A(n22), .B(n20), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Out3) );
  INVX1 U13 ( .A(n11), .Y(Out2) );
  OR2X2 U14 ( .A(n17), .B(n16), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(n14) );
  NOR3X1 U16 ( .A(n18), .B(\S<2> ), .C(n15), .Y(n19) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(\S<2> ), .Y(n16) );
  INVX1 U19 ( .A(In), .Y(n17) );
  INVX1 U20 ( .A(\S<1> ), .Y(n18) );
  INVX1 U21 ( .A(n19), .Y(n22) );
  INVX1 U22 ( .A(n14), .Y(n21) );
  NOR3X1 U23 ( .A(\S<1> ), .B(n21), .C(n20), .Y(Out5) );
  NOR3X1 U24 ( .A(\S<1> ), .B(n1), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U25 ( .A(\S<1> ), .B(n3), .C(n20), .Y(Out1) );
  NOR3X1 U26 ( .A(\S<1> ), .B(n3), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_10 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n2, n3, n4, n5, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20;

  AND2X1 U1 ( .A(n17), .B(n2), .Y(Out2) );
  INVX8 U2 ( .A(\S<0> ), .Y(n2) );
  OR2X1 U3 ( .A(n13), .B(\S<2> ), .Y(n3) );
  OR2X1 U4 ( .A(n4), .B(\S<0> ), .Y(n7) );
  INVX1 U5 ( .A(\S<0> ), .Y(n18) );
  OR2X2 U6 ( .A(n16), .B(n11), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n18), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out7) );
  INVX1 U9 ( .A(n7), .Y(Out6) );
  OR2X2 U10 ( .A(n20), .B(n18), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out3) );
  OR2X2 U12 ( .A(n15), .B(n14), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  NOR3X1 U14 ( .A(n16), .B(\S<2> ), .C(n13), .Y(n17) );
  INVX1 U15 ( .A(In), .Y(n13) );
  INVX1 U16 ( .A(\S<2> ), .Y(n14) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(\S<1> ), .Y(n16) );
  INVX1 U19 ( .A(n17), .Y(n20) );
  INVX1 U20 ( .A(n12), .Y(n19) );
  NOR3X1 U21 ( .A(\S<1> ), .B(n19), .C(n18), .Y(Out5) );
  NOR3X1 U22 ( .A(\S<1> ), .B(n19), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U23 ( .A(\S<1> ), .B(n3), .C(n18), .Y(Out1) );
  NOR3X1 U24 ( .A(\S<1> ), .B(n3), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_11 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n4, n5, n6, n7, n9, n11, n13, n14, n15, n16, n17, n18;

  AND2X1 U1 ( .A(n2), .B(\S<0> ), .Y(Out3) );
  OR2X1 U2 ( .A(n5), .B(\S<0> ), .Y(n11) );
  OR2X1 U3 ( .A(n14), .B(\S<2> ), .Y(n4) );
  OR2X1 U4 ( .A(n6), .B(\S<0> ), .Y(n9) );
  INVX1 U5 ( .A(\S<2> ), .Y(n18) );
  AND2X1 U6 ( .A(n18), .B(\S<1> ), .Y(n1) );
  AND2X2 U7 ( .A(In), .B(n1), .Y(n2) );
  INVX1 U8 ( .A(n2), .Y(n5) );
  INVX1 U9 ( .A(\S<0> ), .Y(n17) );
  OR2X2 U10 ( .A(n16), .B(n13), .Y(n6) );
  OR2X2 U11 ( .A(n6), .B(n17), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(Out7) );
  INVX1 U13 ( .A(n9), .Y(Out6) );
  INVX1 U14 ( .A(n11), .Y(Out2) );
  OR2X2 U15 ( .A(n15), .B(n18), .Y(n13) );
  INVX1 U16 ( .A(In), .Y(n14) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(\S<1> ), .Y(n16) );
  NOR3X1 U19 ( .A(\S<1> ), .B(n13), .C(n17), .Y(Out5) );
  NOR3X1 U20 ( .A(\S<1> ), .B(n13), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U21 ( .A(\S<1> ), .B(n4), .C(n17), .Y(Out1) );
  NOR3X1 U22 ( .A(\S<1> ), .B(n4), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_12 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n4, n5, n6, n7, n9, n11, n13, n14, n15, n16, n17, n18, n19,
         n20;

  AND2X1 U1 ( .A(n2), .B(n18), .Y(Out2) );
  OR2X1 U2 ( .A(n15), .B(\S<2> ), .Y(n4) );
  OR2X1 U3 ( .A(n6), .B(\S<0> ), .Y(n9) );
  INVX1 U4 ( .A(\S<0> ), .Y(n18) );
  INVX1 U5 ( .A(\S<2> ), .Y(n19) );
  AND2X1 U6 ( .A(n19), .B(\S<1> ), .Y(n1) );
  AND2X2 U7 ( .A(In), .B(n1), .Y(n2) );
  INVX1 U8 ( .A(n2), .Y(n5) );
  OR2X2 U9 ( .A(n17), .B(n13), .Y(n6) );
  OR2X2 U10 ( .A(n6), .B(n18), .Y(n7) );
  INVX1 U11 ( .A(n7), .Y(Out7) );
  INVX1 U12 ( .A(n9), .Y(Out6) );
  OR2X2 U13 ( .A(n5), .B(n18), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(Out3) );
  OR2X2 U15 ( .A(n16), .B(n19), .Y(n13) );
  INVX1 U16 ( .A(n13), .Y(n14) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(In), .Y(n16) );
  INVX1 U19 ( .A(\S<1> ), .Y(n17) );
  INVX1 U20 ( .A(n14), .Y(n20) );
  NOR3X1 U21 ( .A(\S<1> ), .B(n20), .C(n18), .Y(Out5) );
  NOR3X1 U22 ( .A(\S<1> ), .B(n20), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U23 ( .A(\S<1> ), .B(n4), .C(n18), .Y(Out1) );
  NOR3X1 U24 ( .A(\S<1> ), .B(n4), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_13 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n3, n4, n5, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22;

  INVX1 U1 ( .A(n15), .Y(n1) );
  AND2X2 U2 ( .A(n11), .B(n21), .Y(Out2) );
  AND2X2 U3 ( .A(n1), .B(\S<2> ), .Y(n20) );
  AND2X2 U4 ( .A(\S<1> ), .B(n14), .Y(n11) );
  OR2X1 U5 ( .A(n4), .B(\S<0> ), .Y(n7) );
  OR2X1 U6 ( .A(n19), .B(\S<2> ), .Y(n13) );
  INVX1 U7 ( .A(\S<0> ), .Y(n21) );
  OR2X2 U8 ( .A(n15), .B(n16), .Y(n3) );
  OR2X2 U9 ( .A(n18), .B(n17), .Y(n4) );
  OR2X2 U10 ( .A(n4), .B(n21), .Y(n5) );
  INVX1 U11 ( .A(n5), .Y(Out7) );
  INVX1 U12 ( .A(n7), .Y(Out6) );
  OR2X2 U13 ( .A(n12), .B(n21), .Y(n9) );
  INVX1 U14 ( .A(n9), .Y(Out3) );
  INVX1 U15 ( .A(n11), .Y(n12) );
  INVX1 U16 ( .A(n13), .Y(n14) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(\S<2> ), .Y(n16) );
  INVX1 U19 ( .A(\S<1> ), .Y(n17) );
  INVX1 U20 ( .A(n20), .Y(n18) );
  INVX1 U21 ( .A(In), .Y(n19) );
  INVX1 U22 ( .A(n14), .Y(n22) );
  NOR3X1 U23 ( .A(\S<1> ), .B(n3), .C(n21), .Y(Out5) );
  NOR3X1 U24 ( .A(\S<1> ), .B(n3), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U25 ( .A(\S<1> ), .B(n22), .C(n21), .Y(Out1) );
  NOR3X1 U26 ( .A(\S<1> ), .B(n22), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_14 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n2, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  AND2X1 U1 ( .A(n13), .B(n2), .Y(Out2) );
  INVX8 U2 ( .A(\S<0> ), .Y(n2) );
  AND2X1 U3 ( .A(n13), .B(\S<0> ), .Y(Out3) );
  INVX1 U4 ( .A(n6), .Y(Out6) );
  OR2X1 U5 ( .A(n11), .B(\S<0> ), .Y(n6) );
  OR2X1 U6 ( .A(n14), .B(\S<2> ), .Y(n5) );
  AND2X1 U7 ( .A(\S<1> ), .B(n9), .Y(n10) );
  AND2X2 U8 ( .A(n10), .B(\S<0> ), .Y(Out7) );
  INVX1 U9 ( .A(\S<0> ), .Y(n17) );
  OR2X2 U10 ( .A(n15), .B(n16), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  INVX1 U12 ( .A(n10), .Y(n11) );
  NOR3X1 U13 ( .A(\S<2> ), .B(n12), .C(n14), .Y(n13) );
  INVX1 U14 ( .A(\S<1> ), .Y(n12) );
  INVX1 U15 ( .A(In), .Y(n14) );
  INVX1 U16 ( .A(In), .Y(n15) );
  INVX1 U17 ( .A(\S<2> ), .Y(n16) );
  INVX1 U18 ( .A(n9), .Y(n18) );
  NOR3X1 U19 ( .A(\S<1> ), .B(n18), .C(n17), .Y(Out5) );
  NOR3X1 U20 ( .A(\S<1> ), .B(n18), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U21 ( .A(\S<1> ), .B(n5), .C(n17), .Y(Out1) );
  NOR3X1 U22 ( .A(\S<1> ), .B(n5), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to8_15 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n5, n6, n7, n8, n10, n12, n14, n15, n16, n17, n18, n19;

  AND2X1 U1 ( .A(n3), .B(n18), .Y(Out2) );
  OR2X1 U2 ( .A(n17), .B(\S<0> ), .Y(n1) );
  OR2X1 U3 ( .A(n15), .B(\S<2> ), .Y(n5) );
  INVX1 U4 ( .A(\S<2> ), .Y(n19) );
  INVX1 U5 ( .A(\S<0> ), .Y(n18) );
  AND2X1 U6 ( .A(n19), .B(\S<1> ), .Y(n2) );
  AND2X2 U7 ( .A(In), .B(n2), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(n6) );
  OR2X2 U9 ( .A(n17), .B(n14), .Y(n7) );
  OR2X2 U10 ( .A(n7), .B(n18), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(Out7) );
  OR2X2 U12 ( .A(n1), .B(n14), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(Out6) );
  OR2X2 U14 ( .A(n6), .B(n18), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(Out3) );
  OR2X2 U16 ( .A(n16), .B(n19), .Y(n14) );
  INVX1 U17 ( .A(In), .Y(n15) );
  INVX1 U18 ( .A(In), .Y(n16) );
  INVX1 U19 ( .A(\S<1> ), .Y(n17) );
  NOR3X1 U20 ( .A(\S<1> ), .B(n14), .C(n18), .Y(Out5) );
  NOR3X1 U21 ( .A(\S<1> ), .B(n14), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U22 ( .A(\S<1> ), .B(n5), .C(n18), .Y(Out1) );
  NOR3X1 U23 ( .A(\S<1> ), .B(n5), .C(\S<0> ), .Y(Out0) );
endmodule


module demux1to2_17 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_18 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_19 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_20 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(S), .Y(n2) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_21 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_22 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(S), .Y(n2) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_23 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_24 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(S), .Y(n2) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_25 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_26 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_27 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_28 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_29 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_30 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_31 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_32 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_15 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  BUFX2 U3 ( .A(In), .Y(n1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_14 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_13 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_12 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  BUFX2 U3 ( .A(In), .Y(n1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_11 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_10 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  AND2X2 U1 ( .A(In), .B(S), .Y(Out1) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
endmodule


module demux1to2_9 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_8 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_7 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_6 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_5 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_4 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_3 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_2 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_1 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  AND2X2 U1 ( .A(In), .B(S), .Y(Out1) );
  INVX1 U2 ( .A(In), .Y(n1) );
endmodule


module demux1to2_0 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to4_16_1 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<1> , \S<0> }), .Out0({
        \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , 
        \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , 
        \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , 
        \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , 
        \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , 
        \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , \Out2<14> , 
        \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , 
        \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , 
        \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , \Out3<13> , 
        \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , 
        \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , 
        \Out3<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> ;
  wire   n23, n24, n25, n26, n27, n28, n1, n2, n3, n4, n5, n11, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22;

  demux1to4_17 \demux[0]  ( .In(\In<0> ), .S({n21, n4}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ) );
  demux1to4_18 \demux[1]  ( .In(\In<1> ), .S({n21, n14}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(n28) );
  demux1to4_19 \demux[2]  ( .In(\In<2> ), .S({n1, n15}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ) );
  demux1to4_20 \demux[3]  ( .In(\In<3> ), .S({n21, n19}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(n27) );
  demux1to4_21 \demux[4]  ( .In(\In<4> ), .S({n13, n4}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ) );
  demux1to4_22 \demux[5]  ( .In(\In<5> ), .S({n1, n16}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ) );
  demux1to4_23 \demux[6]  ( .In(\In<6> ), .S({n1, n4}), .Out0(\Out0<6> ), 
        .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ) );
  demux1to4_24 \demux[7]  ( .In(\In<7> ), .S({n21, n4}), .Out0(\Out0<7> ), 
        .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ) );
  demux1to4_25 \demux[8]  ( .In(\In<8> ), .S({n13, n18}), .Out0(\Out0<8> ), 
        .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(n26) );
  demux1to4_26 \demux[9]  ( .In(\In<9> ), .S({n13, n3}), .Out0(\Out0<9> ), 
        .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(n25) );
  demux1to4_27 \demux[10]  ( .In(\In<10> ), .S({n1, n17}), .Out0(\Out0<10> ), 
        .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(n24) );
  demux1to4_28 \demux[11]  ( .In(\In<11> ), .S({n13, n16}), .Out0(\Out0<11> ), 
        .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ) );
  demux1to4_29 \demux[12]  ( .In(\In<12> ), .S({n1, n17}), .Out0(\Out0<12> ), 
        .Out1(\Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ) );
  demux1to4_30 \demux[13]  ( .In(\In<13> ), .S({n1, n4}), .Out0(\Out0<13> ), 
        .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ) );
  demux1to4_31 \demux[14]  ( .In(\In<14> ), .S({n13, n16}), .Out0(\Out0<14> ), 
        .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(n23) );
  demux1to4_32 \demux[15]  ( .In(\In<15> ), .S({n13, n17}), .Out0(\Out0<15> ), 
        .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ) );
  INVX8 U1 ( .A(n22), .Y(n1) );
  INVX2 U2 ( .A(n2), .Y(n17) );
  INVX2 U3 ( .A(n2), .Y(n16) );
  INVX1 U4 ( .A(n2), .Y(n18) );
  INVX1 U5 ( .A(n20), .Y(n15) );
  INVX1 U6 ( .A(\S<0> ), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  INVX4 U8 ( .A(n20), .Y(n4) );
  INVX1 U9 ( .A(\S<0> ), .Y(n5) );
  INVX8 U10 ( .A(n22), .Y(n13) );
  INVX8 U11 ( .A(n22), .Y(n21) );
  INVX1 U12 ( .A(\S<0> ), .Y(n20) );
  BUFX2 U13 ( .A(n23), .Y(\Out3<14> ) );
  BUFX2 U14 ( .A(n25), .Y(\Out3<9> ) );
  BUFX2 U15 ( .A(n26), .Y(\Out3<8> ) );
  BUFX2 U16 ( .A(n27), .Y(\Out3<3> ) );
  BUFX2 U17 ( .A(n28), .Y(\Out3<1> ) );
  INVX1 U18 ( .A(n24), .Y(n11) );
  INVX1 U19 ( .A(n11), .Y(\Out3<10> ) );
  INVX1 U20 ( .A(n5), .Y(n14) );
  INVX1 U21 ( .A(n5), .Y(n19) );
  INVX8 U22 ( .A(\S<1> ), .Y(n22) );
endmodule


module demux1to4_16_0 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<1> , \S<0> }), .Out0({
        \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , 
        \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , 
        \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , 
        \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , 
        \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , 
        \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , \Out2<14> , 
        \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , 
        \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , 
        \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , \Out3<13> , 
        \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , 
        \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , 
        \Out3<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> ;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n1, n2, n3, n27,
         n29, n30, n31, n32, n33;

  demux1to4_15 \demux[0]  ( .In(\In<0> ), .S({n31, n2}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(n43), .Out3(n57) );
  demux1to4_14 \demux[1]  ( .In(\In<1> ), .S({n31, n1}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(n56) );
  demux1to4_13 \demux[2]  ( .In(\In<2> ), .S({n31, n3}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(n42), .Out3(n55) );
  demux1to4_12 \demux[3]  ( .In(\In<3> ), .S({n31, n1}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(n54) );
  demux1to4_11 \demux[4]  ( .In(\In<4> ), .S({n32, n2}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(n41), .Out3(n53) );
  demux1to4_10 \demux[5]  ( .In(\In<5> ), .S({n31, n2}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(n40), .Out3(n52) );
  demux1to4_9 \demux[6]  ( .In(\In<6> ), .S({n31, n2}), .Out0(\Out0<6> ), 
        .Out1(\Out1<6> ), .Out2(n39), .Out3(n51) );
  demux1to4_8 \demux[7]  ( .In(\In<7> ), .S({n31, n3}), .Out0(\Out0<7> ), 
        .Out1(\Out1<7> ), .Out2(n38), .Out3(n50) );
  demux1to4_7 \demux[8]  ( .In(\In<8> ), .S({n32, n2}), .Out0(\Out0<8> ), 
        .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ) );
  demux1to4_6 \demux[9]  ( .In(\In<9> ), .S({n32, n2}), .Out0(\Out0<9> ), 
        .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(n49) );
  demux1to4_5 \demux[10]  ( .In(\In<10> ), .S({n31, n2}), .Out0(\Out0<10> ), 
        .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ) );
  demux1to4_4 \demux[11]  ( .In(\In<11> ), .S({n32, n30}), .Out0(\Out0<11> ), 
        .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(n48) );
  demux1to4_3 \demux[12]  ( .In(\In<12> ), .S({n32, n30}), .Out0(n36), .Out1(
        \Out1<12> ), .Out2(\Out2<12> ), .Out3(n47) );
  demux1to4_2 \demux[13]  ( .In(\In<13> ), .S({n32, n30}), .Out0(n35), .Out1(
        \Out1<13> ), .Out2(\Out2<13> ), .Out3(n46) );
  demux1to4_1 \demux[14]  ( .In(\In<14> ), .S({n32, n2}), .Out0(n34), .Out1(
        \Out1<14> ), .Out2(\Out2<14> ), .Out3(n45) );
  demux1to4_0 \demux[15]  ( .In(\In<15> ), .S({n32, n30}), .Out0(\Out0<15> ), 
        .Out1(\Out1<15> ), .Out2(n37), .Out3(n44) );
  INVX2 U1 ( .A(n29), .Y(n1) );
  INVX2 U2 ( .A(\S<0> ), .Y(n29) );
  INVX2 U3 ( .A(\S<1> ), .Y(n33) );
  INVX1 U4 ( .A(n29), .Y(n3) );
  INVX4 U5 ( .A(n29), .Y(n2) );
  INVX1 U6 ( .A(n29), .Y(n30) );
  BUFX2 U7 ( .A(n44), .Y(\Out3<15> ) );
  BUFX2 U8 ( .A(n45), .Y(\Out3<14> ) );
  BUFX2 U9 ( .A(n46), .Y(\Out3<13> ) );
  BUFX2 U10 ( .A(n47), .Y(\Out3<12> ) );
  BUFX2 U11 ( .A(n48), .Y(\Out3<11> ) );
  BUFX2 U12 ( .A(n49), .Y(\Out3<9> ) );
  BUFX2 U13 ( .A(n50), .Y(\Out3<7> ) );
  BUFX2 U14 ( .A(n51), .Y(\Out3<6> ) );
  BUFX2 U15 ( .A(n52), .Y(\Out3<5> ) );
  BUFX2 U16 ( .A(n53), .Y(\Out3<4> ) );
  BUFX2 U17 ( .A(n54), .Y(\Out3<3> ) );
  BUFX2 U18 ( .A(n55), .Y(\Out3<2> ) );
  BUFX2 U19 ( .A(n56), .Y(\Out3<1> ) );
  BUFX2 U20 ( .A(n57), .Y(\Out3<0> ) );
  BUFX2 U21 ( .A(n34), .Y(\Out0<14> ) );
  BUFX2 U22 ( .A(n35), .Y(\Out0<13> ) );
  BUFX2 U23 ( .A(n36), .Y(\Out0<12> ) );
  BUFX2 U24 ( .A(n37), .Y(\Out2<15> ) );
  BUFX2 U25 ( .A(n39), .Y(\Out2<6> ) );
  BUFX2 U26 ( .A(n40), .Y(\Out2<5> ) );
  BUFX2 U27 ( .A(n41), .Y(\Out2<4> ) );
  BUFX2 U28 ( .A(n42), .Y(\Out2<2> ) );
  BUFX2 U29 ( .A(n43), .Y(\Out2<0> ) );
  INVX1 U30 ( .A(n38), .Y(n27) );
  INVX1 U31 ( .A(n27), .Y(\Out2<7> ) );
  INVX4 U32 ( .A(n33), .Y(n32) );
  INVX8 U33 ( .A(n33), .Y(n31) );
endmodule


module cla16_0 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \P<3> , \P<2> , \P<1> , \P<0> , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  cla4_3 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(n17), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(n28) );
  cla4_2 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n27), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_1 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n29), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_0 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n6), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  INVX1 U1 ( .A(\G<3> ), .Y(n26) );
  INVX1 U2 ( .A(n16), .Y(n1) );
  INVX1 U3 ( .A(n16), .Y(n2) );
  OAI21X1 U4 ( .A(n25), .B(n24), .C(n1), .Y(n3) );
  INVX1 U5 ( .A(n17), .Y(n25) );
  BUFX2 U6 ( .A(n6), .Y(n4) );
  BUFX2 U7 ( .A(\P<2> ), .Y(n5) );
  OR2X2 U8 ( .A(n8), .B(n7), .Y(n6) );
  OR2X2 U9 ( .A(n14), .B(n15), .Y(n7) );
  AND2X2 U10 ( .A(\G<1> ), .B(n5), .Y(n8) );
  AND2X2 U11 ( .A(n26), .B(n19), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Cout) );
  BUFX2 U13 ( .A(n23), .Y(n11) );
  AND2X2 U14 ( .A(n16), .B(\P<1> ), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(n13) );
  INVX1 U16 ( .A(n21), .Y(n14) );
  INVX1 U17 ( .A(n20), .Y(n15) );
  BUFX2 U18 ( .A(n28), .Y(n16) );
  BUFX2 U19 ( .A(Cin), .Y(n17) );
  AND2X2 U20 ( .A(\P<3> ), .B(n4), .Y(n18) );
  INVX1 U21 ( .A(n18), .Y(n19) );
  INVX1 U22 ( .A(\G<2> ), .Y(n20) );
  INVX1 U23 ( .A(\G<1> ), .Y(n22) );
  NAND3X1 U24 ( .A(\P<1> ), .B(\P<2> ), .C(n3), .Y(n21) );
  NAND3X1 U25 ( .A(n17), .B(\P<1> ), .C(\P<0> ), .Y(n23) );
  NAND3X1 U26 ( .A(n11), .B(n13), .C(n22), .Y(n29) );
  INVX2 U27 ( .A(\P<0> ), .Y(n24) );
  OAI21X1 U28 ( .A(n25), .B(n24), .C(n2), .Y(n27) );
endmodule


module mux4to1_16_0 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n3, n5, n7, n9, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135;

  AND2X1 U1 ( .A(n35), .B(n41), .Y(n64) );
  AND2X1 U2 ( .A(n27), .B(n39), .Y(n56) );
  AND2X1 U3 ( .A(n54), .B(n75), .Y(n13) );
  AND2X1 U4 ( .A(n55), .B(n49), .Y(n14) );
  AND2X2 U5 ( .A(n82), .B(n13), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(\Out<1> ) );
  AND2X2 U7 ( .A(n14), .B(n51), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(\Out<8> ) );
  AND2X2 U9 ( .A(n15), .B(n47), .Y(n5) );
  INVX1 U10 ( .A(n5), .Y(\Out<6> ) );
  AND2X2 U11 ( .A(n78), .B(n42), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(\Out<5> ) );
  AND2X2 U13 ( .A(n79), .B(n45), .Y(n9) );
  INVX1 U14 ( .A(n9), .Y(\Out<7> ) );
  AND2X2 U15 ( .A(n80), .B(n53), .Y(n11) );
  INVX1 U16 ( .A(n11), .Y(\Out<11> ) );
  AND2X2 U17 ( .A(n19), .B(n43), .Y(n15) );
  AND2X2 U18 ( .A(\S<0> ), .B(\S<1> ), .Y(n16) );
  AND2X2 U19 ( .A(\S<0> ), .B(n109), .Y(n17) );
  AND2X2 U20 ( .A(\InB<6> ), .B(n17), .Y(n18) );
  INVX1 U21 ( .A(n18), .Y(n19) );
  AND2X2 U22 ( .A(\InB<10> ), .B(n17), .Y(n20) );
  INVX1 U23 ( .A(n20), .Y(n21) );
  AND2X2 U24 ( .A(\InD<11> ), .B(n16), .Y(n22) );
  INVX1 U25 ( .A(n22), .Y(n23) );
  AND2X2 U26 ( .A(\InB<13> ), .B(n17), .Y(n24) );
  INVX1 U27 ( .A(n24), .Y(n25) );
  AND2X2 U28 ( .A(\InD<9> ), .B(n16), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  AND2X2 U30 ( .A(\InD<10> ), .B(n16), .Y(n28) );
  INVX1 U31 ( .A(n28), .Y(n29) );
  AND2X2 U32 ( .A(\InB<11> ), .B(n17), .Y(n30) );
  INVX1 U33 ( .A(n30), .Y(n31) );
  AND2X2 U34 ( .A(\InD<13> ), .B(n16), .Y(n32) );
  INVX1 U35 ( .A(n32), .Y(n33) );
  AND2X2 U36 ( .A(\InD<14> ), .B(n16), .Y(n34) );
  INVX1 U37 ( .A(n34), .Y(n35) );
  AND2X2 U38 ( .A(\InD<15> ), .B(n16), .Y(n36) );
  INVX1 U39 ( .A(n36), .Y(n37) );
  AND2X2 U40 ( .A(\InB<9> ), .B(n17), .Y(n38) );
  INVX1 U41 ( .A(n38), .Y(n39) );
  AND2X2 U42 ( .A(\InB<14> ), .B(n17), .Y(n40) );
  INVX1 U43 ( .A(n40), .Y(n41) );
  BUFX2 U44 ( .A(n117), .Y(n42) );
  BUFX2 U45 ( .A(n118), .Y(n43) );
  OR2X2 U46 ( .A(n107), .B(n108), .Y(n44) );
  INVX1 U47 ( .A(n44), .Y(n45) );
  AND2X2 U48 ( .A(\InA<6> ), .B(n126), .Y(n46) );
  INVX1 U49 ( .A(n46), .Y(n47) );
  AND2X2 U50 ( .A(\InC<8> ), .B(n132), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n49) );
  AND2X2 U52 ( .A(\InA<8> ), .B(n126), .Y(n50) );
  INVX1 U53 ( .A(n50), .Y(n51) );
  AND2X2 U54 ( .A(\InA<11> ), .B(n126), .Y(n52) );
  INVX1 U55 ( .A(n52), .Y(n53) );
  BUFX2 U56 ( .A(n112), .Y(n54) );
  BUFX2 U57 ( .A(n120), .Y(n55) );
  INVX1 U58 ( .A(n56), .Y(n57) );
  AND2X2 U59 ( .A(n29), .B(n21), .Y(n58) );
  INVX1 U60 ( .A(n58), .Y(n59) );
  AND2X2 U61 ( .A(n31), .B(n23), .Y(n60) );
  INVX1 U62 ( .A(n60), .Y(n61) );
  AND2X2 U63 ( .A(n33), .B(n25), .Y(n62) );
  INVX1 U64 ( .A(n62), .Y(n63) );
  INVX1 U65 ( .A(n64), .Y(n65) );
  AND2X2 U66 ( .A(n37), .B(n77), .Y(n66) );
  INVX1 U67 ( .A(n66), .Y(n67) );
  AND2X2 U68 ( .A(\InA<3> ), .B(n126), .Y(n68) );
  INVX1 U69 ( .A(n68), .Y(n69) );
  AND2X2 U70 ( .A(\InA<4> ), .B(n126), .Y(n70) );
  INVX1 U71 ( .A(n70), .Y(n71) );
  AND2X2 U72 ( .A(n126), .B(\InA<12> ), .Y(n72) );
  INVX1 U73 ( .A(n72), .Y(n73) );
  AND2X2 U74 ( .A(\InB<1> ), .B(n17), .Y(n74) );
  INVX1 U75 ( .A(n74), .Y(n75) );
  AND2X2 U76 ( .A(\InB<15> ), .B(n17), .Y(n76) );
  INVX1 U77 ( .A(n76), .Y(n77) );
  BUFX2 U78 ( .A(n116), .Y(n78) );
  BUFX2 U79 ( .A(n119), .Y(n79) );
  BUFX2 U80 ( .A(n125), .Y(n80) );
  AND2X2 U81 ( .A(\InA<1> ), .B(n126), .Y(n81) );
  INVX1 U82 ( .A(n81), .Y(n82) );
  BUFX2 U83 ( .A(n111), .Y(n83) );
  BUFX2 U84 ( .A(n113), .Y(n84) );
  BUFX2 U85 ( .A(n114), .Y(n85) );
  BUFX2 U86 ( .A(n115), .Y(n86) );
  BUFX2 U87 ( .A(n127), .Y(n87) );
  AND2X2 U88 ( .A(\InA<0> ), .B(n126), .Y(n88) );
  INVX1 U89 ( .A(n88), .Y(n89) );
  AND2X2 U90 ( .A(\InA<2> ), .B(n126), .Y(n90) );
  INVX1 U91 ( .A(n90), .Y(n91) );
  AND2X2 U92 ( .A(\InB<12> ), .B(n17), .Y(n92) );
  INVX1 U93 ( .A(n92), .Y(n93) );
  AND2X2 U94 ( .A(\InB<0> ), .B(n17), .Y(n94) );
  INVX1 U95 ( .A(n94), .Y(n95) );
  AND2X2 U96 ( .A(\InB<2> ), .B(n17), .Y(n96) );
  INVX1 U97 ( .A(n96), .Y(n97) );
  AND2X2 U98 ( .A(\InB<3> ), .B(n17), .Y(n98) );
  INVX1 U99 ( .A(n98), .Y(n99) );
  AND2X2 U100 ( .A(\InB<4> ), .B(n17), .Y(n100) );
  INVX1 U101 ( .A(n100), .Y(n101) );
  BUFX2 U102 ( .A(n122), .Y(n102) );
  BUFX2 U103 ( .A(n124), .Y(n103) );
  BUFX2 U104 ( .A(n129), .Y(n104) );
  BUFX2 U105 ( .A(n131), .Y(n105) );
  BUFX2 U106 ( .A(n134), .Y(n106) );
  INVX1 U107 ( .A(\InA<14> ), .Y(n130) );
  INVX1 U108 ( .A(\S<1> ), .Y(n109) );
  AND2X2 U109 ( .A(\InA<7> ), .B(n126), .Y(n107) );
  AND2X2 U110 ( .A(\InB<7> ), .B(n17), .Y(n108) );
  INVX1 U111 ( .A(\InA<15> ), .Y(n133) );
  INVX1 U112 ( .A(\InA<9> ), .Y(n121) );
  INVX1 U113 ( .A(\InA<10> ), .Y(n123) );
  INVX1 U114 ( .A(\InA<13> ), .Y(n128) );
  INVX8 U115 ( .A(n110), .Y(n132) );
  INVX4 U116 ( .A(n135), .Y(n126) );
  OR2X2 U117 ( .A(n109), .B(\S<0> ), .Y(n110) );
  AOI22X1 U118 ( .A(\InD<0> ), .B(n16), .C(\InC<0> ), .D(n132), .Y(n111) );
  OR2X2 U119 ( .A(\S<1> ), .B(\S<0> ), .Y(n135) );
  NAND3X1 U120 ( .A(n83), .B(n89), .C(n95), .Y(\Out<0> ) );
  AOI22X1 U121 ( .A(\InD<1> ), .B(n16), .C(\InC<1> ), .D(n132), .Y(n112) );
  AOI22X1 U122 ( .A(\InD<2> ), .B(n16), .C(\InC<2> ), .D(n132), .Y(n113) );
  NAND3X1 U123 ( .A(n84), .B(n91), .C(n97), .Y(\Out<2> ) );
  AOI22X1 U124 ( .A(\InD<3> ), .B(n16), .C(\InC<3> ), .D(n132), .Y(n114) );
  NAND3X1 U125 ( .A(n85), .B(n69), .C(n99), .Y(\Out<3> ) );
  AOI22X1 U126 ( .A(\InD<4> ), .B(n16), .C(\InC<4> ), .D(n132), .Y(n115) );
  NAND3X1 U127 ( .A(n86), .B(n101), .C(n71), .Y(\Out<4> ) );
  AOI22X1 U128 ( .A(n126), .B(\InA<5> ), .C(\InB<5> ), .D(n17), .Y(n117) );
  AOI22X1 U129 ( .A(\InD<5> ), .B(n16), .C(\InC<5> ), .D(n132), .Y(n116) );
  AOI22X1 U130 ( .A(\InD<6> ), .B(n16), .C(\InC<6> ), .D(n132), .Y(n118) );
  AOI22X1 U131 ( .A(\InD<7> ), .B(n16), .C(\InC<7> ), .D(n132), .Y(n119) );
  AOI22X1 U132 ( .A(\InD<8> ), .B(n16), .C(\InB<8> ), .D(n17), .Y(n120) );
  AOI21X1 U133 ( .A(\InC<9> ), .B(n132), .C(n57), .Y(n122) );
  AOI22X1 U134 ( .A(n135), .B(n102), .C(n102), .D(n121), .Y(\Out<9> ) );
  AOI21X1 U135 ( .A(\InC<10> ), .B(n132), .C(n59), .Y(n124) );
  AOI22X1 U136 ( .A(n135), .B(n103), .C(n103), .D(n123), .Y(\Out<10> ) );
  AOI21X1 U137 ( .A(\InC<11> ), .B(n132), .C(n61), .Y(n125) );
  AOI22X1 U138 ( .A(\InD<12> ), .B(n16), .C(\InC<12> ), .D(n132), .Y(n127) );
  NAND3X1 U139 ( .A(n87), .B(n93), .C(n73), .Y(\Out<12> ) );
  AOI21X1 U140 ( .A(\InC<13> ), .B(n132), .C(n63), .Y(n129) );
  AOI22X1 U141 ( .A(n135), .B(n104), .C(n104), .D(n128), .Y(\Out<13> ) );
  AOI21X1 U142 ( .A(\InC<14> ), .B(n132), .C(n65), .Y(n131) );
  AOI22X1 U143 ( .A(n135), .B(n105), .C(n105), .D(n130), .Y(\Out<14> ) );
  AOI21X1 U144 ( .A(\InC<15> ), .B(n132), .C(n67), .Y(n134) );
  AOI22X1 U145 ( .A(n135), .B(n106), .C(n106), .D(n133), .Y(\Out<15> ) );
endmodule


module lshifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), Rot_sel, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , Rot_sel;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n20, n21, n22, n23, n25, n27, n29, n31, n33, n34, n35, n37, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n128, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248;

  INVX1 U2 ( .A(\Cnt<2> ), .Y(n179) );
  INVX1 U3 ( .A(\Cnt<1> ), .Y(n184) );
  INVX1 U4 ( .A(\In<2> ), .Y(n208) );
  INVX1 U5 ( .A(\In<1> ), .Y(n195) );
  INVX1 U6 ( .A(Rot_sel), .Y(n172) );
  INVX2 U7 ( .A(n172), .Y(n171) );
  AND2X2 U8 ( .A(\Cnt<3> ), .B(n179), .Y(n1) );
  AND2X2 U9 ( .A(n70), .B(n122), .Y(n2) );
  INVX1 U10 ( .A(n2), .Y(\Out<1> ) );
  AND2X2 U11 ( .A(n11), .B(n97), .Y(n4) );
  INVX1 U12 ( .A(n4), .Y(n5) );
  AND2X2 U13 ( .A(\Cnt<0> ), .B(n184), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(n7) );
  AND2X2 U15 ( .A(n171), .B(n115), .Y(n8) );
  AND2X2 U16 ( .A(n171), .B(n1), .Y(n9) );
  AND2X2 U17 ( .A(n184), .B(n206), .Y(n10) );
  INVX1 U18 ( .A(n10), .Y(n11) );
  AND2X2 U19 ( .A(n71), .B(n59), .Y(n12) );
  AND2X2 U20 ( .A(n73), .B(n60), .Y(n13) );
  AND2X2 U21 ( .A(n72), .B(n61), .Y(n14) );
  INVX1 U22 ( .A(n14), .Y(\Out<2> ) );
  AND2X2 U23 ( .A(n75), .B(n62), .Y(n16) );
  AND2X2 U24 ( .A(n74), .B(n63), .Y(n17) );
  INVX1 U25 ( .A(n17), .Y(\Out<3> ) );
  AND2X2 U26 ( .A(n8), .B(n137), .Y(n19) );
  INVX1 U27 ( .A(n19), .Y(n20) );
  AND2X2 U28 ( .A(n245), .B(n5), .Y(n21) );
  INVX1 U29 ( .A(n21), .Y(n22) );
  AND2X2 U30 ( .A(n76), .B(n64), .Y(n23) );
  INVX1 U31 ( .A(n23), .Y(\Out<7> ) );
  AND2X2 U32 ( .A(n77), .B(n65), .Y(n25) );
  INVX1 U33 ( .A(n25), .Y(\Out<8> ) );
  AND2X2 U34 ( .A(n78), .B(n66), .Y(n27) );
  INVX1 U35 ( .A(n27), .Y(\Out<10> ) );
  AND2X2 U36 ( .A(n79), .B(n118), .Y(n29) );
  INVX1 U37 ( .A(n29), .Y(\Out<11> ) );
  AND2X2 U38 ( .A(n80), .B(n67), .Y(n31) );
  INVX1 U39 ( .A(n31), .Y(\Out<12> ) );
  AND2X2 U40 ( .A(n1), .B(n114), .Y(n33) );
  INVX1 U41 ( .A(n33), .Y(n34) );
  AND2X2 U42 ( .A(n81), .B(n68), .Y(n35) );
  INVX1 U43 ( .A(n35), .Y(\Out<14> ) );
  AND2X2 U44 ( .A(n123), .B(n69), .Y(n37) );
  INVX1 U45 ( .A(n37), .Y(\Out<15> ) );
  BUFX2 U46 ( .A(n187), .Y(n39) );
  BUFX2 U47 ( .A(n191), .Y(n40) );
  BUFX2 U48 ( .A(n213), .Y(n41) );
  BUFX2 U49 ( .A(n217), .Y(n42) );
  BUFX2 U50 ( .A(n228), .Y(n43) );
  INVX1 U51 ( .A(n96), .Y(n44) );
  BUFX2 U52 ( .A(n175), .Y(n45) );
  BUFX2 U53 ( .A(n177), .Y(n46) );
  BUFX2 U54 ( .A(n180), .Y(n47) );
  BUFX2 U55 ( .A(n186), .Y(n48) );
  BUFX2 U56 ( .A(n190), .Y(n49) );
  BUFX2 U57 ( .A(n200), .Y(n50) );
  BUFX2 U58 ( .A(n202), .Y(n51) );
  BUFX2 U59 ( .A(n212), .Y(n52) );
  BUFX2 U60 ( .A(n216), .Y(n53) );
  BUFX2 U61 ( .A(n227), .Y(n54) );
  BUFX2 U62 ( .A(n194), .Y(n55) );
  BUFX2 U63 ( .A(n207), .Y(n56) );
  AND2X2 U64 ( .A(\In<15> ), .B(n220), .Y(n57) );
  INVX1 U65 ( .A(n57), .Y(n58) );
  BUFX2 U66 ( .A(n196), .Y(n59) );
  BUFX2 U67 ( .A(n204), .Y(n60) );
  BUFX2 U68 ( .A(n210), .Y(n61) );
  BUFX2 U69 ( .A(n221), .Y(n62) );
  BUFX2 U70 ( .A(n223), .Y(n63) );
  BUFX2 U71 ( .A(n229), .Y(n64) );
  BUFX2 U72 ( .A(n231), .Y(n65) );
  BUFX2 U73 ( .A(n234), .Y(n66) );
  BUFX2 U74 ( .A(n238), .Y(n67) );
  BUFX2 U75 ( .A(n243), .Y(n68) );
  BUFX2 U76 ( .A(n247), .Y(n69) );
  BUFX2 U77 ( .A(n199), .Y(n70) );
  BUFX2 U78 ( .A(n197), .Y(n71) );
  BUFX2 U79 ( .A(n211), .Y(n72) );
  BUFX2 U80 ( .A(n205), .Y(n73) );
  BUFX2 U81 ( .A(n224), .Y(n74) );
  BUFX2 U82 ( .A(n222), .Y(n75) );
  BUFX2 U83 ( .A(n230), .Y(n76) );
  BUFX2 U84 ( .A(n232), .Y(n77) );
  BUFX2 U85 ( .A(n235), .Y(n78) );
  BUFX2 U86 ( .A(n237), .Y(n79) );
  BUFX2 U87 ( .A(n239), .Y(n80) );
  BUFX2 U88 ( .A(n244), .Y(n81) );
  AND2X2 U89 ( .A(n1), .B(n240), .Y(n82) );
  INVX1 U90 ( .A(n82), .Y(n83) );
  AND2X2 U91 ( .A(n115), .B(n240), .Y(n84) );
  INVX1 U92 ( .A(n84), .Y(n85) );
  AND2X2 U93 ( .A(n95), .B(n94), .Y(n86) );
  INVX1 U94 ( .A(n86), .Y(n87) );
  AND2X2 U95 ( .A(\In<15> ), .B(n171), .Y(n88) );
  INVX1 U96 ( .A(n88), .Y(n89) );
  AND2X2 U97 ( .A(n245), .B(n240), .Y(n90) );
  INVX1 U98 ( .A(n90), .Y(n91) );
  BUFX2 U99 ( .A(n225), .Y(n92) );
  BUFX2 U100 ( .A(n241), .Y(n93) );
  BUFX2 U101 ( .A(n214), .Y(n94) );
  BUFX2 U102 ( .A(n215), .Y(n95) );
  AND2X2 U103 ( .A(n170), .B(n171), .Y(n96) );
  INVX1 U104 ( .A(n96), .Y(n97) );
  AND2X2 U105 ( .A(n44), .B(n11), .Y(n98) );
  INVX1 U106 ( .A(n98), .Y(n99) );
  INVX1 U107 ( .A(n98), .Y(n100) );
  AND2X1 U108 ( .A(\Cnt<0> ), .B(\Cnt<1> ), .Y(n101) );
  INVX2 U109 ( .A(n101), .Y(n102) );
  AND2X2 U110 ( .A(n171), .B(n245), .Y(n103) );
  INVX1 U111 ( .A(n176), .Y(n104) );
  INVX1 U112 ( .A(n104), .Y(n105) );
  INVX1 U113 ( .A(n178), .Y(n106) );
  INVX1 U114 ( .A(n106), .Y(n107) );
  INVX1 U115 ( .A(n181), .Y(n108) );
  INVX1 U116 ( .A(n108), .Y(n109) );
  INVX1 U117 ( .A(n201), .Y(n110) );
  INVX1 U118 ( .A(n110), .Y(n111) );
  INVX1 U119 ( .A(n203), .Y(n112) );
  INVX1 U120 ( .A(n112), .Y(n113) );
  OR2X2 U121 ( .A(n168), .B(n169), .Y(n114) );
  AND2X2 U122 ( .A(\Cnt<3> ), .B(\Cnt<2> ), .Y(n115) );
  INVX1 U123 ( .A(n4), .Y(n116) );
  INVX1 U124 ( .A(n236), .Y(n117) );
  INVX1 U125 ( .A(n117), .Y(n118) );
  INVX1 U126 ( .A(n233), .Y(n119) );
  INVX1 U127 ( .A(n119), .Y(n120) );
  INVX1 U128 ( .A(n198), .Y(n121) );
  INVX1 U129 ( .A(n121), .Y(n122) );
  BUFX2 U130 ( .A(n248), .Y(n123) );
  AND2X2 U131 ( .A(n8), .B(n143), .Y(n124) );
  INVX1 U132 ( .A(n124), .Y(n125) );
  AND2X2 U133 ( .A(n39), .B(n48), .Y(n126) );
  INVX1 U134 ( .A(n126), .Y(\Out<0> ) );
  AND2X2 U135 ( .A(n43), .B(n54), .Y(n128) );
  INVX1 U136 ( .A(n128), .Y(\Out<6> ) );
  AND2X2 U137 ( .A(n8), .B(n140), .Y(n130) );
  INVX1 U138 ( .A(n130), .Y(n131) );
  INVX1 U139 ( .A(n226), .Y(n132) );
  INVX1 U140 ( .A(n132), .Y(n133) );
  INVX8 U141 ( .A(n7), .Y(n134) );
  INVX1 U142 ( .A(n86), .Y(n135) );
  BUFX2 U143 ( .A(n102), .Y(n136) );
  INVX1 U144 ( .A(n139), .Y(n137) );
  INVX1 U145 ( .A(n139), .Y(n138) );
  AND2X2 U146 ( .A(n109), .B(n47), .Y(n139) );
  INVX1 U147 ( .A(n142), .Y(n140) );
  INVX1 U148 ( .A(n142), .Y(n141) );
  AND2X2 U149 ( .A(n40), .B(n49), .Y(n142) );
  INVX1 U150 ( .A(n12), .Y(n143) );
  INVX1 U151 ( .A(n12), .Y(n144) );
  INVX1 U152 ( .A(n147), .Y(n145) );
  INVX1 U153 ( .A(n147), .Y(n146) );
  AND2X2 U154 ( .A(n111), .B(n50), .Y(n147) );
  INVX1 U155 ( .A(n151), .Y(n148) );
  INVX1 U156 ( .A(n151), .Y(n149) );
  INVX1 U157 ( .A(n151), .Y(n150) );
  AND2X2 U158 ( .A(n41), .B(n52), .Y(n151) );
  INVX1 U159 ( .A(n154), .Y(n152) );
  INVX1 U160 ( .A(n154), .Y(n153) );
  AND2X2 U161 ( .A(n105), .B(n45), .Y(n154) );
  INVX1 U162 ( .A(n13), .Y(n155) );
  INVX1 U163 ( .A(n13), .Y(n156) );
  INVX1 U164 ( .A(n159), .Y(n157) );
  INVX1 U165 ( .A(n159), .Y(n158) );
  AND2X2 U166 ( .A(n42), .B(n53), .Y(n159) );
  INVX1 U167 ( .A(n162), .Y(n160) );
  INVX1 U168 ( .A(n162), .Y(n161) );
  AND2X2 U169 ( .A(n107), .B(n46), .Y(n162) );
  INVX1 U170 ( .A(n165), .Y(n163) );
  INVX1 U171 ( .A(n165), .Y(n164) );
  AND2X2 U172 ( .A(n113), .B(n51), .Y(n165) );
  INVX1 U173 ( .A(n16), .Y(n166) );
  INVX1 U174 ( .A(n16), .Y(n167) );
  INVX1 U175 ( .A(n189), .Y(n168) );
  INVX1 U176 ( .A(n188), .Y(n169) );
  INVX1 U177 ( .A(n185), .Y(n170) );
  INVX4 U178 ( .A(n173), .Y(n245) );
  INVX8 U179 ( .A(n209), .Y(n218) );
  INVX8 U180 ( .A(n174), .Y(n220) );
  INVX4 U181 ( .A(n102), .Y(n219) );
  INVX8 U182 ( .A(n182), .Y(n246) );
  OR2X2 U183 ( .A(n179), .B(\Cnt<3> ), .Y(n173) );
  OR2X2 U184 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n209) );
  AOI22X1 U185 ( .A(\In<12> ), .B(n218), .C(\In<11> ), .D(n134), .Y(n176) );
  OR2X2 U186 ( .A(n184), .B(\Cnt<0> ), .Y(n174) );
  AOI22X1 U187 ( .A(\In<10> ), .B(n220), .C(\In<9> ), .D(n219), .Y(n175) );
  AOI22X1 U188 ( .A(\In<4> ), .B(n218), .C(\In<3> ), .D(n134), .Y(n178) );
  AOI22X1 U189 ( .A(\In<2> ), .B(n220), .C(\In<1> ), .D(n219), .Y(n177) );
  AOI22X1 U190 ( .A(n103), .B(n153), .C(n8), .D(n161), .Y(n187) );
  AOI22X1 U191 ( .A(\In<8> ), .B(n218), .C(\In<7> ), .D(n134), .Y(n181) );
  AOI22X1 U192 ( .A(\In<6> ), .B(n220), .C(\In<5> ), .D(n219), .Y(n180) );
  OR2X2 U193 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n182) );
  AOI22X1 U194 ( .A(\In<14> ), .B(n220), .C(\In<13> ), .D(n219), .Y(n185) );
  INVX2 U195 ( .A(\In<0> ), .Y(n183) );
  MUX2X1 U196 ( .B(n183), .A(n89), .S(\Cnt<0> ), .Y(n206) );
  AOI22X1 U197 ( .A(n9), .B(n138), .C(n246), .D(n116), .Y(n186) );
  AOI22X1 U198 ( .A(\In<5> ), .B(n218), .C(\In<4> ), .D(n134), .Y(n189) );
  AOI22X1 U199 ( .A(\In<3> ), .B(n220), .C(\In<2> ), .D(n219), .Y(n188) );
  AOI22X1 U200 ( .A(\In<13> ), .B(n218), .C(\In<12> ), .D(n134), .Y(n191) );
  AOI22X1 U201 ( .A(\In<11> ), .B(n220), .C(\In<10> ), .D(n219), .Y(n190) );
  AOI22X1 U202 ( .A(n8), .B(n114), .C(n103), .D(n141), .Y(n199) );
  INVX2 U203 ( .A(\In<14> ), .Y(n192) );
  OAI21X1 U204 ( .A(n136), .B(n192), .C(n58), .Y(n193) );
  AOI22X1 U205 ( .A(\In<0> ), .B(n134), .C(n171), .D(n193), .Y(n194) );
  OAI21X1 U206 ( .A(n209), .B(n195), .C(n55), .Y(n240) );
  AOI22X1 U207 ( .A(\In<9> ), .B(n218), .C(\In<8> ), .D(n134), .Y(n197) );
  AOI22X1 U208 ( .A(\In<7> ), .B(n220), .C(\In<6> ), .D(n219), .Y(n196) );
  AOI22X1 U209 ( .A(n246), .B(n240), .C(n9), .D(n144), .Y(n198) );
  AOI22X1 U210 ( .A(\In<14> ), .B(n218), .C(\In<13> ), .D(n134), .Y(n201) );
  AOI22X1 U211 ( .A(\In<12> ), .B(n220), .C(\In<11> ), .D(n219), .Y(n200) );
  AOI22X1 U212 ( .A(\In<6> ), .B(n218), .C(\In<5> ), .D(n134), .Y(n203) );
  AOI22X1 U213 ( .A(\In<4> ), .B(n220), .C(\In<3> ), .D(n219), .Y(n202) );
  AOI22X1 U214 ( .A(n103), .B(n145), .C(n8), .D(n163), .Y(n211) );
  AOI22X1 U215 ( .A(\In<10> ), .B(n218), .C(\In<9> ), .D(n134), .Y(n205) );
  AOI22X1 U216 ( .A(\In<8> ), .B(n220), .C(\In<7> ), .D(n219), .Y(n204) );
  AOI22X1 U217 ( .A(\In<1> ), .B(n134), .C(\Cnt<1> ), .D(n206), .Y(n207) );
  OAI21X1 U218 ( .A(n209), .B(n208), .C(n56), .Y(n242) );
  AOI22X1 U219 ( .A(n9), .B(n155), .C(n246), .D(n242), .Y(n210) );
  AOI22X1 U220 ( .A(\In<15> ), .B(n218), .C(\In<14> ), .D(n134), .Y(n213) );
  AOI22X1 U221 ( .A(\In<13> ), .B(n220), .C(\In<12> ), .D(n219), .Y(n212) );
  AOI22X1 U222 ( .A(\In<7> ), .B(n218), .C(\In<6> ), .D(n134), .Y(n215) );
  AOI22X1 U223 ( .A(\In<5> ), .B(n220), .C(\In<4> ), .D(n219), .Y(n214) );
  AOI22X1 U224 ( .A(n103), .B(n149), .C(n87), .D(n8), .Y(n224) );
  AOI22X1 U225 ( .A(\In<11> ), .B(n218), .C(\In<10> ), .D(n134), .Y(n217) );
  AOI22X1 U226 ( .A(\In<9> ), .B(n220), .C(\In<8> ), .D(n219), .Y(n216) );
  AOI22X1 U227 ( .A(\In<3> ), .B(n218), .C(\In<2> ), .D(n134), .Y(n222) );
  AOI22X1 U228 ( .A(\In<1> ), .B(n220), .C(\In<0> ), .D(n219), .Y(n221) );
  AOI22X1 U229 ( .A(n9), .B(n158), .C(n246), .D(n167), .Y(n223) );
  AOI22X1 U230 ( .A(n152), .B(n9), .C(n160), .D(n246), .Y(n225) );
  NAND3X1 U231 ( .A(n20), .B(n22), .C(n92), .Y(\Out<4> ) );
  AOI22X1 U232 ( .A(n9), .B(n140), .C(n246), .D(n114), .Y(n226) );
  NAND3X1 U233 ( .A(n125), .B(n91), .C(n133), .Y(\Out<5> ) );
  AOI22X1 U234 ( .A(n245), .B(n242), .C(n8), .D(n156), .Y(n228) );
  AOI22X1 U235 ( .A(n9), .B(n146), .C(n246), .D(n164), .Y(n227) );
  AOI22X1 U236 ( .A(n245), .B(n166), .C(n8), .D(n157), .Y(n230) );
  AOI22X1 U237 ( .A(n9), .B(n148), .C(n246), .D(n135), .Y(n229) );
  AOI22X1 U238 ( .A(n8), .B(n153), .C(n99), .D(n1), .Y(n232) );
  AOI22X1 U239 ( .A(n246), .B(n138), .C(n160), .D(n245), .Y(n231) );
  AOI22X1 U240 ( .A(n246), .B(n144), .C(n245), .D(n114), .Y(n233) );
  NAND3X1 U241 ( .A(n83), .B(n131), .C(n120), .Y(\Out<9> ) );
  AOI22X1 U242 ( .A(n8), .B(n145), .C(n1), .D(n242), .Y(n235) );
  AOI22X1 U243 ( .A(n246), .B(n155), .C(n245), .D(n164), .Y(n234) );
  AOI22X1 U244 ( .A(n8), .B(n150), .C(n1), .D(n166), .Y(n237) );
  AOI22X1 U245 ( .A(n246), .B(n157), .C(n245), .D(n135), .Y(n236) );
  AOI22X1 U246 ( .A(n161), .B(n1), .C(n115), .D(n100), .Y(n239) );
  AOI22X1 U247 ( .A(n152), .B(n246), .C(n245), .D(n137), .Y(n238) );
  AOI22X1 U248 ( .A(n246), .B(n141), .C(n245), .D(n144), .Y(n241) );
  NAND3X1 U249 ( .A(n85), .B(n34), .C(n93), .Y(\Out<13> ) );
  AOI22X1 U250 ( .A(n1), .B(n163), .C(n115), .D(n242), .Y(n244) );
  AOI22X1 U251 ( .A(n246), .B(n146), .C(n245), .D(n156), .Y(n243) );
  AOI22X1 U252 ( .A(n1), .B(n87), .C(n115), .D(n167), .Y(n248) );
  AOI22X1 U253 ( .A(n246), .B(n148), .C(n245), .D(n157), .Y(n247) );
endmodule


module rshifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), Rot_sel, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , Rot_sel;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n33,
         n35, n36, n38, n39, n40, n41, n42, n43, n44, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254;

  INVX1 U2 ( .A(\Cnt<2> ), .Y(n190) );
  INVX1 U3 ( .A(\In<1> ), .Y(n210) );
  INVX1 U4 ( .A(\Cnt<1> ), .Y(n220) );
  INVX1 U5 ( .A(Rot_sel), .Y(n184) );
  INVX1 U6 ( .A(\In<13> ), .Y(n203) );
  AND2X1 U7 ( .A(n125), .B(n111), .Y(n31) );
  INVX4 U8 ( .A(n212), .Y(n227) );
  AND2X2 U9 ( .A(\Cnt<3> ), .B(n190), .Y(n1) );
  INVX1 U10 ( .A(n1), .Y(n2) );
  AND2X2 U11 ( .A(\Cnt<0> ), .B(\Cnt<1> ), .Y(n3) );
  AND2X2 U12 ( .A(n70), .B(n57), .Y(n4) );
  AND2X2 U13 ( .A(n71), .B(n58), .Y(n5) );
  AND2X2 U14 ( .A(n73), .B(n109), .Y(n6) );
  INVX1 U15 ( .A(n6), .Y(n7) );
  AND2X2 U16 ( .A(n74), .B(n59), .Y(n8) );
  AND2X2 U17 ( .A(n72), .B(n60), .Y(n9) );
  INVX1 U18 ( .A(n9), .Y(\Out<0> ) );
  AND2X2 U19 ( .A(n75), .B(n61), .Y(n11) );
  AND2X2 U20 ( .A(n76), .B(n62), .Y(n12) );
  AND2X2 U21 ( .A(\In<15> ), .B(n226), .Y(n13) );
  AND2X2 U22 ( .A(n183), .B(n211), .Y(n14) );
  AND2X2 U23 ( .A(n77), .B(n63), .Y(n15) );
  AND2X2 U24 ( .A(n78), .B(n64), .Y(n16) );
  AND2X2 U25 ( .A(n220), .B(n219), .Y(n17) );
  INVX1 U26 ( .A(n17), .Y(n18) );
  AND2X2 U27 ( .A(n79), .B(n65), .Y(n19) );
  AND2X2 U28 ( .A(n104), .B(n159), .Y(n20) );
  INVX1 U29 ( .A(n20), .Y(n21) );
  AND2X2 U30 ( .A(n80), .B(n66), .Y(n22) );
  AND2X2 U31 ( .A(n81), .B(n67), .Y(n23) );
  AND2X2 U32 ( .A(n183), .B(n103), .Y(n24) );
  AND2X2 U33 ( .A(n166), .B(n24), .Y(n25) );
  INVX1 U34 ( .A(n25), .Y(n26) );
  AND2X2 U35 ( .A(n164), .B(n244), .Y(n27) );
  INVX1 U36 ( .A(n27), .Y(n28) );
  AND2X2 U37 ( .A(n82), .B(n68), .Y(n29) );
  INVX1 U38 ( .A(n29), .Y(\Out<5> ) );
  INVX1 U39 ( .A(n31), .Y(\Out<6> ) );
  AND2X2 U40 ( .A(n127), .B(n69), .Y(n33) );
  INVX1 U41 ( .A(n33), .Y(\Out<7> ) );
  AND2X2 U42 ( .A(n183), .B(n1), .Y(n35) );
  AND2X2 U43 ( .A(n83), .B(n113), .Y(n36) );
  INVX1 U44 ( .A(n36), .Y(\Out<8> ) );
  AND2X2 U45 ( .A(n163), .B(n35), .Y(n38) );
  INVX1 U46 ( .A(n38), .Y(n39) );
  AND2X2 U47 ( .A(n160), .B(n24), .Y(n40) );
  INVX1 U48 ( .A(n40), .Y(n41) );
  AND2X2 U49 ( .A(n253), .B(n158), .Y(n42) );
  INVX1 U50 ( .A(n42), .Y(n43) );
  AND2X2 U51 ( .A(n84), .B(n100), .Y(n44) );
  INVX1 U52 ( .A(n44), .Y(\Out<12> ) );
  AND2X2 U53 ( .A(n253), .B(n252), .Y(n46) );
  INVX1 U54 ( .A(n46), .Y(n47) );
  BUFX2 U55 ( .A(n200), .Y(n48) );
  BUFX2 U56 ( .A(n209), .Y(n49) );
  BUFX2 U57 ( .A(n199), .Y(n50) );
  BUFX2 U58 ( .A(n208), .Y(n51) );
  OR2X2 U59 ( .A(n102), .B(n120), .Y(n52) );
  INVX1 U60 ( .A(n52), .Y(n53) );
  BUFX2 U61 ( .A(n202), .Y(n54) );
  AND2X2 U62 ( .A(\In<0> ), .B(n228), .Y(n55) );
  INVX1 U63 ( .A(n55), .Y(n56) );
  BUFX2 U64 ( .A(n186), .Y(n57) );
  BUFX2 U65 ( .A(n188), .Y(n58) );
  BUFX2 U66 ( .A(n195), .Y(n59) );
  BUFX2 U67 ( .A(n197), .Y(n60) );
  BUFX2 U68 ( .A(n204), .Y(n61) );
  BUFX2 U69 ( .A(n206), .Y(n62) );
  BUFX2 U70 ( .A(n213), .Y(n63) );
  BUFX2 U71 ( .A(n215), .Y(n64) );
  BUFX2 U72 ( .A(n222), .Y(n65) );
  BUFX2 U73 ( .A(n224), .Y(n66) );
  BUFX2 U74 ( .A(n229), .Y(n67) );
  BUFX2 U75 ( .A(n233), .Y(n68) );
  BUFX2 U76 ( .A(n237), .Y(n69) );
  BUFX2 U77 ( .A(n187), .Y(n70) );
  BUFX2 U78 ( .A(n189), .Y(n71) );
  BUFX2 U79 ( .A(n198), .Y(n72) );
  BUFX2 U80 ( .A(n193), .Y(n73) );
  BUFX2 U81 ( .A(n196), .Y(n74) );
  BUFX2 U82 ( .A(n205), .Y(n75) );
  BUFX2 U83 ( .A(n207), .Y(n76) );
  BUFX2 U84 ( .A(n214), .Y(n77) );
  BUFX2 U85 ( .A(n216), .Y(n78) );
  BUFX2 U86 ( .A(n223), .Y(n79) );
  BUFX2 U87 ( .A(n225), .Y(n80) );
  BUFX2 U88 ( .A(n230), .Y(n81) );
  BUFX2 U89 ( .A(n234), .Y(n82) );
  BUFX2 U90 ( .A(n240), .Y(n83) );
  BUFX2 U91 ( .A(n246), .Y(n84) );
  BUFX2 U92 ( .A(n254), .Y(n85) );
  AND2X2 U93 ( .A(n103), .B(n250), .Y(n86) );
  INVX1 U94 ( .A(n86), .Y(n87) );
  AND2X2 U95 ( .A(n103), .B(n252), .Y(n88) );
  INVX1 U96 ( .A(n88), .Y(n89) );
  BUFX2 U97 ( .A(n221), .Y(n90) );
  AND2X2 U98 ( .A(n244), .B(n252), .Y(n91) );
  INVX1 U99 ( .A(n91), .Y(n92) );
  BUFX2 U100 ( .A(n232), .Y(n93) );
  BUFX2 U101 ( .A(n241), .Y(n94) );
  BUFX2 U102 ( .A(n249), .Y(n95) );
  AND2X1 U103 ( .A(\Cnt<0> ), .B(n220), .Y(n96) );
  INVX1 U104 ( .A(n96), .Y(n97) );
  AND2X2 U105 ( .A(n49), .B(n51), .Y(n138) );
  AND2X2 U106 ( .A(n183), .B(n244), .Y(n98) );
  INVX1 U107 ( .A(n245), .Y(n99) );
  INVX1 U108 ( .A(n99), .Y(n100) );
  OR2X2 U109 ( .A(n212), .B(n121), .Y(n101) );
  INVX1 U110 ( .A(n101), .Y(n102) );
  AND2X2 U111 ( .A(\Cnt<3> ), .B(\Cnt<2> ), .Y(n103) );
  INVX1 U112 ( .A(n2), .Y(n104) );
  INVX1 U113 ( .A(n2), .Y(n105) );
  INVX1 U114 ( .A(\In<15> ), .Y(n201) );
  INVX1 U115 ( .A(n217), .Y(n106) );
  INVX1 U116 ( .A(n106), .Y(n107) );
  INVX1 U117 ( .A(n192), .Y(n108) );
  INVX1 U118 ( .A(n108), .Y(n109) );
  INVX1 U119 ( .A(n235), .Y(n110) );
  INVX1 U120 ( .A(n110), .Y(n111) );
  INVX1 U121 ( .A(n239), .Y(n112) );
  INVX1 U122 ( .A(n112), .Y(n113) );
  AND2X2 U123 ( .A(n244), .B(n250), .Y(n114) );
  INVX1 U124 ( .A(n114), .Y(n115) );
  AND2X2 U125 ( .A(n253), .B(n250), .Y(n116) );
  INVX1 U126 ( .A(n116), .Y(n117) );
  AND2X2 U127 ( .A(\In<14> ), .B(n227), .Y(n118) );
  OR2X2 U128 ( .A(n122), .B(n123), .Y(n119) );
  INVX1 U129 ( .A(n119), .Y(n120) );
  INVX1 U130 ( .A(\In<2> ), .Y(n121) );
  INVX1 U131 ( .A(n226), .Y(n122) );
  INVX1 U132 ( .A(\In<3> ), .Y(n123) );
  INVX4 U133 ( .A(n97), .Y(n226) );
  INVX2 U134 ( .A(n182), .Y(n247) );
  INVX1 U135 ( .A(n236), .Y(n124) );
  INVX1 U136 ( .A(n124), .Y(n125) );
  INVX1 U137 ( .A(n238), .Y(n126) );
  INVX1 U138 ( .A(n126), .Y(n127) );
  AND2X2 U139 ( .A(n253), .B(n156), .Y(n128) );
  INVX1 U140 ( .A(n128), .Y(n129) );
  AND2X2 U141 ( .A(n163), .B(n98), .Y(n130) );
  INVX1 U142 ( .A(n130), .Y(n131) );
  AND2X2 U143 ( .A(n157), .B(n24), .Y(n132) );
  INVX1 U144 ( .A(n132), .Y(n133) );
  AND2X2 U145 ( .A(n159), .B(n24), .Y(n134) );
  INVX1 U146 ( .A(n134), .Y(n135) );
  AND2X2 U147 ( .A(n183), .B(\In<0> ), .Y(n136) );
  INVX1 U148 ( .A(n136), .Y(n137) );
  INVX1 U149 ( .A(n138), .Y(\Out<1> ) );
  AND2X2 U150 ( .A(n104), .B(n156), .Y(n140) );
  INVX1 U151 ( .A(n140), .Y(n141) );
  AND2X2 U152 ( .A(n161), .B(n35), .Y(n142) );
  INVX1 U153 ( .A(n142), .Y(n143) );
  INVX1 U154 ( .A(n218), .Y(n144) );
  INVX1 U155 ( .A(n144), .Y(n145) );
  INVX1 U156 ( .A(n231), .Y(n146) );
  INVX1 U157 ( .A(n146), .Y(n147) );
  INVX1 U158 ( .A(n242), .Y(n148) );
  INVX1 U159 ( .A(n148), .Y(n149) );
  INVX1 U160 ( .A(n243), .Y(n150) );
  INVX1 U161 ( .A(n150), .Y(n151) );
  INVX1 U162 ( .A(n251), .Y(n152) );
  INVX1 U163 ( .A(n152), .Y(n153) );
  INVX2 U164 ( .A(n3), .Y(n154) );
  INVX8 U165 ( .A(n154), .Y(n155) );
  INVX1 U166 ( .A(n15), .Y(n156) );
  INVX1 U167 ( .A(n15), .Y(n157) );
  INVX1 U168 ( .A(n19), .Y(n158) );
  INVX1 U169 ( .A(n19), .Y(n159) );
  INVX1 U170 ( .A(n11), .Y(n160) );
  INVX1 U171 ( .A(n11), .Y(n161) );
  INVX1 U172 ( .A(n12), .Y(n162) );
  INVX1 U173 ( .A(n12), .Y(n163) );
  INVX1 U174 ( .A(n4), .Y(n164) );
  INVX1 U175 ( .A(n4), .Y(n165) );
  INVX1 U176 ( .A(n8), .Y(n166) );
  INVX1 U177 ( .A(n8), .Y(n167) );
  INVX1 U178 ( .A(n16), .Y(n168) );
  INVX1 U179 ( .A(n16), .Y(n169) );
  INVX1 U180 ( .A(n22), .Y(n170) );
  INVX1 U181 ( .A(n22), .Y(n171) );
  INVX1 U182 ( .A(n5), .Y(n172) );
  INVX1 U183 ( .A(n5), .Y(n173) );
  INVX1 U184 ( .A(n176), .Y(n174) );
  INVX1 U185 ( .A(n176), .Y(n175) );
  AND2X2 U186 ( .A(n107), .B(n53), .Y(n176) );
  INVX1 U187 ( .A(n23), .Y(n177) );
  INVX1 U188 ( .A(n23), .Y(n178) );
  NOR3X1 U189 ( .A(n118), .B(n14), .C(n13), .Y(n179) );
  INVX1 U190 ( .A(n179), .Y(n250) );
  INVX1 U191 ( .A(n248), .Y(n180) );
  INVX1 U192 ( .A(n180), .Y(n181) );
  AND2X2 U193 ( .A(n48), .B(n50), .Y(n182) );
  INVX8 U194 ( .A(n185), .Y(n228) );
  INVX4 U195 ( .A(n191), .Y(n244) );
  INVX8 U196 ( .A(n194), .Y(n253) );
  INVX8 U197 ( .A(n184), .Y(n183) );
  OR2X2 U198 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n212) );
  AOI22X1 U199 ( .A(\In<8> ), .B(n227), .C(\In<9> ), .D(n226), .Y(n187) );
  OR2X2 U200 ( .A(n220), .B(\Cnt<0> ), .Y(n185) );
  AOI22X1 U201 ( .A(\In<10> ), .B(n228), .C(\In<11> ), .D(n155), .Y(n186) );
  AOI22X1 U202 ( .A(\In<12> ), .B(n227), .C(\In<13> ), .D(n226), .Y(n189) );
  AOI22X1 U203 ( .A(\In<14> ), .B(n228), .C(\In<15> ), .D(n155), .Y(n188) );
  AOI22X1 U204 ( .A(n104), .B(n164), .C(n103), .D(n173), .Y(n198) );
  OR2X2 U205 ( .A(n190), .B(\Cnt<3> ), .Y(n191) );
  AOI22X1 U206 ( .A(\In<5> ), .B(n226), .C(\In<4> ), .D(n227), .Y(n193) );
  AOI22X1 U207 ( .A(\In<7> ), .B(n155), .C(\In<6> ), .D(n228), .Y(n192) );
  OR2X2 U208 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n194) );
  AOI22X1 U209 ( .A(\In<0> ), .B(n227), .C(\In<1> ), .D(n226), .Y(n196) );
  AOI22X1 U210 ( .A(\In<2> ), .B(n228), .C(\In<3> ), .D(n155), .Y(n195) );
  AOI22X1 U211 ( .A(n244), .B(n7), .C(n253), .D(n167), .Y(n197) );
  AOI22X1 U212 ( .A(\In<10> ), .B(n226), .C(\In<9> ), .D(n227), .Y(n200) );
  AOI22X1 U213 ( .A(\In<12> ), .B(n155), .C(\In<11> ), .D(n228), .Y(n199) );
  MUX2X1 U214 ( .B(n201), .A(n137), .S(\Cnt<0> ), .Y(n219) );
  AOI22X1 U215 ( .A(\In<14> ), .B(n226), .C(\Cnt<1> ), .D(n219), .Y(n202) );
  OAI21X1 U216 ( .A(n212), .B(n203), .C(n54), .Y(n248) );
  AOI22X1 U217 ( .A(n105), .B(n247), .C(n103), .D(n248), .Y(n209) );
  AOI22X1 U218 ( .A(\In<5> ), .B(n227), .C(\In<6> ), .D(n226), .Y(n205) );
  AOI22X1 U219 ( .A(\In<7> ), .B(n228), .C(\In<8> ), .D(n155), .Y(n204) );
  AOI22X1 U220 ( .A(\In<1> ), .B(n227), .C(\In<2> ), .D(n226), .Y(n207) );
  AOI22X1 U221 ( .A(\In<3> ), .B(n228), .C(\In<4> ), .D(n155), .Y(n206) );
  AOI22X1 U222 ( .A(n244), .B(n160), .C(n253), .D(n162), .Y(n208) );
  OAI21X1 U223 ( .A(n154), .B(n210), .C(n56), .Y(n211) );
  AOI22X1 U224 ( .A(\In<10> ), .B(n227), .C(\In<11> ), .D(n226), .Y(n214) );
  AOI22X1 U225 ( .A(\In<12> ), .B(n228), .C(\In<13> ), .D(n155), .Y(n213) );
  AOI22X1 U226 ( .A(\In<6> ), .B(n227), .C(\In<7> ), .D(n226), .Y(n216) );
  AOI22X1 U227 ( .A(\In<8> ), .B(n228), .C(\In<9> ), .D(n155), .Y(n215) );
  AOI22X1 U228 ( .A(\In<4> ), .B(n228), .C(\In<5> ), .D(n155), .Y(n217) );
  AOI22X1 U229 ( .A(n244), .B(n168), .C(n253), .D(n174), .Y(n218) );
  NAND3X1 U230 ( .A(n87), .B(n141), .C(n145), .Y(\Out<2> ) );
  AOI22X1 U231 ( .A(\In<1> ), .B(n228), .C(\In<2> ), .D(n155), .Y(n221) );
  OAI21X1 U232 ( .A(n90), .B(n184), .C(n18), .Y(n252) );
  AOI22X1 U233 ( .A(\In<11> ), .B(n227), .C(\In<12> ), .D(n226), .Y(n223) );
  AOI22X1 U234 ( .A(\In<13> ), .B(n228), .C(\In<14> ), .D(n155), .Y(n222) );
  AOI22X1 U235 ( .A(\In<7> ), .B(n227), .C(\In<8> ), .D(n226), .Y(n225) );
  AOI22X1 U236 ( .A(\In<9> ), .B(n228), .C(\In<10> ), .D(n155), .Y(n224) );
  AOI22X1 U237 ( .A(\In<3> ), .B(n227), .C(\In<4> ), .D(n226), .Y(n230) );
  AOI22X1 U238 ( .A(\In<5> ), .B(n228), .C(\In<6> ), .D(n155), .Y(n229) );
  AOI22X1 U239 ( .A(n244), .B(n171), .C(n253), .D(n178), .Y(n231) );
  NAND3X1 U240 ( .A(n89), .B(n21), .C(n147), .Y(\Out<3> ) );
  AOI22X1 U241 ( .A(n253), .B(n7), .C(n172), .D(n105), .Y(n232) );
  NAND3X1 U242 ( .A(n26), .B(n28), .C(n93), .Y(\Out<4> ) );
  AOI22X1 U243 ( .A(n244), .B(n247), .C(n162), .D(n24), .Y(n234) );
  AOI22X1 U244 ( .A(n253), .B(n161), .C(n104), .D(n181), .Y(n233) );
  AOI22X1 U245 ( .A(n244), .B(n157), .C(n175), .D(n24), .Y(n236) );
  AOI22X1 U246 ( .A(n253), .B(n169), .C(n105), .D(n250), .Y(n235) );
  AOI22X1 U247 ( .A(n244), .B(n158), .C(n177), .D(n24), .Y(n238) );
  AOI22X1 U248 ( .A(n253), .B(n170), .C(n105), .D(n252), .Y(n237) );
  AOI22X1 U249 ( .A(n7), .B(n24), .C(n167), .D(n35), .Y(n240) );
  AOI22X1 U250 ( .A(n172), .B(n244), .C(n165), .D(n253), .Y(n239) );
  AOI22X1 U251 ( .A(n244), .B(n248), .C(n253), .D(n247), .Y(n241) );
  NAND3X1 U252 ( .A(n39), .B(n41), .C(n94), .Y(\Out<9> ) );
  AOI22X1 U253 ( .A(n168), .B(n24), .C(n174), .D(n35), .Y(n242) );
  NAND3X1 U254 ( .A(n129), .B(n115), .C(n149), .Y(\Out<10> ) );
  AOI22X1 U255 ( .A(n171), .B(n24), .C(n177), .D(n35), .Y(n243) );
  NAND3X1 U256 ( .A(n43), .B(n92), .C(n151), .Y(\Out<11> ) );
  AOI22X1 U257 ( .A(n7), .B(n35), .C(n167), .D(n98), .Y(n246) );
  AOI22X1 U258 ( .A(n173), .B(n253), .C(n165), .D(n24), .Y(n245) );
  AOI22X1 U259 ( .A(n253), .B(n181), .C(n247), .D(n24), .Y(n249) );
  NAND3X1 U260 ( .A(n131), .B(n143), .C(n95), .Y(\Out<13> ) );
  AOI22X1 U261 ( .A(n169), .B(n35), .C(n175), .D(n98), .Y(n251) );
  NAND3X1 U262 ( .A(n133), .B(n117), .C(n153), .Y(\Out<14> ) );
  AOI22X1 U263 ( .A(n170), .B(n35), .C(n178), .D(n98), .Y(n254) );
  NAND3X1 U264 ( .A(n85), .B(n47), .C(n135), .Y(\Out<15> ) );
endmodule


module fulladder1_31 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  INVX1 U2 ( .A(Cin), .Y(n2) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(P) );
  XNOR2X1 U5 ( .A(P), .B(n2), .Y(S) );
endmodule


module fulladder1_30 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_29 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_28 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_27 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_26 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_25 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_24 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_23 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_22 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_21 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_20 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_19 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_18 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_17 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX1 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_16 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module cla4_11 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  fulladder1_44 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n45), .G(n41) );
  fulladder1_45 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n14), .S(\S<1> ), .P(
        n46), .G(n42) );
  fulladder1_46 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n40), .S(\S<2> ), .P(
        n47), .G(n43) );
  fulladder1_47 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n39), .S(\S<3> ), .P(
        n48), .G(n44) );
  INVX1 U1 ( .A(n22), .Y(n34) );
  INVX1 U2 ( .A(n39), .Y(n38) );
  AND2X2 U3 ( .A(n46), .B(n24), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X2 U5 ( .A(n47), .B(n25), .Y(n3) );
  AND2X2 U6 ( .A(n34), .B(n11), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n5) );
  OR2X2 U8 ( .A(n5), .B(n9), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(PG) );
  BUFX2 U10 ( .A(n23), .Y(n8) );
  BUFX2 U11 ( .A(n36), .Y(n9) );
  BUFX2 U12 ( .A(n33), .Y(n10) );
  AND2X2 U13 ( .A(n48), .B(n32), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(n12) );
  AND2X2 U15 ( .A(n8), .B(n19), .Y(n13) );
  INVX1 U16 ( .A(n13), .Y(n14) );
  BUFX2 U17 ( .A(n27), .Y(n15) );
  BUFX2 U18 ( .A(n37), .Y(n16) );
  INVX1 U19 ( .A(n30), .Y(n17) );
  INVX1 U20 ( .A(n29), .Y(n30) );
  INVX1 U21 ( .A(n28), .Y(n18) );
  INVX1 U22 ( .A(n18), .Y(n19) );
  INVX1 U23 ( .A(n3), .Y(n20) );
  INVX1 U24 ( .A(n35), .Y(n21) );
  INVX1 U25 ( .A(n2), .Y(n35) );
  XNOR2X1 U26 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  NAND3X1 U27 ( .A(Cin), .B(n45), .C(n34), .Y(n23) );
  NAND3X1 U28 ( .A(\A<0> ), .B(\B<0> ), .C(n41), .Y(n28) );
  XOR2X1 U29 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  NAND3X1 U30 ( .A(\A<1> ), .B(\B<1> ), .C(n42), .Y(n27) );
  OAI21X1 U31 ( .A(n21), .B(n13), .C(n15), .Y(n40) );
  XOR2X1 U32 ( .A(\A<2> ), .B(\B<2> ), .Y(n25) );
  INVX2 U33 ( .A(n40), .Y(n26) );
  NAND3X1 U34 ( .A(\A<2> ), .B(\B<2> ), .C(n43), .Y(n29) );
  OAI21X1 U35 ( .A(n20), .B(n26), .C(n17), .Y(n39) );
  OAI21X1 U36 ( .A(n2), .B(n19), .C(n15), .Y(n31) );
  AOI21X1 U37 ( .A(n3), .B(n31), .C(n30), .Y(n33) );
  XOR2X1 U38 ( .A(\A<3> ), .B(\B<3> ), .Y(n32) );
  NAND3X1 U39 ( .A(\A<3> ), .B(\B<3> ), .C(n44), .Y(n37) );
  OAI21X1 U40 ( .A(n10), .B(n12), .C(n16), .Y(GG) );
  NAND3X1 U41 ( .A(n45), .B(n35), .C(n3), .Y(n36) );
  OAI21X1 U42 ( .A(n12), .B(n38), .C(n16), .Y(Cout) );
endmodule


module cla4_10 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  fulladder1_43 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n45), .G(n41) );
  fulladder1_42 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n20), .S(\S<1> ), .P(
        n46), .G(n42) );
  fulladder1_41 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n40), .S(\S<2> ), .P(
        n47), .G(n43) );
  fulladder1_40 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n39), .S(\S<3> ), .P(
        n48), .G(n44) );
  INVX1 U1 ( .A(n22), .Y(n34) );
  INVX1 U2 ( .A(n39), .Y(n38) );
  AND2X2 U3 ( .A(n46), .B(n24), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X2 U5 ( .A(n47), .B(n25), .Y(n3) );
  AND2X2 U6 ( .A(n34), .B(n11), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n5) );
  OR2X2 U8 ( .A(n5), .B(n9), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(PG) );
  BUFX2 U10 ( .A(n23), .Y(n8) );
  BUFX2 U11 ( .A(n36), .Y(n9) );
  BUFX2 U12 ( .A(n33), .Y(n10) );
  AND2X2 U13 ( .A(n48), .B(n32), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(n12) );
  BUFX2 U15 ( .A(n27), .Y(n13) );
  BUFX2 U16 ( .A(n37), .Y(n14) );
  INVX1 U17 ( .A(n30), .Y(n15) );
  INVX1 U18 ( .A(n29), .Y(n30) );
  INVX1 U19 ( .A(n28), .Y(n16) );
  INVX1 U20 ( .A(n16), .Y(n17) );
  INVX1 U21 ( .A(n3), .Y(n18) );
  AND2X2 U22 ( .A(n8), .B(n17), .Y(n19) );
  INVX1 U23 ( .A(n19), .Y(n20) );
  INVX1 U24 ( .A(n35), .Y(n21) );
  INVX1 U25 ( .A(n2), .Y(n35) );
  XNOR2X1 U26 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  NAND3X1 U27 ( .A(n45), .B(n34), .C(Cin), .Y(n23) );
  NAND3X1 U28 ( .A(\A<0> ), .B(\B<0> ), .C(n41), .Y(n28) );
  XOR2X1 U29 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  NAND3X1 U30 ( .A(\A<1> ), .B(\B<1> ), .C(n42), .Y(n27) );
  OAI21X1 U31 ( .A(n21), .B(n19), .C(n13), .Y(n40) );
  XOR2X1 U32 ( .A(\A<2> ), .B(\B<2> ), .Y(n25) );
  INVX2 U33 ( .A(n40), .Y(n26) );
  NAND3X1 U34 ( .A(\A<2> ), .B(\B<2> ), .C(n43), .Y(n29) );
  OAI21X1 U35 ( .A(n18), .B(n26), .C(n15), .Y(n39) );
  OAI21X1 U36 ( .A(n2), .B(n17), .C(n13), .Y(n31) );
  AOI21X1 U37 ( .A(n3), .B(n31), .C(n30), .Y(n33) );
  XOR2X1 U38 ( .A(\A<3> ), .B(\B<3> ), .Y(n32) );
  NAND3X1 U39 ( .A(\A<3> ), .B(\B<3> ), .C(n44), .Y(n37) );
  OAI21X1 U40 ( .A(n10), .B(n12), .C(n14), .Y(GG) );
  NAND3X1 U41 ( .A(n45), .B(n35), .C(n3), .Y(n36) );
  OAI21X1 U42 ( .A(n12), .B(n38), .C(n14), .Y(Cout) );
endmodule


module cla4_9 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \G<3> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48;

  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n41) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n46) );
  OAI21X1 U10 ( .A(n4), .B(n37), .C(n36), .Y(GG) );
  fulladder1_39 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n43), .G(n38) );
  fulladder1_38 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n20), .S(\S<1> ), .P(
        n44), .G(n39) );
  fulladder1_37 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n22), .S(\S<2> ), .P(
        n45), .G(n40) );
  fulladder1_36 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n35), .S(\S<3> ), .P(
        n47), .G(n42) );
  INVX1 U1 ( .A(n17), .Y(n34) );
  AND2X1 U2 ( .A(n45), .B(n26), .Y(n16) );
  INVX1 U3 ( .A(\G<3> ), .Y(n36) );
  INVX1 U4 ( .A(\P<3> ), .Y(n37) );
  BUFX2 U5 ( .A(n24), .Y(n1) );
  AND2X2 U6 ( .A(n21), .B(n5), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  BUFX2 U8 ( .A(n48), .Y(n4) );
  AND2X2 U9 ( .A(n44), .B(n25), .Y(n5) );
  INVX1 U11 ( .A(n5), .Y(n6) );
  BUFX2 U12 ( .A(n28), .Y(n7) );
  AND2X2 U13 ( .A(n12), .B(n3), .Y(n8) );
  AND2X2 U14 ( .A(\P<3> ), .B(n35), .Y(n9) );
  INVX1 U15 ( .A(n9), .Y(n10) );
  BUFX2 U16 ( .A(n29), .Y(n12) );
  INVX1 U17 ( .A(n30), .Y(n13) );
  INVX1 U18 ( .A(n13), .Y(n14) );
  INVX1 U19 ( .A(n32), .Y(n15) );
  INVX1 U20 ( .A(n31), .Y(n32) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  INVX1 U22 ( .A(n16), .Y(n18) );
  AND2X2 U23 ( .A(n14), .B(n1), .Y(n19) );
  INVX1 U24 ( .A(n19), .Y(n20) );
  INVX1 U25 ( .A(n19), .Y(n21) );
  INVX1 U26 ( .A(n8), .Y(n22) );
  NAND3X1 U27 ( .A(\A<0> ), .B(\B<0> ), .C(n38), .Y(n30) );
  XNOR2X1 U28 ( .A(\A<0> ), .B(\B<0> ), .Y(n27) );
  INVX2 U29 ( .A(n27), .Y(n23) );
  NAND3X1 U30 ( .A(n43), .B(n23), .C(Cin), .Y(n24) );
  NAND3X1 U31 ( .A(\A<1> ), .B(\B<1> ), .C(n39), .Y(n29) );
  XOR2X1 U32 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  XOR2X1 U33 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  NAND3X1 U34 ( .A(\A<2> ), .B(\B<2> ), .C(n40), .Y(n31) );
  OAI21X1 U35 ( .A(n18), .B(n8), .C(n15), .Y(n35) );
  NAND3X1 U36 ( .A(n43), .B(n5), .C(n34), .Y(n28) );
  NOR3X1 U37 ( .A(n7), .B(n27), .C(n37), .Y(PG) );
  NAND2X1 U38 ( .A(n36), .B(n10), .Y(Cout) );
  OAI21X1 U39 ( .A(n14), .B(n6), .C(n12), .Y(n33) );
  AOI21X1 U40 ( .A(n34), .B(n33), .C(n32), .Y(n48) );
  AND2X1 U41 ( .A(n46), .B(n47), .Y(\P<3> ) );
  AND2X1 U42 ( .A(n41), .B(n42), .Y(\G<3> ) );
endmodule


module cla4_8 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \G<3> , \G<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53;

  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n50) );
  NOR3X1 U8 ( .A(n16), .B(n27), .C(n41), .Y(PG) );
  OAI21X1 U10 ( .A(n14), .B(n41), .C(n40), .Y(GG) );
  AOI21X1 U11 ( .A(n26), .B(n39), .C(n22), .Y(n53) );
  AOI21X1 U12 ( .A(n24), .B(\G<0> ), .C(n19), .Y(n52) );
  fulladder1_35 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n47), .G(n42) );
  fulladder1_34 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n9), .S(\S<1> ), .P(n48), .G(n43) );
  fulladder1_33 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n38), .S(\S<2> ), .P(
        n49), .G(n44) );
  fulladder1_32 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n6), .S(\S<3> ), .P(n51), .G(n46) );
  INVX1 U1 ( .A(n10), .Y(n31) );
  INVX1 U2 ( .A(n49), .Y(n32) );
  INVX1 U3 ( .A(n21), .Y(\G<0> ) );
  INVX1 U4 ( .A(\G<3> ), .Y(n40) );
  AND2X1 U5 ( .A(\A<3> ), .B(\B<3> ), .Y(n45) );
  INVX1 U6 ( .A(\P<3> ), .Y(n41) );
  AND2X2 U7 ( .A(Cin), .B(n18), .Y(n1) );
  INVX1 U9 ( .A(n1), .Y(n2) );
  AND2X2 U13 ( .A(n38), .B(n26), .Y(n3) );
  INVX1 U14 ( .A(n3), .Y(n4) );
  AND2X2 U15 ( .A(n23), .B(n4), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(n6) );
  INVX1 U17 ( .A(n5), .Y(n7) );
  AND2X2 U18 ( .A(n21), .B(n2), .Y(n8) );
  INVX1 U19 ( .A(n8), .Y(n9) );
  INVX1 U20 ( .A(n8), .Y(n10) );
  BUFX2 U21 ( .A(n52), .Y(n12) );
  INVX1 U22 ( .A(n12), .Y(n39) );
  BUFX2 U23 ( .A(n53), .Y(n14) );
  AND2X1 U24 ( .A(n24), .B(n18), .Y(n15) );
  INVX1 U25 ( .A(n15), .Y(n16) );
  OR2X2 U26 ( .A(n29), .B(n28), .Y(n17) );
  INVX1 U27 ( .A(n17), .Y(n18) );
  INVX1 U28 ( .A(n20), .Y(n19) );
  BUFX2 U29 ( .A(n36), .Y(n20) );
  BUFX2 U30 ( .A(n35), .Y(n21) );
  INVX1 U31 ( .A(n23), .Y(n22) );
  BUFX2 U32 ( .A(n37), .Y(n23) );
  AND2X1 U33 ( .A(n48), .B(n30), .Y(n24) );
  INVX1 U34 ( .A(n24), .Y(n25) );
  INVX1 U35 ( .A(n7), .Y(n34) );
  INVX1 U36 ( .A(n27), .Y(n26) );
  OR2X1 U37 ( .A(n33), .B(n32), .Y(n27) );
  NAND3X1 U38 ( .A(\A<0> ), .B(\B<0> ), .C(n42), .Y(n35) );
  XNOR2X1 U39 ( .A(\A<0> ), .B(\B<0> ), .Y(n29) );
  INVX2 U40 ( .A(n47), .Y(n28) );
  XOR2X1 U41 ( .A(\A<1> ), .B(\B<1> ), .Y(n30) );
  NAND3X1 U42 ( .A(\A<1> ), .B(\B<1> ), .C(n43), .Y(n36) );
  OAI21X1 U43 ( .A(n25), .B(n31), .C(n20), .Y(n38) );
  NAND3X1 U44 ( .A(\A<2> ), .B(\B<2> ), .C(n44), .Y(n37) );
  XNOR2X1 U45 ( .A(\A<2> ), .B(\B<2> ), .Y(n33) );
  OAI21X1 U46 ( .A(n34), .B(n41), .C(n40), .Y(Cout) );
  AND2X1 U47 ( .A(n50), .B(n51), .Y(\P<3> ) );
  AND2X1 U48 ( .A(n45), .B(n46), .Y(\G<3> ) );
endmodule


module register16_0 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_15 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_14 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(n3) );
  dff_13 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(rst) );
  dff_12 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_11 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_10 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_9 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_8 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_7 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_6 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_5 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_4 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_3 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_2 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_1 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_0 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\d<12> ), .Y(n11) );
  INVX1 U2 ( .A(\q<0> ), .Y(n42) );
  INVX1 U3 ( .A(\q<1> ), .Y(n39) );
  INVX1 U4 ( .A(\q<2> ), .Y(n36) );
  INVX1 U5 ( .A(\q<3> ), .Y(n33) );
  INVX1 U6 ( .A(\q<4> ), .Y(n30) );
  INVX1 U7 ( .A(\q<5> ), .Y(n27) );
  INVX1 U8 ( .A(\q<6> ), .Y(n24) );
  INVX1 U9 ( .A(\q<7> ), .Y(n21) );
  INVX1 U10 ( .A(\q<8> ), .Y(n20) );
  INVX1 U11 ( .A(rst), .Y(n4) );
  INVX1 U12 ( .A(n4), .Y(n3) );
  INVX1 U13 ( .A(\d<11> ), .Y(n13) );
  INVX1 U14 ( .A(\d<9> ), .Y(n17) );
  INVX1 U15 ( .A(\d<10> ), .Y(n15) );
  INVX1 U16 ( .A(\d<15> ), .Y(n5) );
  INVX1 U17 ( .A(\d<13> ), .Y(n9) );
  INVX1 U18 ( .A(\d<14> ), .Y(n7) );
  INVX1 U19 ( .A(\d<8> ), .Y(n19) );
  OAI21X1 U20 ( .A(n43), .B(n2), .C(n44), .Y(n52) );
  INVX2 U21 ( .A(wr_en), .Y(n2) );
  INVX1 U22 ( .A(\d<1> ), .Y(n40) );
  INVX1 U23 ( .A(\d<0> ), .Y(n43) );
  INVX1 U24 ( .A(\d<5> ), .Y(n28) );
  INVX1 U25 ( .A(\d<6> ), .Y(n25) );
  INVX1 U26 ( .A(\d<3> ), .Y(n34) );
  INVX1 U27 ( .A(\d<4> ), .Y(n31) );
  INVX1 U28 ( .A(\d<7> ), .Y(n22) );
  INVX1 U29 ( .A(\d<2> ), .Y(n37) );
  INVX8 U30 ( .A(n2), .Y(n1) );
  INVX2 U31 ( .A(\q<15> ), .Y(n6) );
  MUX2X1 U32 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  INVX2 U33 ( .A(\q<14> ), .Y(n8) );
  MUX2X1 U34 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  INVX2 U35 ( .A(\q<13> ), .Y(n10) );
  MUX2X1 U36 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  INVX2 U37 ( .A(\q<12> ), .Y(n12) );
  MUX2X1 U38 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  INVX2 U39 ( .A(\q<11> ), .Y(n14) );
  MUX2X1 U40 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  INVX2 U41 ( .A(\q<10> ), .Y(n16) );
  MUX2X1 U42 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  INVX2 U43 ( .A(\q<9> ), .Y(n18) );
  MUX2X1 U44 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U45 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U46 ( .A(n1), .B(n21), .Y(n23) );
  AOI22X1 U47 ( .A(n23), .B(n2), .C(n23), .D(n22), .Y(n45) );
  OR2X2 U48 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U49 ( .A(n26), .B(n2), .C(n26), .D(n25), .Y(n46) );
  OR2X2 U50 ( .A(n1), .B(n27), .Y(n29) );
  AOI22X1 U51 ( .A(n29), .B(n2), .C(n29), .D(n28), .Y(n47) );
  OR2X2 U52 ( .A(n1), .B(n30), .Y(n32) );
  AOI22X1 U53 ( .A(n32), .B(n2), .C(n32), .D(n31), .Y(n48) );
  OR2X2 U54 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U55 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U56 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U57 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U58 ( .A(n1), .B(n39), .Y(n41) );
  AOI22X1 U59 ( .A(n41), .B(n2), .C(n41), .D(n40), .Y(n51) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_1 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_31 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_30 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(rst) );
  dff_29 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(n3) );
  dff_28 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_27 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_26 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_25 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_24 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_23 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_22 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_21 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_20 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_19 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_18 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_17 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_16 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<2> ), .Y(n36) );
  INVX1 U3 ( .A(\q<3> ), .Y(n33) );
  INVX1 U4 ( .A(\q<4> ), .Y(n30) );
  INVX1 U5 ( .A(\q<6> ), .Y(n24) );
  INVX1 U6 ( .A(\q<1> ), .Y(n39) );
  INVX1 U7 ( .A(\q<5> ), .Y(n27) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(rst), .Y(n4) );
  INVX1 U11 ( .A(n4), .Y(n3) );
  INVX1 U12 ( .A(\d<12> ), .Y(n11) );
  INVX1 U13 ( .A(\d<11> ), .Y(n13) );
  INVX1 U14 ( .A(\d<9> ), .Y(n17) );
  INVX1 U15 ( .A(\d<10> ), .Y(n15) );
  INVX1 U16 ( .A(\d<15> ), .Y(n5) );
  INVX1 U17 ( .A(\d<13> ), .Y(n9) );
  INVX1 U18 ( .A(\d<14> ), .Y(n7) );
  INVX1 U19 ( .A(\d<8> ), .Y(n19) );
  OAI21X1 U20 ( .A(n2), .B(n31), .C(n32), .Y(n48) );
  INVX1 U21 ( .A(\d<4> ), .Y(n31) );
  OAI21X1 U22 ( .A(n43), .B(n2), .C(n44), .Y(n52) );
  INVX2 U23 ( .A(wr_en), .Y(n2) );
  INVX1 U24 ( .A(\d<1> ), .Y(n40) );
  INVX1 U25 ( .A(\d<0> ), .Y(n43) );
  INVX1 U26 ( .A(\d<3> ), .Y(n34) );
  INVX1 U27 ( .A(\d<2> ), .Y(n37) );
  INVX1 U28 ( .A(\d<6> ), .Y(n25) );
  INVX1 U29 ( .A(\d<5> ), .Y(n28) );
  INVX1 U30 ( .A(\d<7> ), .Y(n22) );
  INVX8 U31 ( .A(n2), .Y(n1) );
  INVX2 U32 ( .A(\q<15> ), .Y(n6) );
  MUX2X1 U33 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  INVX2 U34 ( .A(\q<14> ), .Y(n8) );
  MUX2X1 U35 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  INVX2 U36 ( .A(\q<13> ), .Y(n10) );
  MUX2X1 U37 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  INVX2 U38 ( .A(\q<12> ), .Y(n12) );
  MUX2X1 U39 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  INVX2 U40 ( .A(\q<11> ), .Y(n14) );
  MUX2X1 U41 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  INVX2 U42 ( .A(\q<10> ), .Y(n16) );
  MUX2X1 U43 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  INVX2 U44 ( .A(\q<9> ), .Y(n18) );
  MUX2X1 U45 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U46 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U47 ( .A(n1), .B(n21), .Y(n23) );
  AOI22X1 U48 ( .A(n23), .B(n2), .C(n23), .D(n22), .Y(n45) );
  OR2X2 U49 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U50 ( .A(n26), .B(n2), .C(n26), .D(n25), .Y(n46) );
  OR2X2 U51 ( .A(n1), .B(n27), .Y(n29) );
  AOI22X1 U52 ( .A(n29), .B(n2), .C(n29), .D(n28), .Y(n47) );
  OR2X2 U53 ( .A(n1), .B(n30), .Y(n32) );
  OR2X2 U54 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U55 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U56 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U57 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U58 ( .A(n1), .B(n39), .Y(n41) );
  AOI22X1 U59 ( .A(n41), .B(n2), .C(n41), .D(n40), .Y(n51) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_2 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_47 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_46 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(n3) );
  dff_45 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(rst) );
  dff_44 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_43 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_42 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_41 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_40 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_39 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_38 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_37 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_36 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_35 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_34 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_33 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_32 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<1> ), .Y(n39) );
  INVX1 U3 ( .A(\q<2> ), .Y(n36) );
  INVX1 U4 ( .A(\q<3> ), .Y(n33) );
  INVX1 U5 ( .A(\q<4> ), .Y(n30) );
  INVX1 U6 ( .A(\q<6> ), .Y(n24) );
  INVX1 U7 ( .A(\q<5> ), .Y(n27) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(\q<9> ), .Y(n18) );
  INVX1 U11 ( .A(\q<10> ), .Y(n16) );
  INVX1 U12 ( .A(\q<11> ), .Y(n14) );
  INVX1 U13 ( .A(\q<12> ), .Y(n12) );
  INVX1 U14 ( .A(\q<14> ), .Y(n8) );
  INVX1 U15 ( .A(\q<15> ), .Y(n6) );
  INVX1 U16 ( .A(rst), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n3) );
  INVX1 U18 ( .A(\d<6> ), .Y(n25) );
  INVX1 U19 ( .A(\d<13> ), .Y(n9) );
  INVX1 U20 ( .A(\d<11> ), .Y(n13) );
  INVX1 U21 ( .A(\d<10> ), .Y(n15) );
  INVX1 U22 ( .A(\d<9> ), .Y(n17) );
  INVX1 U23 ( .A(\d<8> ), .Y(n19) );
  OAI21X1 U24 ( .A(n2), .B(n31), .C(n32), .Y(n48) );
  INVX1 U25 ( .A(\d<4> ), .Y(n31) );
  OAI21X1 U26 ( .A(n2), .B(n40), .C(n41), .Y(n51) );
  OAI21X1 U27 ( .A(n2), .B(n22), .C(n23), .Y(n45) );
  OAI21X1 U28 ( .A(n43), .B(n2), .C(n44), .Y(n52) );
  INVX2 U29 ( .A(wr_en), .Y(n2) );
  INVX1 U30 ( .A(\d<15> ), .Y(n5) );
  INVX1 U31 ( .A(\d<12> ), .Y(n11) );
  MUX2X1 U32 ( .B(n13), .A(n14), .S(n2), .Y(n56) );
  INVX1 U33 ( .A(\d<14> ), .Y(n7) );
  INVX1 U34 ( .A(\d<1> ), .Y(n40) );
  INVX1 U35 ( .A(\d<0> ), .Y(n43) );
  INVX1 U36 ( .A(\d<2> ), .Y(n37) );
  INVX1 U37 ( .A(\d<5> ), .Y(n28) );
  INVX1 U38 ( .A(\d<3> ), .Y(n34) );
  INVX1 U39 ( .A(\d<7> ), .Y(n22) );
  INVX8 U40 ( .A(n2), .Y(n1) );
  MUX2X1 U41 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  MUX2X1 U42 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  INVX2 U43 ( .A(\q<13> ), .Y(n10) );
  MUX2X1 U44 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  MUX2X1 U45 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  MUX2X1 U46 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  MUX2X1 U47 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U48 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U49 ( .A(n1), .B(n21), .Y(n23) );
  OR2X2 U50 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U51 ( .A(n26), .B(n2), .C(n25), .D(n26), .Y(n46) );
  OR2X2 U52 ( .A(n1), .B(n27), .Y(n29) );
  AOI22X1 U53 ( .A(n29), .B(n2), .C(n29), .D(n28), .Y(n47) );
  OR2X2 U54 ( .A(n1), .B(n30), .Y(n32) );
  OR2X2 U55 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U56 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U57 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U58 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U59 ( .A(n1), .B(n39), .Y(n41) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_3 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_63 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_62 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(rst) );
  dff_61 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(n3) );
  dff_60 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_59 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_58 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_57 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_56 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_55 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_54 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_53 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_52 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_51 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_50 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_49 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_48 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<2> ), .Y(n36) );
  INVX1 U3 ( .A(\q<3> ), .Y(n33) );
  INVX1 U4 ( .A(\q<5> ), .Y(n27) );
  INVX1 U5 ( .A(\q<6> ), .Y(n24) );
  INVX1 U6 ( .A(\q<1> ), .Y(n39) );
  INVX1 U7 ( .A(\q<4> ), .Y(n30) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(\q<9> ), .Y(n18) );
  INVX1 U11 ( .A(\q<10> ), .Y(n16) );
  INVX1 U12 ( .A(\q<11> ), .Y(n14) );
  INVX1 U13 ( .A(\q<12> ), .Y(n12) );
  INVX1 U14 ( .A(\q<13> ), .Y(n10) );
  INVX1 U15 ( .A(\q<14> ), .Y(n8) );
  INVX1 U16 ( .A(\q<15> ), .Y(n6) );
  INVX1 U17 ( .A(rst), .Y(n4) );
  INVX1 U18 ( .A(n4), .Y(n3) );
  INVX1 U19 ( .A(\d<6> ), .Y(n25) );
  INVX1 U20 ( .A(\d<15> ), .Y(n5) );
  INVX1 U21 ( .A(\d<13> ), .Y(n9) );
  INVX1 U22 ( .A(\d<12> ), .Y(n11) );
  INVX1 U23 ( .A(\d<11> ), .Y(n13) );
  INVX1 U24 ( .A(\d<10> ), .Y(n15) );
  INVX1 U25 ( .A(\d<9> ), .Y(n17) );
  INVX1 U26 ( .A(\d<8> ), .Y(n19) );
  OAI21X1 U27 ( .A(n2), .B(n28), .C(n29), .Y(n47) );
  INVX1 U28 ( .A(\d<5> ), .Y(n28) );
  OAI21X1 U29 ( .A(n2), .B(n22), .C(n23), .Y(n45) );
  OAI21X1 U30 ( .A(n43), .B(n2), .C(n44), .Y(n52) );
  INVX2 U31 ( .A(wr_en), .Y(n2) );
  INVX1 U32 ( .A(\d<14> ), .Y(n7) );
  INVX1 U33 ( .A(\d<1> ), .Y(n40) );
  INVX1 U34 ( .A(\d<0> ), .Y(n43) );
  INVX1 U35 ( .A(\d<2> ), .Y(n37) );
  INVX1 U36 ( .A(\d<4> ), .Y(n31) );
  INVX1 U37 ( .A(\d<3> ), .Y(n34) );
  INVX1 U38 ( .A(\d<7> ), .Y(n22) );
  INVX8 U39 ( .A(n2), .Y(n1) );
  MUX2X1 U40 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  MUX2X1 U41 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  MUX2X1 U42 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  MUX2X1 U43 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  MUX2X1 U44 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  MUX2X1 U45 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  MUX2X1 U46 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U47 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U48 ( .A(n1), .B(n21), .Y(n23) );
  OR2X2 U49 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U50 ( .A(n26), .B(n2), .C(n25), .D(n26), .Y(n46) );
  OR2X2 U51 ( .A(n1), .B(n27), .Y(n29) );
  OR2X2 U52 ( .A(n1), .B(n30), .Y(n32) );
  AOI22X1 U53 ( .A(n32), .B(n2), .C(n32), .D(n31), .Y(n48) );
  OR2X2 U54 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U55 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U56 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U57 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U58 ( .A(n1), .B(n39), .Y(n41) );
  AOI22X1 U59 ( .A(n41), .B(n2), .C(n41), .D(n40), .Y(n51) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_4 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_79 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_78 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(n3) );
  dff_77 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(rst) );
  dff_76 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_75 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_74 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_73 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_72 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_71 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_70 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_69 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_68 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_67 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_66 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_65 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_64 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<1> ), .Y(n39) );
  INVX1 U3 ( .A(\q<2> ), .Y(n36) );
  INVX1 U4 ( .A(\q<3> ), .Y(n33) );
  INVX1 U5 ( .A(\q<5> ), .Y(n27) );
  INVX1 U6 ( .A(\q<4> ), .Y(n30) );
  INVX1 U7 ( .A(\q<6> ), .Y(n24) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(\q<14> ), .Y(n8) );
  INVX1 U11 ( .A(rst), .Y(n4) );
  INVX1 U12 ( .A(n4), .Y(n3) );
  INVX1 U13 ( .A(\d<8> ), .Y(n19) );
  INVX1 U14 ( .A(\d<12> ), .Y(n11) );
  INVX1 U15 ( .A(\d<11> ), .Y(n13) );
  INVX1 U16 ( .A(\d<9> ), .Y(n17) );
  INVX1 U17 ( .A(\d<10> ), .Y(n15) );
  INVX1 U18 ( .A(\d<15> ), .Y(n5) );
  INVX1 U19 ( .A(\d<13> ), .Y(n9) );
  INVX1 U20 ( .A(\d<14> ), .Y(n7) );
  OAI21X1 U21 ( .A(n2), .B(n40), .C(n41), .Y(n51) );
  INVX1 U22 ( .A(\d<1> ), .Y(n40) );
  OAI21X1 U23 ( .A(n2), .B(n28), .C(n29), .Y(n47) );
  INVX1 U24 ( .A(\d<5> ), .Y(n28) );
  OAI21X1 U25 ( .A(n43), .B(n2), .C(n44), .Y(n52) );
  INVX2 U26 ( .A(wr_en), .Y(n2) );
  INVX1 U27 ( .A(\d<0> ), .Y(n43) );
  INVX1 U28 ( .A(\d<2> ), .Y(n37) );
  INVX1 U29 ( .A(\d<4> ), .Y(n31) );
  INVX1 U30 ( .A(\d<6> ), .Y(n25) );
  INVX1 U31 ( .A(\d<3> ), .Y(n34) );
  INVX1 U32 ( .A(\d<7> ), .Y(n22) );
  INVX8 U33 ( .A(n2), .Y(n1) );
  INVX2 U34 ( .A(\q<15> ), .Y(n6) );
  MUX2X1 U35 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  MUX2X1 U36 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  INVX2 U37 ( .A(\q<13> ), .Y(n10) );
  MUX2X1 U38 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  INVX2 U39 ( .A(\q<12> ), .Y(n12) );
  MUX2X1 U40 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  INVX2 U41 ( .A(\q<11> ), .Y(n14) );
  MUX2X1 U42 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  INVX2 U43 ( .A(\q<10> ), .Y(n16) );
  MUX2X1 U44 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  INVX2 U45 ( .A(\q<9> ), .Y(n18) );
  MUX2X1 U46 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U47 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U48 ( .A(n1), .B(n21), .Y(n23) );
  AOI22X1 U49 ( .A(n23), .B(n2), .C(n23), .D(n22), .Y(n45) );
  OR2X2 U50 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U51 ( .A(n26), .B(n2), .C(n26), .D(n25), .Y(n46) );
  OR2X2 U52 ( .A(n1), .B(n27), .Y(n29) );
  OR2X2 U53 ( .A(n1), .B(n30), .Y(n32) );
  AOI22X1 U54 ( .A(n32), .B(n2), .C(n32), .D(n31), .Y(n48) );
  OR2X2 U55 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U56 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U57 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U58 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U59 ( .A(n1), .B(n39), .Y(n41) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_5 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_95 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_94 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(n3) );
  dff_93 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(rst) );
  dff_92 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_91 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_90 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_89 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_88 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_87 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_86 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_85 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_84 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_83 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_82 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_81 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_80 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<1> ), .Y(n39) );
  INVX1 U3 ( .A(\q<2> ), .Y(n36) );
  INVX1 U4 ( .A(\q<3> ), .Y(n33) );
  INVX1 U5 ( .A(\q<5> ), .Y(n27) );
  INVX1 U6 ( .A(\q<6> ), .Y(n24) );
  INVX1 U7 ( .A(\q<4> ), .Y(n30) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(\q<14> ), .Y(n8) );
  INVX1 U11 ( .A(rst), .Y(n4) );
  INVX1 U12 ( .A(n4), .Y(n3) );
  INVX1 U13 ( .A(\d<8> ), .Y(n19) );
  INVX1 U14 ( .A(\d<12> ), .Y(n11) );
  INVX1 U15 ( .A(\d<11> ), .Y(n13) );
  INVX1 U16 ( .A(\d<9> ), .Y(n17) );
  INVX1 U17 ( .A(\d<10> ), .Y(n15) );
  INVX1 U18 ( .A(\d<15> ), .Y(n5) );
  INVX1 U19 ( .A(\d<13> ), .Y(n9) );
  INVX1 U20 ( .A(\d<14> ), .Y(n7) );
  OAI21X1 U21 ( .A(n2), .B(n40), .C(n41), .Y(n51) );
  INVX1 U22 ( .A(\d<1> ), .Y(n40) );
  OAI21X1 U23 ( .A(n2), .B(n28), .C(n29), .Y(n47) );
  INVX1 U24 ( .A(\d<5> ), .Y(n28) );
  OAI21X1 U25 ( .A(n2), .B(n22), .C(n23), .Y(n45) );
  OAI21X1 U26 ( .A(n2), .B(n43), .C(n44), .Y(n52) );
  INVX2 U27 ( .A(wr_en), .Y(n2) );
  INVX1 U28 ( .A(\d<0> ), .Y(n43) );
  INVX1 U29 ( .A(\d<2> ), .Y(n37) );
  INVX1 U30 ( .A(\d<3> ), .Y(n34) );
  INVX1 U31 ( .A(\d<4> ), .Y(n31) );
  INVX1 U32 ( .A(\d<6> ), .Y(n25) );
  INVX1 U33 ( .A(\d<7> ), .Y(n22) );
  INVX8 U34 ( .A(n2), .Y(n1) );
  INVX2 U35 ( .A(\q<15> ), .Y(n6) );
  MUX2X1 U36 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  MUX2X1 U37 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  INVX2 U38 ( .A(\q<13> ), .Y(n10) );
  MUX2X1 U39 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  INVX2 U40 ( .A(\q<12> ), .Y(n12) );
  MUX2X1 U41 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  INVX2 U42 ( .A(\q<11> ), .Y(n14) );
  MUX2X1 U43 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  INVX2 U44 ( .A(\q<10> ), .Y(n16) );
  MUX2X1 U45 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  INVX2 U46 ( .A(\q<9> ), .Y(n18) );
  MUX2X1 U47 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U48 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U49 ( .A(n1), .B(n21), .Y(n23) );
  OR2X2 U50 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U51 ( .A(n26), .B(n2), .C(n26), .D(n25), .Y(n46) );
  OR2X2 U52 ( .A(n1), .B(n27), .Y(n29) );
  OR2X2 U53 ( .A(n1), .B(n30), .Y(n32) );
  AOI22X1 U54 ( .A(n32), .B(n2), .C(n32), .D(n31), .Y(n48) );
  OR2X2 U55 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U56 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U57 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U58 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U59 ( .A(n1), .B(n39), .Y(n41) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_6 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_111 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_110 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(n3) );
  dff_109 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(rst) );
  dff_108 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_107 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_106 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_105 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_104 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_103 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_102 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_101 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_100 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_99 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_98 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_97 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_96 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<1> ), .Y(n39) );
  INVX1 U3 ( .A(\q<2> ), .Y(n36) );
  INVX1 U4 ( .A(\q<3> ), .Y(n33) );
  INVX1 U5 ( .A(\q<4> ), .Y(n30) );
  INVX1 U6 ( .A(\q<5> ), .Y(n27) );
  INVX1 U7 ( .A(\q<6> ), .Y(n24) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(\q<11> ), .Y(n14) );
  INVX1 U11 ( .A(\q<12> ), .Y(n12) );
  INVX1 U12 ( .A(\q<13> ), .Y(n10) );
  INVX1 U13 ( .A(\q<14> ), .Y(n8) );
  INVX1 U14 ( .A(\q<15> ), .Y(n6) );
  INVX1 U15 ( .A(rst), .Y(n4) );
  INVX1 U16 ( .A(n4), .Y(n3) );
  INVX1 U17 ( .A(\d<15> ), .Y(n5) );
  INVX1 U18 ( .A(\d<14> ), .Y(n7) );
  INVX1 U19 ( .A(\d<12> ), .Y(n11) );
  OAI21X1 U20 ( .A(n2), .B(n40), .C(n41), .Y(n51) );
  INVX1 U21 ( .A(\d<1> ), .Y(n40) );
  OAI21X1 U22 ( .A(n2), .B(n31), .C(n32), .Y(n48) );
  INVX1 U23 ( .A(\d<4> ), .Y(n31) );
  OAI21X1 U24 ( .A(n2), .B(n22), .C(n23), .Y(n45) );
  OAI21X1 U25 ( .A(n43), .B(n2), .C(n44), .Y(n52) );
  INVX2 U26 ( .A(wr_en), .Y(n2) );
  MUX2X1 U27 ( .B(n7), .A(n8), .S(n2), .Y(n59) );
  INVX1 U28 ( .A(\d<13> ), .Y(n9) );
  INVX1 U29 ( .A(\d<10> ), .Y(n15) );
  INVX1 U30 ( .A(\d<11> ), .Y(n13) );
  INVX1 U31 ( .A(\d<9> ), .Y(n17) );
  INVX1 U32 ( .A(\d<8> ), .Y(n19) );
  INVX1 U33 ( .A(\d<0> ), .Y(n43) );
  INVX1 U34 ( .A(\d<2> ), .Y(n37) );
  INVX1 U35 ( .A(\d<3> ), .Y(n34) );
  INVX1 U36 ( .A(\d<5> ), .Y(n28) );
  INVX1 U37 ( .A(\d<6> ), .Y(n25) );
  INVX1 U38 ( .A(\d<7> ), .Y(n22) );
  INVX8 U39 ( .A(n2), .Y(n1) );
  MUX2X1 U40 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  MUX2X1 U41 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  MUX2X1 U42 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  MUX2X1 U43 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  INVX2 U44 ( .A(\q<10> ), .Y(n16) );
  MUX2X1 U45 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  INVX2 U46 ( .A(\q<9> ), .Y(n18) );
  MUX2X1 U47 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U48 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U49 ( .A(n1), .B(n21), .Y(n23) );
  OR2X2 U50 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U51 ( .A(n26), .B(n2), .C(n26), .D(n25), .Y(n46) );
  OR2X2 U52 ( .A(n1), .B(n27), .Y(n29) );
  AOI22X1 U53 ( .A(n29), .B(n2), .C(n29), .D(n28), .Y(n47) );
  OR2X2 U54 ( .A(n1), .B(n30), .Y(n32) );
  OR2X2 U55 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U56 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U57 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U58 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U59 ( .A(n1), .B(n39), .Y(n41) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module register16_7 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  dff_112 \dff_arr[0]  ( .q(\q<0> ), .d(n52), .clk(clk), .rst(n3) );
  dff_113 \dff_arr[1]  ( .q(\q<1> ), .d(n51), .clk(clk), .rst(n3) );
  dff_114 \dff_arr[2]  ( .q(\q<2> ), .d(n50), .clk(clk), .rst(rst) );
  dff_115 \dff_arr[3]  ( .q(\q<3> ), .d(n49), .clk(clk), .rst(rst) );
  dff_116 \dff_arr[4]  ( .q(\q<4> ), .d(n48), .clk(clk), .rst(n3) );
  dff_117 \dff_arr[5]  ( .q(\q<5> ), .d(n47), .clk(clk), .rst(n3) );
  dff_118 \dff_arr[6]  ( .q(\q<6> ), .d(n46), .clk(clk), .rst(n3) );
  dff_119 \dff_arr[7]  ( .q(\q<7> ), .d(n45), .clk(clk), .rst(n3) );
  dff_120 \dff_arr[8]  ( .q(\q<8> ), .d(n53), .clk(clk), .rst(n3) );
  dff_121 \dff_arr[9]  ( .q(\q<9> ), .d(n54), .clk(clk), .rst(n3) );
  dff_122 \dff_arr[10]  ( .q(\q<10> ), .d(n55), .clk(clk), .rst(n3) );
  dff_123 \dff_arr[11]  ( .q(\q<11> ), .d(n56), .clk(clk), .rst(n3) );
  dff_124 \dff_arr[12]  ( .q(\q<12> ), .d(n57), .clk(clk), .rst(n3) );
  dff_125 \dff_arr[13]  ( .q(\q<13> ), .d(n58), .clk(clk), .rst(n3) );
  dff_126 \dff_arr[14]  ( .q(\q<14> ), .d(n59), .clk(clk), .rst(n3) );
  dff_127 \dff_arr[15]  ( .q(\q<15> ), .d(n60), .clk(clk), .rst(n3) );
  INVX1 U1 ( .A(\q<0> ), .Y(n42) );
  INVX1 U2 ( .A(\q<1> ), .Y(n39) );
  INVX1 U3 ( .A(\q<2> ), .Y(n36) );
  INVX1 U4 ( .A(\q<3> ), .Y(n33) );
  INVX1 U5 ( .A(\q<4> ), .Y(n30) );
  INVX1 U6 ( .A(\q<5> ), .Y(n27) );
  INVX1 U7 ( .A(\q<6> ), .Y(n24) );
  INVX1 U8 ( .A(\q<7> ), .Y(n21) );
  INVX1 U9 ( .A(\q<8> ), .Y(n20) );
  INVX1 U10 ( .A(\q<9> ), .Y(n18) );
  INVX1 U11 ( .A(\q<10> ), .Y(n16) );
  INVX1 U12 ( .A(\q<11> ), .Y(n14) );
  INVX1 U13 ( .A(\q<12> ), .Y(n12) );
  INVX1 U14 ( .A(\q<13> ), .Y(n10) );
  INVX1 U15 ( .A(\q<15> ), .Y(n6) );
  INVX1 U16 ( .A(rst), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n3) );
  INVX1 U18 ( .A(\d<15> ), .Y(n5) );
  INVX1 U19 ( .A(\d<13> ), .Y(n9) );
  INVX1 U20 ( .A(\d<12> ), .Y(n11) );
  INVX1 U21 ( .A(\d<11> ), .Y(n13) );
  INVX1 U22 ( .A(\d<10> ), .Y(n15) );
  INVX1 U23 ( .A(\d<9> ), .Y(n17) );
  INVX1 U24 ( .A(\d<8> ), .Y(n19) );
  OAI21X1 U25 ( .A(n2), .B(n40), .C(n41), .Y(n51) );
  INVX1 U26 ( .A(\d<1> ), .Y(n40) );
  OAI21X1 U27 ( .A(n2), .B(n28), .C(n29), .Y(n47) );
  INVX1 U28 ( .A(\d<5> ), .Y(n28) );
  OAI21X1 U29 ( .A(n2), .B(n31), .C(n32), .Y(n48) );
  INVX1 U30 ( .A(\d<4> ), .Y(n31) );
  OAI21X1 U31 ( .A(n2), .B(n22), .C(n23), .Y(n45) );
  OAI21X1 U32 ( .A(n2), .B(n43), .C(n44), .Y(n52) );
  INVX2 U33 ( .A(wr_en), .Y(n2) );
  INVX1 U34 ( .A(\d<14> ), .Y(n7) );
  INVX1 U35 ( .A(\d<0> ), .Y(n43) );
  INVX1 U36 ( .A(\d<2> ), .Y(n37) );
  INVX1 U37 ( .A(\d<3> ), .Y(n34) );
  INVX1 U38 ( .A(\d<6> ), .Y(n25) );
  INVX1 U39 ( .A(\d<7> ), .Y(n22) );
  INVX8 U40 ( .A(n2), .Y(n1) );
  MUX2X1 U41 ( .B(n6), .A(n5), .S(n1), .Y(n60) );
  INVX2 U42 ( .A(\q<14> ), .Y(n8) );
  MUX2X1 U43 ( .B(n8), .A(n7), .S(n1), .Y(n59) );
  MUX2X1 U44 ( .B(n10), .A(n9), .S(n1), .Y(n58) );
  MUX2X1 U45 ( .B(n12), .A(n11), .S(n1), .Y(n57) );
  MUX2X1 U46 ( .B(n14), .A(n13), .S(n1), .Y(n56) );
  MUX2X1 U47 ( .B(n16), .A(n15), .S(n1), .Y(n55) );
  MUX2X1 U48 ( .B(n18), .A(n17), .S(n1), .Y(n54) );
  MUX2X1 U49 ( .B(n20), .A(n19), .S(n1), .Y(n53) );
  OR2X2 U50 ( .A(n1), .B(n21), .Y(n23) );
  OR2X2 U51 ( .A(n1), .B(n24), .Y(n26) );
  AOI22X1 U52 ( .A(n26), .B(n2), .C(n26), .D(n25), .Y(n46) );
  OR2X2 U53 ( .A(n1), .B(n27), .Y(n29) );
  OR2X2 U54 ( .A(n1), .B(n30), .Y(n32) );
  OR2X2 U55 ( .A(n1), .B(n33), .Y(n35) );
  AOI22X1 U56 ( .A(n35), .B(n2), .C(n35), .D(n34), .Y(n49) );
  OR2X2 U57 ( .A(n1), .B(n36), .Y(n38) );
  AOI22X1 U58 ( .A(n38), .B(n2), .C(n38), .D(n37), .Y(n50) );
  OR2X2 U59 ( .A(n1), .B(n39), .Y(n41) );
  OR2X2 U60 ( .A(n1), .B(n42), .Y(n44) );
endmodule


module decoder3to8 ( .In({\In<2> , \In<1> , \In<0> }), .Out({\Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<2> , \In<1> , \In<0> ;
  output \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> ,
         \Out<0> ;
  wire   n1, n2, n3;

  NOR3X1 U4 ( .A(n3), .B(n1), .C(n2), .Y(\Out<7> ) );
  NOR3X1 U5 ( .A(n3), .B(\In<0> ), .C(n2), .Y(\Out<6> ) );
  NOR3X1 U6 ( .A(n3), .B(\In<1> ), .C(n1), .Y(\Out<5> ) );
  NOR3X1 U7 ( .A(n3), .B(\In<1> ), .C(\In<0> ), .Y(\Out<4> ) );
  NOR3X1 U8 ( .A(n2), .B(\In<2> ), .C(n1), .Y(\Out<3> ) );
  NOR3X1 U9 ( .A(n2), .B(\In<2> ), .C(\In<0> ), .Y(\Out<2> ) );
  NOR3X1 U10 ( .A(n1), .B(\In<2> ), .C(\In<1> ), .Y(\Out<1> ) );
  NOR3X1 U11 ( .A(\In<0> ), .B(\In<2> ), .C(\In<1> ), .Y(\Out<0> ) );
  INVX1 U1 ( .A(\In<0> ), .Y(n1) );
  INVX1 U2 ( .A(\In<1> ), .Y(n2) );
  INVX1 U3 ( .A(\In<2> ), .Y(n3) );
endmodule


module mux8to1_16_1 ( .In({\In<127> , \In<126> , \In<125> , \In<124> , 
        \In<123> , \In<122> , \In<121> , \In<120> , \In<119> , \In<118> , 
        \In<117> , \In<116> , \In<115> , \In<114> , \In<113> , \In<112> , 
        \In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , 
        \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , 
        \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , 
        \In<78> , \In<77> , \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , 
        \In<71> , \In<70> , \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , 
        \In<64> , \In<63> , \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , 
        \In<57> , \In<56> , \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , 
        \In<50> , \In<49> , \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , 
        \In<43> , \In<42> , \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , 
        \In<36> , \In<35> , \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , 
        \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , 
        \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , 
        \In<0> }), .Sel({\Sel<2> , \Sel<1> , \Sel<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<127> , \In<126> , \In<125> , \In<124> , \In<123> , \In<122> ,
         \In<121> , \In<120> , \In<119> , \In<118> , \In<117> , \In<116> ,
         \In<115> , \In<114> , \In<113> , \In<112> , \In<111> , \In<110> ,
         \In<109> , \In<108> , \In<107> , \In<106> , \In<105> , \In<104> ,
         \In<103> , \In<102> , \In<101> , \In<100> , \In<99> , \In<98> ,
         \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , \In<92> , \In<91> ,
         \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , \In<85> , \In<84> ,
         \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , \In<78> , \In<77> ,
         \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , \In<71> , \In<70> ,
         \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , \In<64> , \In<63> ,
         \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , \In<57> , \In<56> ,
         \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , \In<50> , \In<49> ,
         \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> ,
         \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> ,
         \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , \In<29> , \In<28> ,
         \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , \In<22> , \In<21> ,
         \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , \In<15> , \In<14> ,
         \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , \In<8> , \In<7> ,
         \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , \In<0> ,
         \Sel<2> , \Sel<1> , \Sel<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \mux0_out<15> , \mux0_out<14> , \mux0_out<13> , \mux0_out<12> ,
         \mux0_out<11> , \mux0_out<10> , \mux0_out<9> , \mux0_out<8> ,
         \mux0_out<7> , \mux0_out<6> , \mux0_out<5> , \mux0_out<4> ,
         \mux0_out<3> , \mux0_out<2> , \mux0_out<1> , \mux0_out<0> ,
         \mux1_out<15> , \mux1_out<14> , \mux1_out<13> , \mux1_out<12> ,
         \mux1_out<11> , \mux1_out<10> , \mux1_out<9> , \mux1_out<8> ,
         \mux1_out<7> , \mux1_out<6> , \mux1_out<5> , \mux1_out<4> ,
         \mux1_out<3> , \mux1_out<2> , \mux1_out<1> , \mux1_out<0> , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38;

  mux4to1_16_4 mux0 ( .InA({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .InB({\In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> }), 
        .InC({\In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> , 
        \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> , 
        \In<34> , \In<33> , \In<32> }), .InD({\In<63> , \In<62> , \In<61> , 
        \In<60> , \In<59> , \In<58> , \In<57> , \In<56> , \In<55> , \In<54> , 
        \In<53> , \In<52> , \In<51> , \In<50> , \In<49> , \In<48> }), .S({
        \Sel<1> , \Sel<0> }), .Out({\mux0_out<15> , \mux0_out<14> , 
        \mux0_out<13> , \mux0_out<12> , \mux0_out<11> , \mux0_out<10> , 
        \mux0_out<9> , \mux0_out<8> , \mux0_out<7> , \mux0_out<6> , 
        \mux0_out<5> , \mux0_out<4> , \mux0_out<3> , \mux0_out<2> , 
        \mux0_out<1> , \mux0_out<0> }) );
  mux4to1_16_3 mux1 ( .InA({\In<79> , \In<78> , \In<77> , \In<76> , \In<75> , 
        \In<74> , \In<73> , \In<72> , \In<71> , \In<70> , \In<69> , \In<68> , 
        \In<67> , \In<66> , \In<65> , \In<64> }), .InB({\In<95> , \In<94> , 
        \In<93> , \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , 
        \In<86> , \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> }), 
        .InC({\In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> }), .InD({\In<127> , \In<126> , 
        \In<125> , \In<124> , \In<123> , \In<122> , \In<121> , \In<120> , 
        \In<119> , \In<118> , \In<117> , \In<116> , \In<115> , \In<114> , 
        \In<113> , \In<112> }), .S({\Sel<1> , \Sel<0> }), .Out({\mux1_out<15> , 
        \mux1_out<14> , \mux1_out<13> , \mux1_out<12> , \mux1_out<11> , 
        \mux1_out<10> , \mux1_out<9> , \mux1_out<8> , \mux1_out<7> , 
        \mux1_out<6> , \mux1_out<5> , \mux1_out<4> , \mux1_out<3> , 
        \mux1_out<2> , \mux1_out<1> , \mux1_out<0> }) );
  INVX1 U1 ( .A(n6), .Y(n3) );
  INVX1 U2 ( .A(n4), .Y(n2) );
  INVX1 U3 ( .A(n4), .Y(n1) );
  MUX2X1 U4 ( .B(n22), .A(n21), .S(n1), .Y(\Out<7> ) );
  MUX2X1 U5 ( .B(n16), .A(n15), .S(n2), .Y(\Out<4> ) );
  MUX2X1 U6 ( .B(n27), .A(n28), .S(n3), .Y(\Out<10> ) );
  INVX1 U7 ( .A(\mux1_out<8> ), .Y(n23) );
  INVX1 U8 ( .A(\mux1_out<9> ), .Y(n25) );
  INVX1 U9 ( .A(\mux1_out<11> ), .Y(n29) );
  INVX1 U10 ( .A(\mux1_out<12> ), .Y(n31) );
  INVX1 U11 ( .A(\mux1_out<13> ), .Y(n33) );
  INVX1 U12 ( .A(\mux1_out<14> ), .Y(n35) );
  INVX1 U13 ( .A(\mux1_out<15> ), .Y(n37) );
  INVX1 U14 ( .A(\mux0_out<8> ), .Y(n24) );
  INVX1 U15 ( .A(\mux0_out<12> ), .Y(n32) );
  INVX1 U16 ( .A(\mux0_out<13> ), .Y(n34) );
  INVX1 U17 ( .A(\mux0_out<14> ), .Y(n36) );
  INVX1 U18 ( .A(\mux0_out<15> ), .Y(n38) );
  INVX1 U19 ( .A(\mux1_out<10> ), .Y(n27) );
  MUX2X1 U20 ( .B(n19), .A(n20), .S(n4), .Y(\Out<6> ) );
  INVX4 U21 ( .A(n5), .Y(n4) );
  INVX1 U22 ( .A(\mux1_out<7> ), .Y(n21) );
  INVX1 U23 ( .A(\mux0_out<7> ), .Y(n22) );
  INVX1 U24 ( .A(\mux0_out<9> ), .Y(n26) );
  INVX1 U25 ( .A(\mux1_out<4> ), .Y(n15) );
  INVX1 U26 ( .A(\mux1_out<5> ), .Y(n17) );
  INVX1 U27 ( .A(\mux0_out<4> ), .Y(n16) );
  INVX1 U28 ( .A(\mux0_out<11> ), .Y(n30) );
  INVX1 U29 ( .A(\mux0_out<5> ), .Y(n18) );
  INVX1 U30 ( .A(\mux0_out<2> ), .Y(n12) );
  INVX1 U31 ( .A(\mux0_out<10> ), .Y(n28) );
  INVX1 U32 ( .A(\mux0_out<6> ), .Y(n20) );
  INVX1 U33 ( .A(\mux1_out<6> ), .Y(n19) );
  INVX1 U34 ( .A(\mux1_out<2> ), .Y(n11) );
  INVX1 U35 ( .A(\mux1_out<3> ), .Y(n13) );
  INVX1 U36 ( .A(\mux0_out<3> ), .Y(n14) );
  INVX1 U37 ( .A(\mux1_out<0> ), .Y(n7) );
  INVX1 U38 ( .A(\mux0_out<0> ), .Y(n8) );
  INVX1 U39 ( .A(\mux1_out<1> ), .Y(n9) );
  INVX1 U40 ( .A(\mux0_out<1> ), .Y(n10) );
  BUFX4 U41 ( .A(\Sel<2> ), .Y(n5) );
  BUFX4 U42 ( .A(\Sel<2> ), .Y(n6) );
  MUX2X1 U43 ( .B(n8), .A(n7), .S(n5), .Y(\Out<0> ) );
  MUX2X1 U44 ( .B(n10), .A(n9), .S(n5), .Y(\Out<1> ) );
  MUX2X1 U45 ( .B(n12), .A(n11), .S(n5), .Y(\Out<2> ) );
  MUX2X1 U46 ( .B(n14), .A(n13), .S(n5), .Y(\Out<3> ) );
  MUX2X1 U47 ( .B(n18), .A(n17), .S(n5), .Y(\Out<5> ) );
  MUX2X1 U48 ( .B(n24), .A(n23), .S(n6), .Y(\Out<8> ) );
  MUX2X1 U49 ( .B(n26), .A(n25), .S(n6), .Y(\Out<9> ) );
  MUX2X1 U50 ( .B(n30), .A(n29), .S(n6), .Y(\Out<11> ) );
  MUX2X1 U51 ( .B(n32), .A(n31), .S(n6), .Y(\Out<12> ) );
  MUX2X1 U52 ( .B(n34), .A(n33), .S(n6), .Y(\Out<13> ) );
  MUX2X1 U53 ( .B(n36), .A(n35), .S(n6), .Y(\Out<14> ) );
  MUX2X1 U54 ( .B(n38), .A(n37), .S(n6), .Y(\Out<15> ) );
endmodule


module mux8to1_16_0 ( .In({\In<127> , \In<126> , \In<125> , \In<124> , 
        \In<123> , \In<122> , \In<121> , \In<120> , \In<119> , \In<118> , 
        \In<117> , \In<116> , \In<115> , \In<114> , \In<113> , \In<112> , 
        \In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , 
        \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , 
        \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , 
        \In<78> , \In<77> , \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , 
        \In<71> , \In<70> , \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , 
        \In<64> , \In<63> , \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , 
        \In<57> , \In<56> , \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , 
        \In<50> , \In<49> , \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , 
        \In<43> , \In<42> , \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , 
        \In<36> , \In<35> , \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , 
        \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , 
        \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , 
        \In<0> }), .Sel({\Sel<2> , \Sel<1> , \Sel<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<127> , \In<126> , \In<125> , \In<124> , \In<123> , \In<122> ,
         \In<121> , \In<120> , \In<119> , \In<118> , \In<117> , \In<116> ,
         \In<115> , \In<114> , \In<113> , \In<112> , \In<111> , \In<110> ,
         \In<109> , \In<108> , \In<107> , \In<106> , \In<105> , \In<104> ,
         \In<103> , \In<102> , \In<101> , \In<100> , \In<99> , \In<98> ,
         \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , \In<92> , \In<91> ,
         \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , \In<85> , \In<84> ,
         \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , \In<78> , \In<77> ,
         \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , \In<71> , \In<70> ,
         \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , \In<64> , \In<63> ,
         \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , \In<57> , \In<56> ,
         \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , \In<50> , \In<49> ,
         \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> ,
         \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> ,
         \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , \In<29> , \In<28> ,
         \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , \In<22> , \In<21> ,
         \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , \In<15> , \In<14> ,
         \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , \In<8> , \In<7> ,
         \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , \In<0> ,
         \Sel<2> , \Sel<1> , \Sel<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \mux0_out<15> , \mux0_out<14> , \mux0_out<13> , \mux0_out<12> ,
         \mux0_out<11> , \mux0_out<10> , \mux0_out<9> , \mux0_out<8> ,
         \mux0_out<7> , \mux0_out<6> , \mux0_out<5> , \mux0_out<4> ,
         \mux0_out<3> , \mux0_out<2> , \mux0_out<1> , \mux0_out<0> ,
         \mux1_out<15> , \mux1_out<14> , \mux1_out<13> , \mux1_out<12> ,
         \mux1_out<11> , \mux1_out<10> , \mux1_out<9> , \mux1_out<8> ,
         \mux1_out<7> , \mux1_out<6> , \mux1_out<5> , \mux1_out<4> ,
         \mux1_out<3> , \mux1_out<2> , \mux1_out<1> , \mux1_out<0> , n1, n2,
         n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n32, n33, n34, n35, n36, n37, n38, n39;

  mux4to1_16_2 mux0 ( .InA({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .InB({\In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> }), 
        .InC({\In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> , 
        \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> , 
        \In<34> , \In<33> , \In<32> }), .InD({\In<63> , \In<62> , \In<61> , 
        \In<60> , \In<59> , \In<58> , \In<57> , \In<56> , \In<55> , \In<54> , 
        \In<53> , \In<52> , \In<51> , \In<50> , \In<49> , \In<48> }), .S({
        \Sel<1> , \Sel<0> }), .Out({\mux0_out<15> , \mux0_out<14> , 
        \mux0_out<13> , \mux0_out<12> , \mux0_out<11> , \mux0_out<10> , 
        \mux0_out<9> , \mux0_out<8> , \mux0_out<7> , \mux0_out<6> , 
        \mux0_out<5> , \mux0_out<4> , \mux0_out<3> , \mux0_out<2> , 
        \mux0_out<1> , \mux0_out<0> }) );
  mux4to1_16_1 mux1 ( .InA({\In<79> , \In<78> , \In<77> , \In<76> , \In<75> , 
        \In<74> , \In<73> , \In<72> , \In<71> , \In<70> , \In<69> , \In<68> , 
        \In<67> , \In<66> , \In<65> , \In<64> }), .InB({\In<95> , \In<94> , 
        \In<93> , \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , 
        \In<86> , \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> }), 
        .InC({\In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> }), .InD({\In<127> , \In<126> , 
        \In<125> , \In<124> , \In<123> , \In<122> , \In<121> , \In<120> , 
        \In<119> , \In<118> , \In<117> , \In<116> , \In<115> , \In<114> , 
        \In<113> , \In<112> }), .S({\Sel<1> , \Sel<0> }), .Out({\mux1_out<15> , 
        \mux1_out<14> , \mux1_out<13> , \mux1_out<12> , \mux1_out<11> , 
        \mux1_out<10> , \mux1_out<9> , \mux1_out<8> , \mux1_out<7> , 
        \mux1_out<6> , \mux1_out<5> , \mux1_out<4> , \mux1_out<3> , 
        \mux1_out<2> , \mux1_out<1> , \mux1_out<0> }) );
  MUX2X1 U1 ( .B(n34), .A(n35), .S(n2), .Y(\Out<3> ) );
  INVX4 U2 ( .A(\Sel<2> ), .Y(n2) );
  MUX2X1 U3 ( .B(\mux0_out<9> ), .A(\mux1_out<9> ), .S(n1), .Y(n13) );
  INVX8 U4 ( .A(n2), .Y(n1) );
  MUX2X1 U5 ( .B(\mux0_out<0> ), .A(\mux1_out<0> ), .S(n21), .Y(n18) );
  MUX2X1 U6 ( .B(\mux1_out<14> ), .A(\mux0_out<14> ), .S(n2), .Y(n12) );
  INVX1 U7 ( .A(n17), .Y(\Out<4> ) );
  MUX2X1 U8 ( .B(\mux1_out<4> ), .A(\mux0_out<4> ), .S(n2), .Y(n17) );
  MUX2X1 U9 ( .B(\mux0_out<10> ), .A(\mux1_out<10> ), .S(n21), .Y(n14) );
  MUX2X1 U10 ( .B(n37), .A(n36), .S(n20), .Y(\Out<5> ) );
  INVX1 U11 ( .A(n11), .Y(\Out<13> ) );
  INVX1 U12 ( .A(n12), .Y(\Out<14> ) );
  MUX2X1 U13 ( .B(n33), .A(n32), .S(n20), .Y(\Out<2> ) );
  INVX1 U14 ( .A(n10), .Y(\Out<12> ) );
  MUX2X1 U15 ( .B(n4), .A(n5), .S(n20), .Y(\Out<6> ) );
  INVX1 U16 ( .A(\mux0_out<6> ), .Y(n4) );
  INVX1 U17 ( .A(\mux1_out<6> ), .Y(n5) );
  MUX2X1 U18 ( .B(n7), .A(n8), .S(n20), .Y(\Out<1> ) );
  INVX1 U19 ( .A(\mux0_out<1> ), .Y(n7) );
  INVX1 U20 ( .A(\mux1_out<1> ), .Y(n8) );
  BUFX2 U21 ( .A(\mux0_out<13> ), .Y(n9) );
  INVX1 U22 ( .A(\mux1_out<15> ), .Y(n38) );
  INVX1 U23 ( .A(\mux0_out<15> ), .Y(n39) );
  INVX1 U24 ( .A(n15), .Y(\Out<8> ) );
  INVX1 U25 ( .A(n13), .Y(\Out<9> ) );
  INVX1 U26 ( .A(n14), .Y(\Out<10> ) );
  INVX1 U27 ( .A(n16), .Y(\Out<11> ) );
  MUX2X1 U28 ( .B(\mux0_out<12> ), .A(\mux1_out<12> ), .S(n21), .Y(n10) );
  MUX2X1 U29 ( .B(n9), .A(\mux1_out<13> ), .S(n21), .Y(n11) );
  INVX1 U30 ( .A(n19), .Y(\Out<7> ) );
  MUX2X1 U31 ( .B(\mux0_out<11> ), .A(\mux1_out<11> ), .S(n21), .Y(n16) );
  INVX1 U32 ( .A(n18), .Y(\Out<0> ) );
  MUX2X1 U33 ( .B(\mux0_out<8> ), .A(\mux1_out<8> ), .S(n21), .Y(n15) );
  INVX1 U34 ( .A(\mux1_out<3> ), .Y(n34) );
  MUX2X1 U35 ( .B(\mux0_out<7> ), .A(\mux1_out<7> ), .S(n20), .Y(n19) );
  INVX1 U36 ( .A(\mux1_out<5> ), .Y(n36) );
  INVX1 U37 ( .A(\mux0_out<5> ), .Y(n37) );
  INVX1 U38 ( .A(\mux1_out<2> ), .Y(n32) );
  INVX1 U39 ( .A(\mux0_out<2> ), .Y(n33) );
  INVX1 U40 ( .A(\mux0_out<3> ), .Y(n35) );
  BUFX4 U41 ( .A(\Sel<2> ), .Y(n20) );
  BUFX4 U42 ( .A(\Sel<2> ), .Y(n21) );
  MUX2X1 U43 ( .B(n39), .A(n38), .S(n21), .Y(\Out<15> ) );
endmodule


module demux1to8_16 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<2> , \S<1> , \S<0> }), 
    .Out0({\Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , 
        \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , 
        \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({
        \Out1<15> , \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , 
        \Out1<9> , \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , 
        \Out1<3> , \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , 
        \Out2<14> , \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , 
        \Out2<8> , \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , 
        \Out2<2> , \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , 
        \Out3<13> , \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , 
        \Out3<7> , \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , 
        \Out3<1> , \Out3<0> }), .Out4({\Out4<15> , \Out4<14> , \Out4<13> , 
        \Out4<12> , \Out4<11> , \Out4<10> , \Out4<9> , \Out4<8> , \Out4<7> , 
        \Out4<6> , \Out4<5> , \Out4<4> , \Out4<3> , \Out4<2> , \Out4<1> , 
        \Out4<0> }), .Out5({\Out5<15> , \Out5<14> , \Out5<13> , \Out5<12> , 
        \Out5<11> , \Out5<10> , \Out5<9> , \Out5<8> , \Out5<7> , \Out5<6> , 
        \Out5<5> , \Out5<4> , \Out5<3> , \Out5<2> , \Out5<1> , \Out5<0> }), 
    .Out6({\Out6<15> , \Out6<14> , \Out6<13> , \Out6<12> , \Out6<11> , 
        \Out6<10> , \Out6<9> , \Out6<8> , \Out6<7> , \Out6<6> , \Out6<5> , 
        \Out6<4> , \Out6<3> , \Out6<2> , \Out6<1> , \Out6<0> }), .Out7({
        \Out7<15> , \Out7<14> , \Out7<13> , \Out7<12> , \Out7<11> , \Out7<10> , 
        \Out7<9> , \Out7<8> , \Out7<7> , \Out7<6> , \Out7<5> , \Out7<4> , 
        \Out7<3> , \Out7<2> , \Out7<1> , \Out7<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<2> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> , \Out4<15> ,
         \Out4<14> , \Out4<13> , \Out4<12> , \Out4<11> , \Out4<10> , \Out4<9> ,
         \Out4<8> , \Out4<7> , \Out4<6> , \Out4<5> , \Out4<4> , \Out4<3> ,
         \Out4<2> , \Out4<1> , \Out4<0> , \Out5<15> , \Out5<14> , \Out5<13> ,
         \Out5<12> , \Out5<11> , \Out5<10> , \Out5<9> , \Out5<8> , \Out5<7> ,
         \Out5<6> , \Out5<5> , \Out5<4> , \Out5<3> , \Out5<2> , \Out5<1> ,
         \Out5<0> , \Out6<15> , \Out6<14> , \Out6<13> , \Out6<12> , \Out6<11> ,
         \Out6<10> , \Out6<9> , \Out6<8> , \Out6<7> , \Out6<6> , \Out6<5> ,
         \Out6<4> , \Out6<3> , \Out6<2> , \Out6<1> , \Out6<0> , \Out7<15> ,
         \Out7<14> , \Out7<13> , \Out7<12> , \Out7<11> , \Out7<10> , \Out7<9> ,
         \Out7<8> , \Out7<7> , \Out7<6> , \Out7<5> , \Out7<4> , \Out7<3> ,
         \Out7<2> , \Out7<1> , \Out7<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7;

  demux1to8_0 \demux[0]  ( .In(\In<0> ), .S({n6, n3, n1}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ), .Out4(\Out4<0> ), 
        .Out5(\Out5<0> ), .Out6(\Out6<0> ), .Out7(\Out7<0> ) );
  demux1to8_1 \demux[1]  ( .In(\In<1> ), .S({n5, n3, n1}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ), .Out4(\Out4<1> ), 
        .Out5(\Out5<1> ), .Out6(\Out6<1> ), .Out7(\Out7<1> ) );
  demux1to8_2 \demux[2]  ( .In(\In<2> ), .S({n6, n3, \S<0> }), .Out0(\Out0<2> ), .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ), .Out4(\Out4<2> ), 
        .Out5(\Out5<2> ), .Out6(\Out6<2> ), .Out7(\Out7<2> ) );
  demux1to8_3 \demux[3]  ( .In(\In<3> ), .S({n6, n3, \S<0> }), .Out0(\Out0<3> ), .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ), .Out4(\Out4<3> ), 
        .Out5(\Out5<3> ), .Out6(\Out6<3> ), .Out7(\Out7<3> ) );
  demux1to8_4 \demux[4]  ( .In(\In<4> ), .S({n5, n3, n1}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ), .Out4(\Out4<4> ), 
        .Out5(\Out5<4> ), .Out6(\Out6<4> ), .Out7(\Out7<4> ) );
  demux1to8_5 \demux[5]  ( .In(\In<5> ), .S({n5, n3, n1}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ), .Out4(\Out4<5> ), 
        .Out5(\Out5<5> ), .Out6(\Out6<5> ), .Out7(\Out7<5> ) );
  demux1to8_6 \demux[6]  ( .In(\In<6> ), .S({n5, \S<1> , \S<0> }), .Out0(
        \Out0<6> ), .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ), 
        .Out4(\Out4<6> ), .Out5(\Out5<6> ), .Out6(\Out6<6> ), .Out7(\Out7<6> )
         );
  demux1to8_7 \demux[7]  ( .In(\In<7> ), .S({n5, \S<1> , \S<0> }), .Out0(
        \Out0<7> ), .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ), 
        .Out4(\Out4<7> ), .Out5(\Out5<7> ), .Out6(\Out6<7> ), .Out7(\Out7<7> )
         );
  demux1to8_8 \demux[8]  ( .In(\In<8> ), .S({n5, \S<1> , n1}), .Out0(\Out0<8> ), .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ), .Out4(\Out4<8> ), 
        .Out5(\Out5<8> ), .Out6(\Out6<8> ), .Out7(\Out7<8> ) );
  demux1to8_9 \demux[9]  ( .In(\In<9> ), .S({n5, \S<1> , \S<0> }), .Out0(
        \Out0<9> ), .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ), 
        .Out4(\Out4<9> ), .Out5(\Out5<9> ), .Out6(\Out6<9> ), .Out7(\Out7<9> )
         );
  demux1to8_10 \demux[10]  ( .In(\In<10> ), .S({n5, \S<1> , \S<0> }), .Out0(
        \Out0<10> ), .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ), 
        .Out4(\Out4<10> ), .Out5(\Out5<10> ), .Out6(\Out6<10> ), .Out7(
        \Out7<10> ) );
  demux1to8_11 \demux[11]  ( .In(\In<11> ), .S({n5, n3, \S<0> }), .Out0(
        \Out0<11> ), .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ), 
        .Out4(\Out4<11> ), .Out5(\Out5<11> ), .Out6(\Out6<11> ), .Out7(
        \Out7<11> ) );
  demux1to8_12 \demux[12]  ( .In(\In<12> ), .S({n5, \S<1> , n1}), .Out0(
        \Out0<12> ), .Out1(\Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ), 
        .Out4(\Out4<12> ), .Out5(\Out5<12> ), .Out6(\Out6<12> ), .Out7(
        \Out7<12> ) );
  demux1to8_13 \demux[13]  ( .In(\In<13> ), .S({n5, \S<1> , n1}), .Out0(
        \Out0<13> ), .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ), 
        .Out4(\Out4<13> ), .Out5(\Out5<13> ), .Out6(\Out6<13> ), .Out7(
        \Out7<13> ) );
  demux1to8_14 \demux[14]  ( .In(\In<14> ), .S({n5, n3, n1}), .Out0(\Out0<14> ), .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ), .Out4(\Out4<14> ), 
        .Out5(\Out5<14> ), .Out6(\Out6<14> ), .Out7(\Out7<14> ) );
  demux1to8_15 \demux[15]  ( .In(\In<15> ), .S({n5, \S<1> , n1}), .Out0(
        \Out0<15> ), .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ), 
        .Out4(\Out4<15> ), .Out5(\Out5<15> ), .Out6(\Out6<15> ), .Out7(
        \Out7<15> ) );
  INVX1 U1 ( .A(\S<2> ), .Y(n7) );
  INVX1 U2 ( .A(n7), .Y(n6) );
  INVX1 U3 ( .A(n4), .Y(n3) );
  INVX1 U4 ( .A(\S<0> ), .Y(n2) );
  INVX1 U5 ( .A(n7), .Y(n5) );
  INVX1 U6 ( .A(n2), .Y(n1) );
  INVX1 U7 ( .A(\S<1> ), .Y(n4) );
endmodule


module demux1to2_16_1 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), S, .Out0({\Out0<15> , \Out0<14> , 
        \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , \Out0<9> , \Out0<8> , 
        \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , \Out0<3> , \Out0<2> , 
        \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , \Out1<14> , \Out1<13> , 
        \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , \Out1<8> , \Out1<7> , 
        \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , \Out1<2> , \Out1<1> , 
        \Out1<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , S;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> ;


  demux1to2_17 \d[0]  ( .In(\In<0> ), .S(S), .Out0(\Out0<0> ), .Out1(\Out1<0> ) );
  demux1to2_18 \d[1]  ( .In(\In<1> ), .S(S), .Out0(\Out0<1> ), .Out1(\Out1<1> ) );
  demux1to2_19 \d[2]  ( .In(\In<2> ), .S(S), .Out0(\Out0<2> ), .Out1(\Out1<2> ) );
  demux1to2_20 \d[3]  ( .In(\In<3> ), .S(S), .Out0(\Out0<3> ), .Out1(\Out1<3> ) );
  demux1to2_21 \d[4]  ( .In(\In<4> ), .S(S), .Out0(\Out0<4> ), .Out1(\Out1<4> ) );
  demux1to2_22 \d[5]  ( .In(\In<5> ), .S(S), .Out0(\Out0<5> ), .Out1(\Out1<5> ) );
  demux1to2_23 \d[6]  ( .In(\In<6> ), .S(S), .Out0(\Out0<6> ), .Out1(\Out1<6> ) );
  demux1to2_24 \d[7]  ( .In(\In<7> ), .S(S), .Out0(\Out0<7> ), .Out1(\Out1<7> ) );
  demux1to2_25 \d[8]  ( .In(\In<8> ), .S(S), .Out0(\Out0<8> ), .Out1(\Out1<8> ) );
  demux1to2_26 \d[9]  ( .In(\In<9> ), .S(S), .Out0(\Out0<9> ), .Out1(\Out1<9> ) );
  demux1to2_27 \d[10]  ( .In(\In<10> ), .S(S), .Out0(\Out0<10> ), .Out1(
        \Out1<10> ) );
  demux1to2_28 \d[11]  ( .In(\In<11> ), .S(S), .Out0(\Out0<11> ), .Out1(
        \Out1<11> ) );
  demux1to2_29 \d[12]  ( .In(\In<12> ), .S(S), .Out0(\Out0<12> ), .Out1(
        \Out1<12> ) );
  demux1to2_30 \d[13]  ( .In(\In<13> ), .S(S), .Out0(\Out0<13> ), .Out1(
        \Out1<13> ) );
  demux1to2_31 \d[14]  ( .In(\In<14> ), .S(S), .Out0(\Out0<14> ), .Out1(
        \Out1<14> ) );
  demux1to2_32 \d[15]  ( .In(\In<15> ), .S(S), .Out0(\Out0<15> ), .Out1(
        \Out1<15> ) );
endmodule


module demux1to2_16_0 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), S, .Out0({\Out0<15> , \Out0<14> , 
        \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , \Out0<9> , \Out0<8> , 
        \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , \Out0<3> , \Out0<2> , 
        \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , \Out1<14> , \Out1<13> , 
        \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , \Out1<8> , \Out1<7> , 
        \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , \Out1<2> , \Out1<1> , 
        \Out1<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , S;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> ;


  demux1to2_15 \d[0]  ( .In(\In<0> ), .S(S), .Out0(\Out0<0> ), .Out1(\Out1<0> ) );
  demux1to2_14 \d[1]  ( .In(\In<1> ), .S(S), .Out0(\Out0<1> ), .Out1(\Out1<1> ) );
  demux1to2_13 \d[2]  ( .In(\In<2> ), .S(S), .Out0(\Out0<2> ), .Out1(\Out1<2> ) );
  demux1to2_12 \d[3]  ( .In(\In<3> ), .S(S), .Out0(\Out0<3> ), .Out1(\Out1<3> ) );
  demux1to2_11 \d[4]  ( .In(\In<4> ), .S(S), .Out0(\Out0<4> ), .Out1(\Out1<4> ) );
  demux1to2_10 \d[5]  ( .In(\In<5> ), .S(S), .Out0(\Out0<5> ), .Out1(\Out1<5> ) );
  demux1to2_9 \d[6]  ( .In(\In<6> ), .S(S), .Out0(\Out0<6> ), .Out1(\Out1<6> )
         );
  demux1to2_8 \d[7]  ( .In(\In<7> ), .S(S), .Out0(\Out0<7> ), .Out1(\Out1<7> )
         );
  demux1to2_7 \d[8]  ( .In(\In<8> ), .S(S), .Out0(\Out0<8> ), .Out1(\Out1<8> )
         );
  demux1to2_6 \d[9]  ( .In(\In<9> ), .S(S), .Out0(\Out0<9> ), .Out1(\Out1<9> )
         );
  demux1to2_5 \d[10]  ( .In(\In<10> ), .S(S), .Out0(\Out0<10> ), .Out1(
        \Out1<10> ) );
  demux1to2_4 \d[11]  ( .In(\In<11> ), .S(S), .Out0(\Out0<11> ), .Out1(
        \Out1<11> ) );
  demux1to2_3 \d[12]  ( .In(\In<12> ), .S(S), .Out0(\Out0<12> ), .Out1(
        \Out1<12> ) );
  demux1to2_2 \d[13]  ( .In(\In<13> ), .S(S), .Out0(\Out0<13> ), .Out1(
        \Out1<13> ) );
  demux1to2_1 \d[14]  ( .In(\In<14> ), .S(S), .Out0(\Out0<14> ), .Out1(
        \Out1<14> ) );
  demux1to2_0 \d[15]  ( .In(\In<15> ), .S(S), .Out0(\Out0<15> ), .Out1(
        \Out1<15> ) );
endmodule


module cla_or_xor_and ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , 
        \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , 
        \B<3> , \B<2> , \B<1> , \B<0> }), Cin, .Op({\Op<1> , \Op<0> }), .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<1> , \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Cout;
  wire   cla_cout, \op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> ,
         \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> ,
         \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> ,
         \op0_A<1> , \op0_A<0> , \op1_A<15> , \op1_A<14> , \op1_A<13> ,
         \op1_A<12> , \op1_A<11> , \op1_A<10> , \op1_A<9> , \op1_A<8> ,
         \op1_A<7> , \op1_A<6> , \op1_A<5> , \op1_A<4> , \op1_A<3> ,
         \op1_A<2> , \op1_A<1> , \op1_A<0> , \op2_A<15> , \op2_A<14> ,
         \op2_A<13> , \op2_A<12> , \op2_A<11> , \op2_A<10> , \op2_A<9> ,
         \op2_A<8> , \op2_A<7> , \op2_A<6> , \op2_A<5> , \op2_A<4> ,
         \op2_A<3> , \op2_A<2> , \op2_A<1> , \op2_A<0> , \op3_A<15> ,
         \op3_A<14> , \op3_A<13> , \op3_A<12> , \op3_A<11> , \op3_A<10> ,
         \op3_A<9> , \op3_A<8> , \op3_A<7> , \op3_A<6> , \op3_A<5> ,
         \op3_A<4> , \op3_A<3> , \op3_A<2> , \op3_A<1> , \op3_A<0> ,
         \op0_B<15> , \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> ,
         \op0_B<10> , \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> ,
         \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , \op0_B<1> ,
         \op0_B<0> , \op1_B<15> , \op1_B<14> , \op1_B<13> , \op1_B<12> ,
         \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , \op1_B<7> ,
         \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> ,
         \op1_B<1> , \op1_B<0> , \op2_B<15> , \op2_B<14> , \op2_B<13> ,
         \op2_B<12> , \op2_B<11> , \op2_B<10> , \op2_B<9> , \op2_B<8> ,
         \op2_B<7> , \op2_B<6> , \op2_B<5> , \op2_B<4> , \op2_B<3> ,
         \op2_B<2> , \op2_B<1> , \op2_B<0> , \op3_B<15> , \op3_B<14> ,
         \op3_B<13> , \op3_B<12> , \op3_B<11> , \op3_B<10> , \op3_B<9> ,
         \op3_B<8> , \op3_B<7> , \op3_B<6> , \op3_B<5> , \op3_B<4> ,
         \op3_B<3> , \op3_B<2> , \op3_B<1> , \op3_B<0> , \op0_out<15> ,
         \op0_out<14> , \op0_out<13> , \op0_out<12> , \op0_out<11> ,
         \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , \op0_out<6> ,
         \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , \op0_out<1> ,
         \op0_out<0> , \op2_out<15> , \op2_out<14> , \op2_out<13> ,
         \op2_out<12> , \op2_out<11> , \op2_out<10> , \op2_out<9> ,
         \op2_out<8> , \op2_out<7> , \op2_out<6> , \op2_out<5> , \op2_out<4> ,
         \op2_out<3> , \op2_out<2> , \op2_out<1> , \op2_out<0> , \op3_out<15> ,
         \op3_out<14> , \op3_out<13> , \op3_out<12> , \op3_out<11> ,
         \op3_out<10> , \op3_out<9> , \op3_out<8> , \op3_out<7> , \op3_out<6> ,
         \op3_out<5> , \op3_out<4> , \op3_out<3> , \op3_out<2> , \op3_out<1> ,
         \op3_out<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;

  demux1to4_16_1 demux0 ( .In({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .S({\Op<1> , \Op<0> }), .Out0({\op0_A<15> , 
        \op0_A<14> , \op0_A<13> , \op0_A<12> , \op0_A<11> , \op0_A<10> , 
        \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , \op0_A<5> , \op0_A<4> , 
        \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .Out1({\op1_A<15> , 
        \op1_A<14> , \op1_A<13> , \op1_A<12> , \op1_A<11> , \op1_A<10> , 
        \op1_A<9> , \op1_A<8> , \op1_A<7> , \op1_A<6> , \op1_A<5> , \op1_A<4> , 
        \op1_A<3> , \op1_A<2> , \op1_A<1> , \op1_A<0> }), .Out2({\op2_A<15> , 
        \op2_A<14> , \op2_A<13> , \op2_A<12> , \op2_A<11> , \op2_A<10> , 
        \op2_A<9> , \op2_A<8> , \op2_A<7> , \op2_A<6> , \op2_A<5> , \op2_A<4> , 
        \op2_A<3> , \op2_A<2> , \op2_A<1> , \op2_A<0> }), .Out3({\op3_A<15> , 
        \op3_A<14> , \op3_A<13> , \op3_A<12> , \op3_A<11> , \op3_A<10> , 
        \op3_A<9> , \op3_A<8> , \op3_A<7> , \op3_A<6> , \op3_A<5> , \op3_A<4> , 
        \op3_A<3> , \op3_A<2> , \op3_A<1> , \op3_A<0> }) );
  demux1to4_16_0 demux1 ( .In({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , 
        \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , 
        \B<2> , \B<1> , \B<0> }), .S({\Op<1> , \Op<0> }), .Out0({\op0_B<15> , 
        \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , \op0_B<10> , 
        \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , 
        \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }), .Out1({\op1_B<15> , 
        \op1_B<14> , \op1_B<13> , \op1_B<12> , \op1_B<11> , \op1_B<10> , 
        \op1_B<9> , \op1_B<8> , \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , 
        \op1_B<3> , \op1_B<2> , \op1_B<1> , \op1_B<0> }), .Out2({\op2_B<15> , 
        \op2_B<14> , \op2_B<13> , \op2_B<12> , \op2_B<11> , \op2_B<10> , 
        \op2_B<9> , \op2_B<8> , \op2_B<7> , \op2_B<6> , \op2_B<5> , \op2_B<4> , 
        \op2_B<3> , \op2_B<2> , \op2_B<1> , \op2_B<0> }), .Out3({\op3_B<15> , 
        \op3_B<14> , \op3_B<13> , \op3_B<12> , \op3_B<11> , \op3_B<10> , 
        \op3_B<9> , \op3_B<8> , \op3_B<7> , \op3_B<6> , \op3_B<5> , \op3_B<4> , 
        \op3_B<3> , \op3_B<2> , \op3_B<1> , \op3_B<0> }) );
  cla16_0 cla0 ( .A({\op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> , 
        \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> , 
        \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> , \op0_A<1> , 
        \op0_A<0> }), .B({\op0_B<15> , \op0_B<14> , \op0_B<13> , \op0_B<12> , 
        \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> , \op0_B<7> , 
        \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , \op0_B<1> , 
        \op0_B<0> }), .Cin(Cin), .S({\op0_out<15> , \op0_out<14> , 
        \op0_out<13> , \op0_out<12> , \op0_out<11> , \op0_out<10> , 
        \op0_out<9> , \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , 
        \op0_out<4> , \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> }), 
        .Cout(cla_cout) );
  mux4to1_16_0 mux0 ( .InA({\op0_out<15> , \op0_out<14> , \op0_out<13> , 
        \op0_out<12> , \op0_out<11> , \op0_out<10> , \op0_out<9> , 
        \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , \op0_out<4> , 
        \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> }), .InB({n29, 
        n27, n25, n23, n21, n19, n17, n15, n13, n31, n33, n11, n9, n7, n5, n3}), .InC({\op2_out<15> , \op2_out<14> , \op2_out<13> , \op2_out<12> , 
        \op2_out<11> , \op2_out<10> , \op2_out<9> , \op2_out<8> , \op2_out<7> , 
        \op2_out<6> , \op2_out<5> , \op2_out<4> , \op2_out<3> , \op2_out<2> , 
        \op2_out<1> , \op2_out<0> }), .InD({\op3_out<15> , \op3_out<14> , 
        \op3_out<13> , \op3_out<12> , \op3_out<11> , \op3_out<10> , 
        \op3_out<9> , \op3_out<8> , \op3_out<7> , \op3_out<6> , \op3_out<5> , 
        \op3_out<4> , \op3_out<3> , \op3_out<2> , \op3_out<1> , \op3_out<0> }), 
        .S({\Op<1> , n1}), .Out({\Out<15> , \Out<14> , \Out<13> , \Out<12> , 
        \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , 
        \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> }) );
  AND2X1 U2 ( .A(n67), .B(n66), .Y(n14) );
  AND2X1 U3 ( .A(n65), .B(n64), .Y(n12) );
  AND2X1 U4 ( .A(n61), .B(n60), .Y(n32) );
  BUFX2 U5 ( .A(\Op<0> ), .Y(n1) );
  AND2X2 U6 ( .A(n51), .B(n50), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  AND2X2 U8 ( .A(n53), .B(n52), .Y(n4) );
  INVX1 U9 ( .A(n4), .Y(n5) );
  AND2X2 U10 ( .A(n55), .B(n54), .Y(n6) );
  INVX1 U11 ( .A(n6), .Y(n7) );
  AND2X2 U12 ( .A(n57), .B(n56), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  AND2X2 U14 ( .A(n59), .B(n58), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  INVX1 U16 ( .A(n12), .Y(n13) );
  INVX1 U17 ( .A(n14), .Y(n15) );
  AND2X2 U18 ( .A(n69), .B(n68), .Y(n16) );
  INVX1 U19 ( .A(n16), .Y(n17) );
  AND2X2 U20 ( .A(n71), .B(n70), .Y(n18) );
  INVX1 U21 ( .A(n18), .Y(n19) );
  AND2X2 U22 ( .A(n73), .B(n72), .Y(n20) );
  INVX1 U23 ( .A(n20), .Y(n21) );
  AND2X2 U24 ( .A(n75), .B(n74), .Y(n22) );
  INVX1 U25 ( .A(n22), .Y(n23) );
  AND2X2 U26 ( .A(n77), .B(n76), .Y(n24) );
  INVX1 U27 ( .A(n24), .Y(n25) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  AND2X2 U30 ( .A(n81), .B(n80), .Y(n28) );
  INVX1 U31 ( .A(n28), .Y(n29) );
  AND2X2 U32 ( .A(n63), .B(n62), .Y(n30) );
  INVX1 U33 ( .A(n30), .Y(n31) );
  INVX1 U34 ( .A(cla_cout), .Y(n82) );
  INVX1 U35 ( .A(\op1_B<15> ), .Y(n81) );
  INVX1 U36 ( .A(\op1_B<14> ), .Y(n79) );
  INVX1 U37 ( .A(\op1_B<13> ), .Y(n77) );
  INVX1 U38 ( .A(\op1_B<12> ), .Y(n75) );
  INVX1 U39 ( .A(\op1_B<11> ), .Y(n73) );
  INVX1 U40 ( .A(\op1_B<10> ), .Y(n71) );
  INVX1 U41 ( .A(\op1_B<9> ), .Y(n69) );
  INVX1 U42 ( .A(\op1_B<7> ), .Y(n65) );
  INVX1 U43 ( .A(\op1_B<6> ), .Y(n63) );
  INVX1 U44 ( .A(\op1_B<5> ), .Y(n61) );
  INVX1 U45 ( .A(\op1_B<4> ), .Y(n59) );
  INVX1 U46 ( .A(\op1_B<3> ), .Y(n57) );
  INVX1 U47 ( .A(\op1_B<2> ), .Y(n55) );
  INVX1 U48 ( .A(\op1_B<1> ), .Y(n53) );
  INVX1 U49 ( .A(\op1_B<0> ), .Y(n51) );
  INVX1 U50 ( .A(\op2_A<15> ), .Y(n49) );
  INVX1 U51 ( .A(\op1_A<15> ), .Y(n80) );
  INVX1 U52 ( .A(\op2_A<14> ), .Y(n48) );
  INVX1 U53 ( .A(\op1_A<14> ), .Y(n78) );
  INVX1 U54 ( .A(\op2_A<13> ), .Y(n47) );
  INVX1 U55 ( .A(\op1_A<13> ), .Y(n76) );
  INVX1 U56 ( .A(\op2_A<12> ), .Y(n46) );
  INVX1 U57 ( .A(\op1_A<12> ), .Y(n74) );
  INVX1 U58 ( .A(\op2_A<11> ), .Y(n45) );
  INVX1 U59 ( .A(\op1_A<11> ), .Y(n72) );
  INVX1 U60 ( .A(\op2_A<10> ), .Y(n44) );
  INVX1 U61 ( .A(\op1_A<10> ), .Y(n70) );
  INVX1 U62 ( .A(\op2_A<9> ), .Y(n43) );
  INVX1 U63 ( .A(\op1_A<9> ), .Y(n68) );
  INVX1 U64 ( .A(\op2_A<8> ), .Y(n42) );
  INVX1 U65 ( .A(\op2_A<7> ), .Y(n41) );
  INVX1 U66 ( .A(\op1_A<7> ), .Y(n64) );
  INVX1 U67 ( .A(\op2_A<6> ), .Y(n40) );
  INVX1 U68 ( .A(\op1_A<6> ), .Y(n62) );
  INVX1 U69 ( .A(\op2_A<5> ), .Y(n39) );
  INVX1 U70 ( .A(\op1_A<5> ), .Y(n60) );
  INVX1 U71 ( .A(\op2_A<4> ), .Y(n38) );
  INVX1 U72 ( .A(\op1_A<4> ), .Y(n58) );
  INVX1 U73 ( .A(\op2_A<3> ), .Y(n37) );
  INVX1 U74 ( .A(\op1_A<3> ), .Y(n56) );
  INVX1 U75 ( .A(\op2_A<2> ), .Y(n36) );
  INVX1 U76 ( .A(\op1_A<2> ), .Y(n54) );
  INVX1 U77 ( .A(\op2_A<1> ), .Y(n35) );
  INVX1 U78 ( .A(\op1_A<1> ), .Y(n52) );
  INVX1 U79 ( .A(\op2_A<0> ), .Y(n34) );
  INVX1 U80 ( .A(\op1_A<0> ), .Y(n50) );
  INVX1 U81 ( .A(n32), .Y(n33) );
  INVX1 U82 ( .A(\op1_B<8> ), .Y(n67) );
  INVX1 U83 ( .A(\op1_A<8> ), .Y(n66) );
  AND2X2 U84 ( .A(\op3_A<0> ), .B(\op3_B<0> ), .Y(\op3_out<0> ) );
  AND2X2 U85 ( .A(\op3_A<1> ), .B(\op3_B<1> ), .Y(\op3_out<1> ) );
  AND2X2 U86 ( .A(\op3_A<2> ), .B(\op3_B<2> ), .Y(\op3_out<2> ) );
  AND2X2 U87 ( .A(\op3_A<3> ), .B(\op3_B<3> ), .Y(\op3_out<3> ) );
  AND2X2 U88 ( .A(\op3_A<4> ), .B(\op3_B<4> ), .Y(\op3_out<4> ) );
  AND2X2 U89 ( .A(\op3_A<5> ), .B(\op3_B<5> ), .Y(\op3_out<5> ) );
  AND2X2 U90 ( .A(\op3_A<6> ), .B(\op3_B<6> ), .Y(\op3_out<6> ) );
  AND2X2 U91 ( .A(\op3_A<7> ), .B(\op3_B<7> ), .Y(\op3_out<7> ) );
  AND2X2 U92 ( .A(\op3_A<8> ), .B(\op3_B<8> ), .Y(\op3_out<8> ) );
  AND2X2 U93 ( .A(\op3_A<9> ), .B(\op3_B<9> ), .Y(\op3_out<9> ) );
  AND2X2 U94 ( .A(\op3_A<10> ), .B(\op3_B<10> ), .Y(\op3_out<10> ) );
  AND2X2 U95 ( .A(\op3_A<11> ), .B(\op3_B<11> ), .Y(\op3_out<11> ) );
  AND2X2 U96 ( .A(\op3_A<12> ), .B(\op3_B<12> ), .Y(\op3_out<12> ) );
  AND2X2 U97 ( .A(\op3_A<13> ), .B(\op3_B<13> ), .Y(\op3_out<13> ) );
  AND2X2 U98 ( .A(\op3_A<14> ), .B(\op3_B<14> ), .Y(\op3_out<14> ) );
  AND2X2 U99 ( .A(\op3_A<15> ), .B(\op3_B<15> ), .Y(\op3_out<15> ) );
  XNOR2X1 U100 ( .A(\op2_B<0> ), .B(n34), .Y(\op2_out<0> ) );
  XNOR2X1 U101 ( .A(\op2_B<1> ), .B(n35), .Y(\op2_out<1> ) );
  XNOR2X1 U102 ( .A(\op2_B<2> ), .B(n36), .Y(\op2_out<2> ) );
  XNOR2X1 U103 ( .A(\op2_B<3> ), .B(n37), .Y(\op2_out<3> ) );
  XNOR2X1 U104 ( .A(\op2_B<4> ), .B(n38), .Y(\op2_out<4> ) );
  XNOR2X1 U105 ( .A(\op2_B<5> ), .B(n39), .Y(\op2_out<5> ) );
  XNOR2X1 U106 ( .A(\op2_B<6> ), .B(n40), .Y(\op2_out<6> ) );
  XNOR2X1 U107 ( .A(\op2_B<7> ), .B(n41), .Y(\op2_out<7> ) );
  XNOR2X1 U108 ( .A(\op2_B<8> ), .B(n42), .Y(\op2_out<8> ) );
  XNOR2X1 U109 ( .A(\op2_B<9> ), .B(n43), .Y(\op2_out<9> ) );
  XNOR2X1 U110 ( .A(\op2_B<10> ), .B(n44), .Y(\op2_out<10> ) );
  XNOR2X1 U111 ( .A(\op2_B<11> ), .B(n45), .Y(\op2_out<11> ) );
  XNOR2X1 U112 ( .A(\op2_B<12> ), .B(n46), .Y(\op2_out<12> ) );
  XNOR2X1 U113 ( .A(\op2_B<13> ), .B(n47), .Y(\op2_out<13> ) );
  XNOR2X1 U114 ( .A(\op2_B<14> ), .B(n48), .Y(\op2_out<14> ) );
  XNOR2X1 U115 ( .A(\op2_B<15> ), .B(n49), .Y(\op2_out<15> ) );
  NOR3X1 U116 ( .A(\Op<1> ), .B(n1), .C(n82), .Y(Cout) );
endmodule


module shifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Op({\Op<1> , \Op<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , \Op<1> ,
         \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \ls_out<15> , \ls_out<14> , \ls_out<13> , \ls_out<12> , \ls_out<11> ,
         \ls_out<10> , \ls_out<9> , \ls_out<8> , \ls_out<7> , \ls_out<6> ,
         \ls_out<5> , \ls_out<4> , \ls_out<3> , \ls_out<2> , \ls_out<1> ,
         \ls_out<0> , \rs_out<15> , \rs_out<14> , \rs_out<13> , \rs_out<12> ,
         \rs_out<11> , \rs_out<10> , \rs_out<9> , \rs_out<8> , \rs_out<7> ,
         \rs_out<6> , \rs_out<5> , \rs_out<4> , \rs_out<3> , \rs_out<2> ,
         \rs_out<1> , \rs_out<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;

  lshifter ls ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Rot_sel(n2), .Out({\ls_out<15> , \ls_out<14> , 
        \ls_out<13> , \ls_out<12> , \ls_out<11> , \ls_out<10> , \ls_out<9> , 
        \ls_out<8> , \ls_out<7> , \ls_out<6> , \ls_out<5> , \ls_out<4> , 
        \ls_out<3> , \ls_out<2> , \ls_out<1> , \ls_out<0> }) );
  rshifter rs ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Rot_sel(n2), .Out({\rs_out<15> , \rs_out<14> , 
        \rs_out<13> , \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> , 
        \rs_out<8> , \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> , 
        \rs_out<3> , \rs_out<2> , \rs_out<1> , \rs_out<0> }) );
  INVX1 U1 ( .A(n1), .Y(\Out<1> ) );
  INVX1 U2 ( .A(\rs_out<2> ), .Y(n7) );
  INVX1 U3 ( .A(\rs_out<3> ), .Y(n9) );
  INVX1 U4 ( .A(\rs_out<9> ), .Y(n21) );
  INVX1 U5 ( .A(\rs_out<10> ), .Y(n23) );
  INVX1 U6 ( .A(\rs_out<11> ), .Y(n25) );
  INVX1 U7 ( .A(\rs_out<13> ), .Y(n29) );
  INVX1 U8 ( .A(\rs_out<14> ), .Y(n31) );
  INVX1 U9 ( .A(\rs_out<15> ), .Y(n33) );
  INVX1 U10 ( .A(\ls_out<5> ), .Y(n14) );
  INVX1 U11 ( .A(\ls_out<9> ), .Y(n22) );
  INVX1 U12 ( .A(\ls_out<13> ), .Y(n30) );
  INVX1 U13 ( .A(\rs_out<0> ), .Y(n5) );
  INVX1 U14 ( .A(\rs_out<5> ), .Y(n13) );
  INVX1 U15 ( .A(\rs_out<6> ), .Y(n15) );
  INVX1 U16 ( .A(\rs_out<7> ), .Y(n17) );
  INVX1 U17 ( .A(\rs_out<8> ), .Y(n19) );
  INVX1 U18 ( .A(\rs_out<12> ), .Y(n27) );
  INVX1 U19 ( .A(\ls_out<0> ), .Y(n6) );
  INVX1 U20 ( .A(\ls_out<2> ), .Y(n8) );
  INVX1 U21 ( .A(\ls_out<3> ), .Y(n10) );
  INVX1 U22 ( .A(\ls_out<6> ), .Y(n16) );
  INVX1 U23 ( .A(\ls_out<7> ), .Y(n18) );
  INVX1 U24 ( .A(\ls_out<8> ), .Y(n20) );
  INVX1 U25 ( .A(\ls_out<10> ), .Y(n24) );
  INVX1 U26 ( .A(\ls_out<11> ), .Y(n26) );
  INVX1 U27 ( .A(\ls_out<12> ), .Y(n28) );
  INVX1 U28 ( .A(\ls_out<14> ), .Y(n32) );
  INVX1 U29 ( .A(\ls_out<15> ), .Y(n34) );
  MUX2X1 U30 ( .B(\ls_out<1> ), .A(\rs_out<1> ), .S(\Op<1> ), .Y(n1) );
  INVX1 U31 ( .A(\rs_out<4> ), .Y(n11) );
  INVX1 U32 ( .A(\ls_out<4> ), .Y(n12) );
  INVX2 U33 ( .A(\Op<1> ), .Y(n4) );
  INVX1 U34 ( .A(\Op<0> ), .Y(n2) );
  INVX8 U35 ( .A(n4), .Y(n3) );
  MUX2X1 U36 ( .B(n6), .A(n5), .S(n3), .Y(\Out<0> ) );
  MUX2X1 U37 ( .B(n8), .A(n7), .S(n3), .Y(\Out<2> ) );
  MUX2X1 U38 ( .B(n10), .A(n9), .S(n3), .Y(\Out<3> ) );
  MUX2X1 U39 ( .B(n12), .A(n11), .S(n3), .Y(\Out<4> ) );
  MUX2X1 U40 ( .B(n14), .A(n13), .S(n3), .Y(\Out<5> ) );
  MUX2X1 U41 ( .B(n16), .A(n15), .S(n3), .Y(\Out<6> ) );
  MUX2X1 U42 ( .B(n18), .A(n17), .S(n3), .Y(\Out<7> ) );
  MUX2X1 U43 ( .B(n20), .A(n19), .S(n3), .Y(\Out<8> ) );
  MUX2X1 U44 ( .B(n22), .A(n21), .S(n3), .Y(\Out<9> ) );
  MUX2X1 U45 ( .B(n24), .A(n23), .S(n3), .Y(\Out<10> ) );
  MUX2X1 U46 ( .B(n26), .A(n25), .S(n3), .Y(\Out<11> ) );
  MUX2X1 U47 ( .B(n28), .A(n27), .S(n3), .Y(\Out<12> ) );
  MUX2X1 U48 ( .B(n30), .A(n29), .S(n3), .Y(\Out<13> ) );
  MUX2X1 U49 ( .B(n32), .A(n31), .S(n3), .Y(\Out<14> ) );
  MUX2X1 U50 ( .B(n34), .A(n33), .S(n3), .Y(\Out<15> ) );
endmodule


module cla4_7 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;

  fulladder1_31 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n42), .G(n38) );
  fulladder1_30 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n17), .S(\S<1> ), .P(
        n43), .G(n39) );
  fulladder1_29 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n37), .S(\S<2> ), .P(
        n44), .G(n40) );
  fulladder1_28 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n36), .S(\S<3> ), .P(
        n45), .G(n41) );
  INVX1 U1 ( .A(n33), .Y(n20) );
  INVX1 U2 ( .A(n36), .Y(n35) );
  AND2X2 U3 ( .A(n44), .B(n23), .Y(n1) );
  AND2X2 U4 ( .A(n43), .B(n22), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(n3) );
  AND2X2 U6 ( .A(n45), .B(n30), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n5) );
  AND2X2 U8 ( .A(n43), .B(n22), .Y(n6) );
  BUFX2 U9 ( .A(n21), .Y(n7) );
  BUFX2 U10 ( .A(n31), .Y(n8) );
  AND2X2 U11 ( .A(n45), .B(n30), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(n10) );
  BUFX2 U13 ( .A(n32), .Y(n11) );
  BUFX2 U14 ( .A(n25), .Y(n12) );
  BUFX2 U15 ( .A(n34), .Y(n13) );
  INVX1 U16 ( .A(n28), .Y(n14) );
  INVX1 U17 ( .A(n27), .Y(n28) );
  BUFX2 U18 ( .A(n26), .Y(n15) );
  INVX1 U19 ( .A(n1), .Y(n16) );
  INVX1 U20 ( .A(n18), .Y(n17) );
  AND2X2 U21 ( .A(n7), .B(n15), .Y(n18) );
  INVX1 U22 ( .A(n6), .Y(n19) );
  XNOR2X1 U23 ( .A(\A<0> ), .B(\B<0> ), .Y(n33) );
  NAND3X1 U24 ( .A(Cin), .B(n42), .C(n20), .Y(n21) );
  NAND3X1 U25 ( .A(\A<0> ), .B(\B<0> ), .C(n38), .Y(n26) );
  XOR2X1 U26 ( .A(\A<1> ), .B(\B<1> ), .Y(n22) );
  NAND3X1 U27 ( .A(\A<1> ), .B(\B<1> ), .C(n39), .Y(n25) );
  OAI21X1 U28 ( .A(n19), .B(n18), .C(n12), .Y(n37) );
  XOR2X1 U29 ( .A(\A<2> ), .B(\B<2> ), .Y(n23) );
  INVX2 U30 ( .A(n37), .Y(n24) );
  NAND3X1 U31 ( .A(\A<2> ), .B(\B<2> ), .C(n40), .Y(n27) );
  OAI21X1 U32 ( .A(n16), .B(n24), .C(n14), .Y(n36) );
  OAI21X1 U33 ( .A(n3), .B(n15), .C(n12), .Y(n29) );
  AOI21X1 U34 ( .A(n1), .B(n29), .C(n28), .Y(n31) );
  XOR2X1 U35 ( .A(\A<3> ), .B(\B<3> ), .Y(n30) );
  NAND3X1 U36 ( .A(\A<3> ), .B(\B<3> ), .C(n41), .Y(n34) );
  OAI21X1 U37 ( .A(n8), .B(n10), .C(n13), .Y(GG) );
  NAND3X1 U38 ( .A(n42), .B(n6), .C(n1), .Y(n32) );
  NOR3X1 U39 ( .A(n33), .B(n11), .C(n5), .Y(PG) );
  OAI21X1 U40 ( .A(n10), .B(n35), .C(n13), .Y(Cout) );
endmodule


module cla4_6 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  fulladder1_27 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n41), .G(n37) );
  fulladder1_26 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n9), .S(\S<1> ), .P(n42), .G(n38) );
  fulladder1_25 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n36), .S(\S<2> ), .P(
        n43), .G(n39) );
  fulladder1_24 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n35), .S(\S<3> ), .P(
        n44), .G(n40) );
  INVX1 U1 ( .A(n32), .Y(n18) );
  INVX1 U2 ( .A(n35), .Y(n34) );
  AND2X2 U3 ( .A(n42), .B(n20), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X2 U5 ( .A(n43), .B(n21), .Y(n3) );
  BUFX2 U6 ( .A(n19), .Y(n4) );
  AND2X2 U7 ( .A(n44), .B(n28), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  INVX1 U9 ( .A(n5), .Y(n7) );
  AND2X2 U10 ( .A(n4), .B(n15), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  BUFX2 U12 ( .A(n29), .Y(n10) );
  BUFX2 U13 ( .A(n31), .Y(n11) );
  BUFX2 U14 ( .A(n23), .Y(n12) );
  BUFX2 U15 ( .A(n33), .Y(n13) );
  INVX1 U16 ( .A(n26), .Y(n14) );
  INVX1 U17 ( .A(n25), .Y(n26) );
  BUFX2 U18 ( .A(n24), .Y(n15) );
  INVX1 U19 ( .A(n3), .Y(n16) );
  INVX1 U20 ( .A(n30), .Y(n17) );
  INVX1 U21 ( .A(n2), .Y(n30) );
  XNOR2X1 U22 ( .A(\A<0> ), .B(\B<0> ), .Y(n32) );
  NAND3X1 U23 ( .A(Cin), .B(n41), .C(n18), .Y(n19) );
  NAND3X1 U24 ( .A(\A<0> ), .B(\B<0> ), .C(n37), .Y(n24) );
  XOR2X1 U25 ( .A(\A<1> ), .B(\B<1> ), .Y(n20) );
  NAND3X1 U26 ( .A(\A<1> ), .B(\B<1> ), .C(n38), .Y(n23) );
  OAI21X1 U27 ( .A(n17), .B(n8), .C(n12), .Y(n36) );
  XOR2X1 U28 ( .A(\A<2> ), .B(\B<2> ), .Y(n21) );
  INVX2 U29 ( .A(n36), .Y(n22) );
  NAND3X1 U30 ( .A(\A<2> ), .B(\B<2> ), .C(n39), .Y(n25) );
  OAI21X1 U31 ( .A(n16), .B(n22), .C(n14), .Y(n35) );
  OAI21X1 U32 ( .A(n2), .B(n15), .C(n12), .Y(n27) );
  AOI21X1 U33 ( .A(n3), .B(n27), .C(n26), .Y(n29) );
  XOR2X1 U34 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  NAND3X1 U35 ( .A(\A<3> ), .B(\B<3> ), .C(n40), .Y(n33) );
  OAI21X1 U36 ( .A(n10), .B(n6), .C(n13), .Y(GG) );
  NAND3X1 U37 ( .A(n41), .B(n30), .C(n3), .Y(n31) );
  NOR3X1 U38 ( .A(n32), .B(n11), .C(n7), .Y(PG) );
  OAI21X1 U39 ( .A(n7), .B(n34), .C(n13), .Y(Cout) );
endmodule


module cla4_5 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;

  fulladder1_23 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n42), .G(n38) );
  fulladder1_22 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n9), .S(\S<1> ), .P(n43), .G(n39) );
  fulladder1_21 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n37), .S(\S<2> ), .P(
        n44), .G(n40) );
  fulladder1_20 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n36), .S(\S<3> ), .P(
        n45), .G(n41) );
  INVX1 U1 ( .A(n33), .Y(n20) );
  INVX1 U2 ( .A(n36), .Y(n35) );
  AND2X2 U3 ( .A(n43), .B(n22), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X2 U5 ( .A(n44), .B(n23), .Y(n3) );
  BUFX2 U6 ( .A(n21), .Y(n4) );
  AND2X2 U7 ( .A(n45), .B(n30), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  INVX1 U9 ( .A(n5), .Y(n7) );
  AND2X2 U10 ( .A(n4), .B(n17), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  INVX1 U12 ( .A(n31), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(n11) );
  INVX1 U14 ( .A(n32), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(n13) );
  BUFX2 U16 ( .A(n25), .Y(n14) );
  BUFX2 U17 ( .A(n34), .Y(n15) );
  INVX1 U18 ( .A(n28), .Y(n16) );
  INVX1 U19 ( .A(n27), .Y(n28) );
  BUFX2 U20 ( .A(n26), .Y(n17) );
  INVX1 U21 ( .A(n3), .Y(n18) );
  INVX1 U22 ( .A(n1), .Y(n19) );
  XNOR2X1 U23 ( .A(\A<0> ), .B(\B<0> ), .Y(n33) );
  NAND3X1 U24 ( .A(Cin), .B(n42), .C(n20), .Y(n21) );
  NAND3X1 U25 ( .A(\A<0> ), .B(\B<0> ), .C(n38), .Y(n26) );
  XOR2X1 U26 ( .A(\A<1> ), .B(\B<1> ), .Y(n22) );
  NAND3X1 U27 ( .A(\A<1> ), .B(\B<1> ), .C(n39), .Y(n25) );
  OAI21X1 U28 ( .A(n19), .B(n8), .C(n14), .Y(n37) );
  XOR2X1 U29 ( .A(\A<2> ), .B(\B<2> ), .Y(n23) );
  INVX2 U30 ( .A(n37), .Y(n24) );
  NAND3X1 U31 ( .A(\A<2> ), .B(\B<2> ), .C(n40), .Y(n27) );
  OAI21X1 U32 ( .A(n18), .B(n24), .C(n16), .Y(n36) );
  OAI21X1 U33 ( .A(n2), .B(n17), .C(n14), .Y(n29) );
  AOI21X1 U34 ( .A(n3), .B(n29), .C(n28), .Y(n31) );
  XOR2X1 U35 ( .A(\A<3> ), .B(\B<3> ), .Y(n30) );
  NAND3X1 U36 ( .A(\A<3> ), .B(\B<3> ), .C(n41), .Y(n34) );
  OAI21X1 U37 ( .A(n11), .B(n6), .C(n15), .Y(GG) );
  NAND3X1 U38 ( .A(n42), .B(n1), .C(n3), .Y(n32) );
  NOR3X1 U39 ( .A(n33), .B(n13), .C(n7), .Y(PG) );
  OAI21X1 U40 ( .A(n7), .B(n35), .C(n15), .Y(Cout) );
endmodule


module cla4_4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n50, \P<3> , \G<3> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49;

  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n43) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n48) );
  fulladder1_19 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n45), .G(n40) );
  fulladder1_18 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n4), .S(\S<1> ), .P(n46), .G(n41) );
  fulladder1_17 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n37), .S(\S<2> ), .P(
        n47), .G(n42) );
  fulladder1_16 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n36), .S(\S<3> ), .P(
        n49), .G(n44) );
  XOR2X1 U1 ( .A(\A<0> ), .B(\B<0> ), .Y(n1) );
  INVX1 U2 ( .A(n29), .Y(n35) );
  INVX1 U3 ( .A(n19), .Y(n34) );
  INVX1 U4 ( .A(\G<3> ), .Y(n38) );
  OR2X1 U5 ( .A(n8), .B(n10), .Y(n12) );
  INVX1 U6 ( .A(\P<3> ), .Y(n39) );
  BUFX2 U7 ( .A(n25), .Y(n2) );
  AND2X2 U8 ( .A(n2), .B(n20), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(n4) );
  AND2X2 U10 ( .A(\P<3> ), .B(n36), .Y(n5) );
  INVX1 U11 ( .A(n5), .Y(n6) );
  AND2X2 U12 ( .A(n1), .B(n23), .Y(n7) );
  INVX1 U13 ( .A(n7), .Y(n8) );
  AND2X2 U14 ( .A(n45), .B(n35), .Y(n9) );
  INVX1 U15 ( .A(n9), .Y(n10) );
  BUFX2 U16 ( .A(n50), .Y(GG) );
  INVX1 U17 ( .A(n12), .Y(PG) );
  AND2X1 U18 ( .A(n35), .B(n32), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(n15) );
  AND2X1 U20 ( .A(\P<3> ), .B(n34), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  BUFX2 U22 ( .A(n30), .Y(n18) );
  BUFX2 U23 ( .A(n33), .Y(n19) );
  BUFX2 U24 ( .A(n31), .Y(n20) );
  AND2X2 U25 ( .A(n47), .B(n27), .Y(n21) );
  INVX1 U26 ( .A(n21), .Y(n22) );
  AND2X2 U27 ( .A(n46), .B(n26), .Y(n23) );
  INVX1 U28 ( .A(n23), .Y(n24) );
  NAND3X1 U29 ( .A(n45), .B(n1), .C(Cin), .Y(n25) );
  NAND3X1 U30 ( .A(\A<0> ), .B(\B<0> ), .C(n40), .Y(n31) );
  XOR2X1 U31 ( .A(\A<1> ), .B(\B<1> ), .Y(n26) );
  NAND3X1 U32 ( .A(\A<1> ), .B(\B<1> ), .C(n41), .Y(n30) );
  OAI21X1 U33 ( .A(n24), .B(n3), .C(n18), .Y(n37) );
  XOR2X1 U34 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  INVX2 U35 ( .A(n37), .Y(n28) );
  NAND3X1 U36 ( .A(\A<2> ), .B(\B<2> ), .C(n42), .Y(n33) );
  OAI21X1 U37 ( .A(n22), .B(n28), .C(n19), .Y(n36) );
  OR2X2 U38 ( .A(n22), .B(n39), .Y(n29) );
  OAI21X1 U39 ( .A(n24), .B(n20), .C(n18), .Y(n32) );
  NAND3X1 U40 ( .A(n38), .B(n15), .C(n17), .Y(n50) );
  NAND2X1 U41 ( .A(n38), .B(n6), .Y(Cout) );
  AND2X1 U42 ( .A(n48), .B(n49), .Y(\P<3> ) );
  AND2X1 U43 ( .A(n43), .B(n44), .Y(\G<3> ) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memory2c_1 ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, n5053, n5054, n5055, \mem<0><7> ,
         \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><7> , \mem<1><6> , \mem<1><5> ,
         \mem<1><4> , \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> ,
         \mem<2><7> , \mem<2><6> , \mem<2><5> , \mem<2><4> , \mem<2><3> ,
         \mem<2><2> , \mem<2><1> , \mem<2><0> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><7> , \mem<4><6> , \mem<4><5> , \mem<4><4> ,
         \mem<4><3> , \mem<4><2> , \mem<4><1> , \mem<4><0> , \mem<5><7> ,
         \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><7> , \mem<6><6> , \mem<6><5> ,
         \mem<6><4> , \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> ,
         \mem<7><7> , \mem<7><6> , \mem<7><5> , \mem<7><4> , \mem<7><3> ,
         \mem<7><2> , \mem<7><1> , \mem<7><0> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><7> , \mem<9><6> , \mem<9><5> , \mem<9><4> ,
         \mem<9><3> , \mem<9><2> , \mem<9><1> , \mem<9><0> , \mem<10><7> ,
         \mem<10><6> , \mem<10><5> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><7> , \mem<11><6> , \mem<11><5> ,
         \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> , \mem<11><0> ,
         \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> , \mem<12><3> ,
         \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><7> ,
         \mem<15><6> , \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><7> , \mem<16><6> , \mem<16><5> ,
         \mem<16><4> , \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> ,
         \mem<17><7> , \mem<17><6> , \mem<17><5> , \mem<17><4> , \mem<17><3> ,
         \mem<17><2> , \mem<17><1> , \mem<17><0> , \mem<18><7> , \mem<18><6> ,
         \mem<18><5> , \mem<18><4> , \mem<18><3> , \mem<18><2> , \mem<18><1> ,
         \mem<18><0> , \mem<19><7> , \mem<19><6> , \mem<19><5> , \mem<19><4> ,
         \mem<19><3> , \mem<19><2> , \mem<19><1> , \mem<19><0> , \mem<20><7> ,
         \mem<20><6> , \mem<20><5> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><7> , \mem<21><6> , \mem<21><5> ,
         \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> , \mem<21><0> ,
         \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> , \mem<22><3> ,
         \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><7> ,
         \mem<25><6> , \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><7> , \mem<26><6> , \mem<26><5> ,
         \mem<26><4> , \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> ,
         \mem<27><7> , \mem<27><6> , \mem<27><5> , \mem<27><4> , \mem<27><3> ,
         \mem<27><2> , \mem<27><1> , \mem<27><0> , \mem<28><7> , \mem<28><6> ,
         \mem<28><5> , \mem<28><4> , \mem<28><3> , \mem<28><2> , \mem<28><1> ,
         \mem<28><0> , \mem<29><7> , \mem<29><6> , \mem<29><5> , \mem<29><4> ,
         \mem<29><3> , \mem<29><2> , \mem<29><1> , \mem<29><0> , \mem<30><7> ,
         \mem<30><6> , \mem<30><5> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><7> , \mem<31><6> , \mem<31><5> ,
         \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> , \mem<31><0> ,
         \mem<32><7> , \mem<32><6> , \mem<32><5> , \mem<32><4> , \mem<32><3> ,
         \mem<32><2> , \mem<32><1> , \mem<32><0> , \mem<33><7> , \mem<33><6> ,
         \mem<33><5> , \mem<33><4> , \mem<33><3> , \mem<33><2> , \mem<33><1> ,
         \mem<33><0> , \mem<34><7> , \mem<34><6> , \mem<34><5> , \mem<34><4> ,
         \mem<34><3> , \mem<34><2> , \mem<34><1> , \mem<34><0> , \mem<35><7> ,
         \mem<35><6> , \mem<35><5> , \mem<35><4> , \mem<35><3> , \mem<35><2> ,
         \mem<35><1> , \mem<35><0> , \mem<36><7> , \mem<36><6> , \mem<36><5> ,
         \mem<36><4> , \mem<36><3> , \mem<36><2> , \mem<36><1> , \mem<36><0> ,
         \mem<37><7> , \mem<37><6> , \mem<37><5> , \mem<37><4> , \mem<37><3> ,
         \mem<37><2> , \mem<37><1> , \mem<37><0> , \mem<38><7> , \mem<38><6> ,
         \mem<38><5> , \mem<38><4> , \mem<38><3> , \mem<38><2> , \mem<38><1> ,
         \mem<38><0> , \mem<39><7> , \mem<39><6> , \mem<39><5> , \mem<39><4> ,
         \mem<39><3> , \mem<39><2> , \mem<39><1> , \mem<39><0> , \mem<40><7> ,
         \mem<40><6> , \mem<40><5> , \mem<40><4> , \mem<40><3> , \mem<40><2> ,
         \mem<40><1> , \mem<40><0> , \mem<41><7> , \mem<41><6> , \mem<41><5> ,
         \mem<41><4> , \mem<41><3> , \mem<41><2> , \mem<41><1> , \mem<41><0> ,
         \mem<42><7> , \mem<42><6> , \mem<42><5> , \mem<42><4> , \mem<42><3> ,
         \mem<42><2> , \mem<42><1> , \mem<42><0> , \mem<43><7> , \mem<43><6> ,
         \mem<43><5> , \mem<43><4> , \mem<43><3> , \mem<43><2> , \mem<43><1> ,
         \mem<43><0> , \mem<44><7> , \mem<44><6> , \mem<44><5> , \mem<44><4> ,
         \mem<44><3> , \mem<44><2> , \mem<44><1> , \mem<44><0> , \mem<45><7> ,
         \mem<45><6> , \mem<45><5> , \mem<45><4> , \mem<45><3> , \mem<45><2> ,
         \mem<45><1> , \mem<45><0> , \mem<46><7> , \mem<46><6> , \mem<46><5> ,
         \mem<46><4> , \mem<46><3> , \mem<46><2> , \mem<46><1> , \mem<46><0> ,
         \mem<47><7> , \mem<47><6> , \mem<47><5> , \mem<47><4> , \mem<47><3> ,
         \mem<47><2> , \mem<47><1> , \mem<47><0> , \mem<48><7> , \mem<48><6> ,
         \mem<48><5> , \mem<48><4> , \mem<48><3> , \mem<48><2> , \mem<48><1> ,
         \mem<48><0> , \mem<49><7> , \mem<49><6> , \mem<49><5> , \mem<49><4> ,
         \mem<49><3> , \mem<49><2> , \mem<49><1> , \mem<49><0> , \mem<50><7> ,
         \mem<50><6> , \mem<50><5> , \mem<50><4> , \mem<50><3> , \mem<50><2> ,
         \mem<50><1> , \mem<50><0> , \mem<51><7> , \mem<51><6> , \mem<51><5> ,
         \mem<51><4> , \mem<51><3> , \mem<51><2> , \mem<51><1> , \mem<51><0> ,
         \mem<52><7> , \mem<52><6> , \mem<52><5> , \mem<52><4> , \mem<52><3> ,
         \mem<52><2> , \mem<52><1> , \mem<52><0> , \mem<53><7> , \mem<53><6> ,
         \mem<53><5> , \mem<53><4> , \mem<53><3> , \mem<53><2> , \mem<53><1> ,
         \mem<53><0> , \mem<54><7> , \mem<54><6> , \mem<54><5> , \mem<54><4> ,
         \mem<54><3> , \mem<54><2> , \mem<54><1> , \mem<54><0> , \mem<55><7> ,
         \mem<55><6> , \mem<55><5> , \mem<55><4> , \mem<55><3> , \mem<55><2> ,
         \mem<55><1> , \mem<55><0> , \mem<56><7> , \mem<56><6> , \mem<56><5> ,
         \mem<56><4> , \mem<56><3> , \mem<56><2> , \mem<56><1> , \mem<56><0> ,
         \mem<57><7> , \mem<57><6> , \mem<57><5> , \mem<57><4> , \mem<57><3> ,
         \mem<57><2> , \mem<57><1> , \mem<57><0> , \mem<58><7> , \mem<58><6> ,
         \mem<58><5> , \mem<58><4> , \mem<58><3> , \mem<58><2> , \mem<58><1> ,
         \mem<58><0> , \mem<59><7> , \mem<59><6> , \mem<59><5> , \mem<59><4> ,
         \mem<59><3> , \mem<59><2> , \mem<59><1> , \mem<59><0> , \mem<60><7> ,
         \mem<60><6> , \mem<60><5> , \mem<60><4> , \mem<60><3> , \mem<60><2> ,
         \mem<60><1> , \mem<60><0> , \mem<61><7> , \mem<61><6> , \mem<61><5> ,
         \mem<61><4> , \mem<61><3> , \mem<61><2> , \mem<61><1> , \mem<61><0> ,
         \mem<62><7> , \mem<62><6> , \mem<62><5> , \mem<62><4> , \mem<62><3> ,
         \mem<62><2> , \mem<62><1> , \mem<62><0> , \mem<63><7> , \mem<63><6> ,
         \mem<63><5> , \mem<63><4> , \mem<63><3> , \mem<63><2> , \mem<63><1> ,
         \mem<63><0> , N185, N186, N187, N188, N189, N190, N191, N192, n599,
         n602, n603, n604, n605, n606, n607, n608, n625, n1525, n1526, n1527,
         n1552, n1577, n1578, n1579, n1604, n1629, n1630, n1631, n1656, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n600, n601, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n2327), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2326), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2325), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2324), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2323), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2322), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2321), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2320), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2319), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2318), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2317), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2316), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2315), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2314), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2313), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2312), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2311), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2310), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2309), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2308), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2307), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2306), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2305), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2304), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2303), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2302), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2301), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2300), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2299), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2298), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2297), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2296), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2295), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2294), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2293), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2292), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2291), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2290), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2289), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2288), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2287), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2286), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2285), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2284), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2283), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2282), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2281), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2280), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2279), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2278), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2277), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2276), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2275), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2274), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2273), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2272), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2271), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2270), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2269), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2268), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2267), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2266), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2265), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2264), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2263), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2262), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2261), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2260), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2259), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2258), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2257), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2256), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2255), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2254), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2253), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2252), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2251), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2250), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2249), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2248), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2247), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2246), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2245), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2244), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2243), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2242), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2241), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2240), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2239), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2238), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2237), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2236), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2235), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2234), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2233), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2232), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2231), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2230), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2229), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2228), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2227), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2226), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2225), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2224), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2223), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2222), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2221), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2220), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2219), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2218), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2217), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2216), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2215), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2214), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2213), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2212), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2211), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2210), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2209), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2208), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2207), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2206), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2205), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2204), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2203), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2202), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2201), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2200), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2199), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2198), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2197), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2196), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2195), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2194), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2193), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2192), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2191), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2190), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2189), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2188), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2187), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2186), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2185), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2184), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2183), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2182), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2181), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2180), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2179), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2178), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2177), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2176), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2175), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2174), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2173), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2172), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2171), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2170), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2169), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2168), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2167), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2166), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2165), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2164), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2163), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2162), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2161), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2160), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2159), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2158), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2157), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2156), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2155), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2154), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2153), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2152), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2151), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2150), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2149), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2148), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2147), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2146), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2145), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2144), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2143), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2142), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2141), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2140), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2139), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2138), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2137), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2136), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2135), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2134), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2133), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2132), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2131), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2130), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2129), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2128), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2127), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2126), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2125), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2124), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2123), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2122), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2121), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2120), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2119), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2118), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2117), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2116), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2115), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2114), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2113), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2112), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2111), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2110), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2109), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2108), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2107), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2106), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2105), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2104), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2103), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2102), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2101), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2100), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2099), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2098), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2097), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2096), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2095), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2094), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2093), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2092), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2091), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2090), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2089), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2088), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2087), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2086), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2085), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2084), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2083), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2082), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2081), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2080), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2079), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2078), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2077), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2076), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2075), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2074), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2073), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2072), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n2071), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n2070), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n2069), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n2068), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n2067), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n2066), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n2065), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n2064), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n2063), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n2062), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n2061), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n2060), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n2059), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n2058), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n2057), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n2056), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n2055), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n2054), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n2053), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n2052), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n2051), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n2050), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n2049), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n2048), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n2047), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n2046), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n2045), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n2044), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n2043), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n2042), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n2041), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n2040), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n2039), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n2038), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n2037), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n2036), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n2035), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n2034), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n2033), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n2032), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n2031), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n2030), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n2029), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n2028), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n2027), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n2026), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n2025), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n2024), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n2023), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n2022), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n2021), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n2020), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n2019), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n2018), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n2017), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n2016), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n2015), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n2014), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n2013), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n2012), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n2011), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n2010), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n2009), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n2008), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n2007), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n2006), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n2005), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n2004), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n2003), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n2002), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n2001), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n2000), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n1999), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n1998), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n1997), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n1996), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n1995), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n1994), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n1993), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n1992), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n1991), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n1990), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n1989), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n1988), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n1987), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n1986), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n1985), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n1984), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n1983), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n1982), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n1981), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n1980), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n1979), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n1978), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n1977), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n1976), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n1975), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n1974), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n1973), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n1972), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n1971), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n1970), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n1969), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n1968), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n1967), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n1966), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n1965), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n1964), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n1963), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n1962), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n1961), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n1960), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n1959), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n1958), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n1957), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n1956), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n1955), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n1954), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n1953), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n1952), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n1951), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n1950), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n1949), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n1948), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n1947), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n1946), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n1945), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n1944), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n1943), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n1942), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n1941), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n1940), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n1939), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n1938), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n1937), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n1936), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n1935), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n1934), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n1933), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n1932), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n1931), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n1930), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n1929), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n1928), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n1927), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n1926), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n1925), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n1924), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n1923), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n1922), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n1921), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n1920), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n1919), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n1918), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n1917), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n1916), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n1915), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n1914), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n1913), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n1912), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n1911), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n1910), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n1909), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n1908), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n1907), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n1906), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n1905), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n1904), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n1903), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n1902), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n1901), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n1900), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n1899), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n1898), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n1897), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n1896), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n1895), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n1894), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n1893), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n1892), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n1891), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n1890), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n1889), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n1888), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n1887), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n1886), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n1885), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n1884), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n1883), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n1882), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n1881), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n1880), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n1879), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n1878), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n1877), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n1876), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n1875), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n1874), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n1873), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n1872), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n1871), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n1870), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n1869), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n1868), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n1867), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n1866), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n1865), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n1864), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n1863), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n1862), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n1861), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n1860), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n1859), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n1858), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n1857), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n1856), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n1855), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n1854), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n1853), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n1852), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n1851), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n1850), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n1849), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n1848), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n1847), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n1846), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n1845), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n1844), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n1843), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n1842), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n1841), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n1840), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n1839), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n1838), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n1837), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n1836), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n1835), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n1834), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n1833), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n1832), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n1831), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n1830), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n1829), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n1828), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n1827), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n1826), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n1825), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n1824), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n1823), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n1822), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n1821), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n1820), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n1819), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n1818), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n1817), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n1816), .CLK(clk), .Q(\mem<63><0> ) );
  OAI21X1 U817 ( .A(n4586), .B(n2684), .C(n809), .Y(n1816) );
  OAI21X1 U819 ( .A(n4586), .B(n2747), .C(n808), .Y(n1817) );
  OAI21X1 U821 ( .A(n4586), .B(n5052), .C(n807), .Y(n1818) );
  OAI21X1 U823 ( .A(n4586), .B(n5051), .C(n806), .Y(n1819) );
  OAI21X1 U825 ( .A(n4586), .B(n5050), .C(n805), .Y(n1820) );
  OAI21X1 U827 ( .A(n4586), .B(n5049), .C(n804), .Y(n1821) );
  OAI21X1 U829 ( .A(n4586), .B(n5048), .C(n803), .Y(n1822) );
  OAI21X1 U831 ( .A(n4586), .B(n2882), .C(n802), .Y(n1823) );
  NAND3X1 U1905 ( .A(enable), .B(n2637), .C(wr), .Y(n625) );
  AOI21X1 U2035 ( .A(n1525), .B(n1526), .C(n2623), .Y(n5053) );
  NOR3X1 U2036 ( .A(n1527), .B(n1150), .C(n1164), .Y(n1526) );
  NOR3X1 U2057 ( .A(n1552), .B(n1148), .C(n1162), .Y(n1525) );
  AOI21X1 U2078 ( .A(n1577), .B(n1578), .C(n2623), .Y(n5054) );
  NOR3X1 U2079 ( .A(n1579), .B(n1146), .C(n1160), .Y(n1578) );
  NOR3X1 U2100 ( .A(n1604), .B(n1144), .C(n1158), .Y(n1577) );
  AOI21X1 U2121 ( .A(n1629), .B(n1630), .C(n2623), .Y(n5055) );
  NOR3X1 U2122 ( .A(n1631), .B(n1142), .C(n1156), .Y(n1630) );
  NOR3X1 U2143 ( .A(n1656), .B(n1140), .C(n1154), .Y(n1629) );
  INVX1 U3 ( .A(n70), .Y(n1) );
  INVX1 U4 ( .A(n532), .Y(n2) );
  INVX4 U5 ( .A(n416), .Y(n3849) );
  INVX1 U6 ( .A(n3290), .Y(n3267) );
  INVX1 U7 ( .A(n3370), .Y(n3348) );
  INVX1 U8 ( .A(n3214), .Y(n3192) );
  INVX1 U9 ( .A(n3316), .Y(n3294) );
  INVX1 U10 ( .A(n3344), .Y(n3321) );
  AND2X1 U11 ( .A(n2629), .B(n719), .Y(n1193) );
  AND2X1 U12 ( .A(n1445), .B(\mem<35><6> ), .Y(n138) );
  INVX2 U13 ( .A(n2635), .Y(n2634) );
  AND2X1 U14 ( .A(n2624), .B(n444), .Y(n700) );
  AND2X1 U15 ( .A(n2628), .B(n703), .Y(n1177) );
  AND2X1 U16 ( .A(n3167), .B(n444), .Y(n702) );
  AND2X1 U17 ( .A(n2628), .B(n709), .Y(n1183) );
  AND2X1 U18 ( .A(n2628), .B(n713), .Y(n1187) );
  AND2X1 U19 ( .A(n2629), .B(n715), .Y(n1189) );
  AND2X1 U20 ( .A(n2629), .B(n727), .Y(n1201) );
  INVX1 U21 ( .A(n446), .Y(n3953) );
  AND2X1 U22 ( .A(n2631), .B(n775), .Y(n1249) );
  AND2X1 U23 ( .A(n2631), .B(n777), .Y(n1251) );
  AND2X1 U24 ( .A(n2631), .B(n779), .Y(n1253) );
  INVX1 U25 ( .A(n2963), .Y(n4586) );
  OR2X1 U26 ( .A(n1034), .B(n1048), .Y(n1132) );
  INVX1 U27 ( .A(\mem<62><0> ), .Y(n5047) );
  INVX1 U28 ( .A(\mem<62><1> ), .Y(n5046) );
  INVX1 U29 ( .A(\mem<62><7> ), .Y(n5042) );
  INVX1 U30 ( .A(\mem<61><2> ), .Y(n5041) );
  INVX1 U31 ( .A(\mem<61><3> ), .Y(n5040) );
  INVX1 U32 ( .A(\mem<61><4> ), .Y(n5039) );
  INVX1 U33 ( .A(\mem<61><5> ), .Y(n5038) );
  INVX1 U34 ( .A(\mem<61><6> ), .Y(n5037) );
  INVX1 U35 ( .A(\mem<60><0> ), .Y(n5036) );
  INVX1 U36 ( .A(\mem<60><1> ), .Y(n5035) );
  INVX1 U37 ( .A(\mem<60><7> ), .Y(n5031) );
  INVX1 U38 ( .A(\mem<59><0> ), .Y(n5030) );
  INVX1 U39 ( .A(\mem<59><2> ), .Y(n5029) );
  INVX1 U40 ( .A(\mem<59><3> ), .Y(n5028) );
  INVX1 U41 ( .A(\mem<59><4> ), .Y(n5027) );
  INVX1 U42 ( .A(\mem<59><5> ), .Y(n5026) );
  INVX1 U43 ( .A(\mem<59><6> ), .Y(n5025) );
  INVX1 U44 ( .A(\mem<58><0> ), .Y(n5024) );
  INVX1 U45 ( .A(\mem<58><1> ), .Y(n5023) );
  INVX1 U46 ( .A(\mem<58><5> ), .Y(n2783) );
  INVX1 U47 ( .A(\mem<58><6> ), .Y(n5019) );
  INVX1 U48 ( .A(\mem<58><7> ), .Y(n5018) );
  INVX1 U49 ( .A(\mem<57><0> ), .Y(n5017) );
  INVX1 U50 ( .A(\mem<57><1> ), .Y(n5016) );
  INVX1 U51 ( .A(\mem<57><7> ), .Y(n5012) );
  INVX1 U52 ( .A(\mem<56><0> ), .Y(n5011) );
  INVX1 U53 ( .A(\mem<56><1> ), .Y(n5010) );
  INVX1 U54 ( .A(\mem<56><2> ), .Y(n5009) );
  INVX1 U55 ( .A(\mem<56><3> ), .Y(n5008) );
  INVX1 U56 ( .A(\mem<56><4> ), .Y(n5007) );
  INVX1 U57 ( .A(\mem<56><5> ), .Y(n5006) );
  INVX1 U58 ( .A(\mem<56><6> ), .Y(n5005) );
  INVX1 U59 ( .A(\mem<56><7> ), .Y(n5004) );
  INVX1 U60 ( .A(\mem<55><0> ), .Y(n5003) );
  INVX1 U61 ( .A(\mem<55><1> ), .Y(n5002) );
  INVX1 U62 ( .A(\mem<55><2> ), .Y(n5001) );
  INVX1 U63 ( .A(\mem<55><3> ), .Y(n5000) );
  INVX1 U64 ( .A(\mem<55><4> ), .Y(n4999) );
  INVX1 U65 ( .A(\mem<55><5> ), .Y(n4998) );
  INVX1 U66 ( .A(\mem<55><6> ), .Y(n4997) );
  INVX1 U67 ( .A(\mem<55><7> ), .Y(n4996) );
  INVX1 U68 ( .A(\mem<54><0> ), .Y(n4995) );
  INVX1 U69 ( .A(\mem<54><1> ), .Y(n4994) );
  INVX1 U70 ( .A(\mem<54><5> ), .Y(n4990) );
  INVX1 U71 ( .A(\mem<54><6> ), .Y(n4989) );
  INVX1 U72 ( .A(\mem<54><7> ), .Y(n4988) );
  AND2X1 U73 ( .A(n514), .B(n1179), .Y(n1320) );
  INVX1 U74 ( .A(\mem<53><0> ), .Y(n4987) );
  INVX1 U75 ( .A(\mem<53><1> ), .Y(n4986) );
  INVX1 U76 ( .A(\mem<53><2> ), .Y(n4985) );
  INVX1 U77 ( .A(\mem<53><3> ), .Y(n4984) );
  INVX1 U78 ( .A(\mem<53><4> ), .Y(n4983) );
  INVX1 U79 ( .A(\mem<53><5> ), .Y(n4982) );
  INVX1 U80 ( .A(\mem<53><6> ), .Y(n4981) );
  INVX1 U81 ( .A(\mem<53><7> ), .Y(n4980) );
  AND2X1 U82 ( .A(n482), .B(n1181), .Y(n1322) );
  INVX1 U83 ( .A(\mem<52><0> ), .Y(n4979) );
  INVX1 U84 ( .A(\mem<52><1> ), .Y(n4978) );
  INVX1 U85 ( .A(\mem<52><5> ), .Y(n4974) );
  INVX1 U86 ( .A(\mem<52><6> ), .Y(n4973) );
  INVX1 U87 ( .A(\mem<52><7> ), .Y(n4972) );
  AND2X1 U88 ( .A(n506), .B(n3267), .Y(n1324) );
  INVX1 U89 ( .A(\mem<51><0> ), .Y(n4971) );
  INVX1 U90 ( .A(\mem<51><1> ), .Y(n4970) );
  INVX1 U91 ( .A(\mem<51><2> ), .Y(n4969) );
  INVX1 U92 ( .A(\mem<51><3> ), .Y(n4968) );
  INVX1 U93 ( .A(\mem<51><4> ), .Y(n4967) );
  INVX1 U94 ( .A(\mem<51><5> ), .Y(n4966) );
  INVX1 U95 ( .A(\mem<51><6> ), .Y(n4965) );
  INVX1 U96 ( .A(\mem<51><7> ), .Y(n4964) );
  INVX1 U97 ( .A(\mem<50><0> ), .Y(n4963) );
  INVX1 U98 ( .A(\mem<50><1> ), .Y(n4962) );
  INVX1 U99 ( .A(\mem<50><5> ), .Y(n4958) );
  INVX1 U100 ( .A(\mem<50><6> ), .Y(n4957) );
  INVX1 U101 ( .A(\mem<50><7> ), .Y(n4956) );
  INVX1 U102 ( .A(\mem<49><0> ), .Y(n4955) );
  INVX1 U103 ( .A(\mem<49><1> ), .Y(n4954) );
  INVX1 U104 ( .A(\mem<49><2> ), .Y(n4953) );
  INVX1 U105 ( .A(\mem<49><3> ), .Y(n4952) );
  INVX1 U106 ( .A(\mem<49><4> ), .Y(n4951) );
  INVX1 U107 ( .A(\mem<49><5> ), .Y(n4950) );
  INVX1 U108 ( .A(\mem<49><6> ), .Y(n4949) );
  INVX1 U109 ( .A(\mem<49><7> ), .Y(n4948) );
  AND2X1 U110 ( .A(n440), .B(n3348), .Y(n1330) );
  INVX1 U111 ( .A(\mem<48><0> ), .Y(n4947) );
  INVX1 U112 ( .A(\mem<48><1> ), .Y(n4946) );
  INVX1 U113 ( .A(\mem<48><5> ), .Y(n4942) );
  INVX1 U114 ( .A(\mem<48><6> ), .Y(n4941) );
  INVX1 U115 ( .A(\mem<48><7> ), .Y(n4940) );
  INVX1 U116 ( .A(\mem<47><0> ), .Y(n4939) );
  INVX1 U117 ( .A(\mem<47><1> ), .Y(n4938) );
  INVX1 U118 ( .A(\mem<47><2> ), .Y(n4937) );
  INVX1 U119 ( .A(\mem<47><3> ), .Y(n4936) );
  INVX1 U120 ( .A(\mem<47><4> ), .Y(n4935) );
  INVX1 U121 ( .A(\mem<47><5> ), .Y(n4934) );
  INVX1 U122 ( .A(\mem<47><6> ), .Y(n4933) );
  INVX1 U123 ( .A(\mem<47><7> ), .Y(n4932) );
  INVX1 U124 ( .A(\mem<46><0> ), .Y(n4931) );
  INVX1 U125 ( .A(\mem<46><1> ), .Y(n4930) );
  INVX1 U126 ( .A(\mem<46><5> ), .Y(n4926) );
  INVX1 U127 ( .A(\mem<46><6> ), .Y(n4925) );
  INVX1 U128 ( .A(\mem<46><7> ), .Y(n4924) );
  INVX1 U129 ( .A(\mem<45><0> ), .Y(n4923) );
  INVX1 U130 ( .A(\mem<45><1> ), .Y(n4922) );
  INVX1 U131 ( .A(\mem<45><2> ), .Y(n4921) );
  INVX1 U132 ( .A(\mem<45><3> ), .Y(n4920) );
  INVX1 U133 ( .A(\mem<45><4> ), .Y(n4919) );
  INVX1 U134 ( .A(\mem<45><5> ), .Y(n4918) );
  INVX1 U135 ( .A(\mem<45><6> ), .Y(n4917) );
  INVX1 U136 ( .A(\mem<45><7> ), .Y(n4916) );
  INVX1 U137 ( .A(\mem<44><0> ), .Y(n4915) );
  INVX1 U138 ( .A(\mem<44><1> ), .Y(n4914) );
  INVX1 U139 ( .A(\mem<44><5> ), .Y(n4910) );
  INVX1 U140 ( .A(\mem<44><6> ), .Y(n4909) );
  INVX1 U141 ( .A(\mem<44><7> ), .Y(n4908) );
  AND2X1 U142 ( .A(n2613), .B(n1191), .Y(n1340) );
  INVX1 U143 ( .A(\mem<43><0> ), .Y(n4907) );
  INVX1 U144 ( .A(\mem<43><1> ), .Y(n4906) );
  INVX1 U145 ( .A(\mem<43><2> ), .Y(n4905) );
  INVX1 U146 ( .A(\mem<43><3> ), .Y(n4904) );
  INVX1 U147 ( .A(\mem<43><4> ), .Y(n4903) );
  INVX1 U148 ( .A(\mem<43><6> ), .Y(n4901) );
  INVX1 U149 ( .A(\mem<43><7> ), .Y(n4900) );
  AND2X1 U150 ( .A(n17), .B(n1193), .Y(n1342) );
  INVX1 U151 ( .A(\mem<42><0> ), .Y(n4899) );
  INVX1 U152 ( .A(\mem<42><1> ), .Y(n4898) );
  INVX1 U153 ( .A(\mem<42><6> ), .Y(n4893) );
  INVX1 U154 ( .A(\mem<42><7> ), .Y(n4892) );
  INVX1 U155 ( .A(\mem<41><0> ), .Y(n4891) );
  INVX1 U156 ( .A(\mem<41><1> ), .Y(n4890) );
  INVX1 U157 ( .A(\mem<41><5> ), .Y(n4886) );
  INVX1 U158 ( .A(\mem<41><6> ), .Y(n4885) );
  INVX1 U159 ( .A(\mem<41><7> ), .Y(n4884) );
  AND2X1 U160 ( .A(n7), .B(n1197), .Y(n1346) );
  INVX1 U161 ( .A(\mem<40><0> ), .Y(n4883) );
  INVX1 U162 ( .A(\mem<40><1> ), .Y(n4882) );
  INVX1 U163 ( .A(\mem<40><2> ), .Y(n4881) );
  INVX1 U164 ( .A(\mem<40><3> ), .Y(n4880) );
  INVX1 U165 ( .A(\mem<40><4> ), .Y(n4879) );
  INVX1 U166 ( .A(\mem<40><5> ), .Y(n4878) );
  INVX1 U167 ( .A(\mem<40><6> ), .Y(n4877) );
  INVX1 U168 ( .A(\mem<40><7> ), .Y(n4876) );
  AND2X1 U169 ( .A(n483), .B(n1199), .Y(n1348) );
  INVX1 U170 ( .A(\mem<39><0> ), .Y(n4875) );
  INVX1 U171 ( .A(\mem<39><1> ), .Y(n4874) );
  INVX1 U172 ( .A(\mem<39><2> ), .Y(n4873) );
  INVX1 U173 ( .A(\mem<39><4> ), .Y(n4872) );
  INVX1 U174 ( .A(\mem<39><6> ), .Y(n4870) );
  INVX1 U175 ( .A(\mem<39><7> ), .Y(n4869) );
  INVX1 U176 ( .A(\mem<38><0> ), .Y(n4868) );
  INVX1 U177 ( .A(\mem<38><1> ), .Y(n4867) );
  INVX1 U178 ( .A(\mem<38><6> ), .Y(n4863) );
  INVX1 U179 ( .A(\mem<38><7> ), .Y(n4862) );
  INVX1 U180 ( .A(\mem<37><0> ), .Y(n4861) );
  INVX1 U181 ( .A(\mem<37><1> ), .Y(n4860) );
  INVX1 U182 ( .A(\mem<37><2> ), .Y(n4859) );
  INVX1 U183 ( .A(\mem<37><3> ), .Y(n4858) );
  INVX1 U184 ( .A(\mem<37><4> ), .Y(n4857) );
  INVX1 U185 ( .A(\mem<37><5> ), .Y(n4856) );
  INVX1 U186 ( .A(\mem<37><6> ), .Y(n4855) );
  INVX1 U187 ( .A(\mem<37><7> ), .Y(n4854) );
  INVX1 U188 ( .A(\mem<36><0> ), .Y(n4853) );
  INVX1 U189 ( .A(\mem<36><1> ), .Y(n4852) );
  INVX1 U190 ( .A(\mem<36><5> ), .Y(n4848) );
  INVX1 U191 ( .A(\mem<36><6> ), .Y(n4847) );
  INVX1 U192 ( .A(\mem<36><7> ), .Y(n4846) );
  INVX1 U193 ( .A(\mem<35><0> ), .Y(n4845) );
  INVX1 U194 ( .A(\mem<35><2> ), .Y(n4843) );
  INVX1 U195 ( .A(\mem<35><3> ), .Y(n4842) );
  INVX1 U196 ( .A(\mem<35><4> ), .Y(n4841) );
  INVX1 U197 ( .A(\mem<35><5> ), .Y(n4840) );
  INVX1 U198 ( .A(\mem<35><6> ), .Y(n4839) );
  INVX1 U199 ( .A(\mem<35><7> ), .Y(n4838) );
  INVX1 U200 ( .A(\mem<34><0> ), .Y(n4837) );
  INVX1 U201 ( .A(\mem<34><5> ), .Y(n4832) );
  INVX1 U202 ( .A(\mem<34><6> ), .Y(n4831) );
  INVX1 U203 ( .A(\mem<34><7> ), .Y(n4830) );
  INVX1 U204 ( .A(\mem<33><0> ), .Y(n4829) );
  INVX1 U205 ( .A(\mem<33><1> ), .Y(n4828) );
  INVX1 U206 ( .A(\mem<33><2> ), .Y(n4827) );
  INVX1 U207 ( .A(\mem<33><3> ), .Y(n4826) );
  INVX1 U208 ( .A(\mem<33><4> ), .Y(n4825) );
  INVX1 U209 ( .A(\mem<33><5> ), .Y(n4824) );
  INVX1 U210 ( .A(\mem<33><6> ), .Y(n4823) );
  INVX1 U211 ( .A(\mem<33><7> ), .Y(n4822) );
  INVX1 U212 ( .A(\mem<32><5> ), .Y(n4818) );
  INVX1 U213 ( .A(\mem<32><6> ), .Y(n4817) );
  AND2X1 U214 ( .A(n539), .B(n1215), .Y(n1364) );
  INVX1 U215 ( .A(\mem<31><0> ), .Y(n4816) );
  INVX1 U216 ( .A(\mem<31><1> ), .Y(n4815) );
  INVX1 U217 ( .A(\mem<31><2> ), .Y(n4814) );
  INVX1 U218 ( .A(\mem<31><3> ), .Y(n4813) );
  INVX1 U219 ( .A(\mem<31><4> ), .Y(n4812) );
  INVX1 U220 ( .A(\mem<31><5> ), .Y(n4811) );
  INVX1 U221 ( .A(\mem<31><6> ), .Y(n4810) );
  INVX1 U222 ( .A(\mem<31><7> ), .Y(n4809) );
  AND2X1 U223 ( .A(n433), .B(n1217), .Y(n1366) );
  INVX1 U224 ( .A(\mem<30><0> ), .Y(n4808) );
  INVX1 U225 ( .A(\mem<30><1> ), .Y(n4807) );
  INVX1 U226 ( .A(\mem<30><5> ), .Y(n4803) );
  INVX1 U227 ( .A(\mem<30><6> ), .Y(n4802) );
  INVX1 U228 ( .A(\mem<30><7> ), .Y(n4801) );
  INVX1 U229 ( .A(\mem<29><0> ), .Y(n4800) );
  INVX1 U230 ( .A(\mem<29><1> ), .Y(n4799) );
  INVX1 U231 ( .A(\mem<29><2> ), .Y(n4798) );
  INVX1 U232 ( .A(\mem<29><3> ), .Y(n4797) );
  INVX1 U233 ( .A(\mem<29><4> ), .Y(n4796) );
  INVX1 U234 ( .A(\mem<29><7> ), .Y(n4795) );
  INVX1 U235 ( .A(\mem<28><1> ), .Y(n4794) );
  INVX1 U236 ( .A(\mem<28><5> ), .Y(n4790) );
  INVX1 U237 ( .A(\mem<28><6> ), .Y(n4789) );
  INVX1 U238 ( .A(\mem<27><0> ), .Y(n4788) );
  INVX1 U239 ( .A(\mem<27><1> ), .Y(n4787) );
  INVX1 U240 ( .A(\mem<27><2> ), .Y(n4786) );
  INVX1 U241 ( .A(\mem<27><3> ), .Y(n4785) );
  INVX1 U242 ( .A(\mem<27><4> ), .Y(n4784) );
  INVX1 U243 ( .A(\mem<27><7> ), .Y(n4783) );
  INVX1 U244 ( .A(\mem<26><5> ), .Y(n4779) );
  INVX1 U245 ( .A(\mem<26><6> ), .Y(n4778) );
  INVX1 U246 ( .A(\mem<25><5> ), .Y(n4774) );
  INVX1 U247 ( .A(\mem<25><6> ), .Y(n4773) );
  INVX1 U248 ( .A(\mem<24><0> ), .Y(n4772) );
  INVX1 U249 ( .A(\mem<24><1> ), .Y(n4771) );
  INVX1 U250 ( .A(\mem<24><2> ), .Y(n4770) );
  INVX1 U251 ( .A(\mem<24><3> ), .Y(n4769) );
  INVX1 U252 ( .A(\mem<24><4> ), .Y(n4768) );
  INVX1 U253 ( .A(\mem<24><5> ), .Y(n4767) );
  INVX1 U254 ( .A(\mem<24><6> ), .Y(n4766) );
  INVX1 U255 ( .A(\mem<24><7> ), .Y(n4765) );
  AND2X1 U256 ( .A(n465), .B(n1231), .Y(n1380) );
  INVX1 U257 ( .A(\mem<23><0> ), .Y(n4764) );
  INVX1 U258 ( .A(\mem<23><1> ), .Y(n4763) );
  INVX1 U259 ( .A(\mem<23><2> ), .Y(n4762) );
  INVX1 U260 ( .A(\mem<23><3> ), .Y(n4761) );
  INVX1 U261 ( .A(\mem<23><4> ), .Y(n4760) );
  INVX1 U262 ( .A(\mem<23><5> ), .Y(n4759) );
  INVX1 U263 ( .A(\mem<23><6> ), .Y(n4758) );
  INVX1 U264 ( .A(\mem<23><7> ), .Y(n4757) );
  INVX1 U265 ( .A(\mem<22><0> ), .Y(n4756) );
  INVX1 U266 ( .A(\mem<22><1> ), .Y(n4755) );
  INVX1 U267 ( .A(\mem<22><5> ), .Y(n4751) );
  INVX1 U268 ( .A(\mem<22><6> ), .Y(n4750) );
  INVX1 U269 ( .A(\mem<22><7> ), .Y(n4749) );
  INVX1 U270 ( .A(\mem<21><0> ), .Y(n4748) );
  INVX1 U271 ( .A(\mem<21><1> ), .Y(n4747) );
  INVX1 U272 ( .A(\mem<21><2> ), .Y(n4746) );
  INVX1 U273 ( .A(\mem<21><3> ), .Y(n4745) );
  INVX1 U274 ( .A(\mem<21><4> ), .Y(n4744) );
  INVX1 U275 ( .A(\mem<21><5> ), .Y(n4743) );
  INVX1 U276 ( .A(\mem<21><6> ), .Y(n4742) );
  INVX1 U277 ( .A(\mem<21><7> ), .Y(n4741) );
  AND2X1 U278 ( .A(n461), .B(n1237), .Y(n1386) );
  INVX1 U279 ( .A(\mem<20><0> ), .Y(n4740) );
  INVX1 U280 ( .A(\mem<20><1> ), .Y(n4739) );
  INVX1 U281 ( .A(\mem<20><5> ), .Y(n4735) );
  INVX1 U282 ( .A(\mem<20><6> ), .Y(n4734) );
  INVX1 U283 ( .A(\mem<20><7> ), .Y(n4733) );
  INVX1 U284 ( .A(\mem<19><0> ), .Y(n4732) );
  INVX1 U285 ( .A(\mem<19><1> ), .Y(n4731) );
  INVX1 U286 ( .A(\mem<19><2> ), .Y(n4730) );
  INVX1 U287 ( .A(\mem<19><3> ), .Y(n4729) );
  INVX1 U288 ( .A(\mem<19><4> ), .Y(n4728) );
  INVX1 U289 ( .A(\mem<19><5> ), .Y(n4727) );
  INVX1 U290 ( .A(\mem<19><6> ), .Y(n4726) );
  INVX1 U291 ( .A(\mem<19><7> ), .Y(n4725) );
  AND2X1 U292 ( .A(n566), .B(n1241), .Y(n1390) );
  INVX1 U293 ( .A(\mem<18><0> ), .Y(n4724) );
  INVX1 U294 ( .A(\mem<18><1> ), .Y(n4723) );
  INVX1 U295 ( .A(\mem<18><5> ), .Y(n4719) );
  INVX1 U296 ( .A(\mem<18><6> ), .Y(n4718) );
  INVX1 U297 ( .A(\mem<18><7> ), .Y(n4717) );
  INVX1 U298 ( .A(\mem<17><0> ), .Y(n4716) );
  INVX1 U299 ( .A(\mem<17><1> ), .Y(n4715) );
  INVX1 U300 ( .A(\mem<17><2> ), .Y(n4714) );
  INVX1 U301 ( .A(\mem<17><3> ), .Y(n4713) );
  INVX1 U302 ( .A(\mem<17><4> ), .Y(n4712) );
  INVX1 U303 ( .A(\mem<17><5> ), .Y(n4711) );
  INVX1 U304 ( .A(\mem<17><6> ), .Y(n4710) );
  INVX1 U305 ( .A(\mem<17><7> ), .Y(n4709) );
  AND2X1 U306 ( .A(n77), .B(n1245), .Y(n1394) );
  INVX1 U307 ( .A(\mem<16><0> ), .Y(n4708) );
  INVX1 U308 ( .A(\mem<16><1> ), .Y(n4707) );
  INVX1 U309 ( .A(\mem<16><5> ), .Y(n4703) );
  INVX1 U310 ( .A(\mem<16><6> ), .Y(n4702) );
  INVX1 U311 ( .A(\mem<16><7> ), .Y(n4701) );
  INVX1 U312 ( .A(\mem<15><0> ), .Y(n4700) );
  INVX1 U313 ( .A(\mem<15><1> ), .Y(n4699) );
  INVX1 U314 ( .A(\mem<15><2> ), .Y(n4698) );
  INVX1 U315 ( .A(\mem<15><3> ), .Y(n4697) );
  INVX1 U316 ( .A(\mem<15><4> ), .Y(n4696) );
  INVX1 U317 ( .A(\mem<15><5> ), .Y(n4695) );
  INVX1 U318 ( .A(\mem<15><6> ), .Y(n4694) );
  INVX1 U319 ( .A(\mem<15><7> ), .Y(n4693) );
  INVX1 U320 ( .A(\mem<14><0> ), .Y(n4692) );
  INVX1 U321 ( .A(\mem<14><1> ), .Y(n4691) );
  INVX1 U322 ( .A(\mem<14><5> ), .Y(n4687) );
  INVX1 U323 ( .A(\mem<14><6> ), .Y(n4686) );
  INVX1 U324 ( .A(\mem<14><7> ), .Y(n4685) );
  INVX1 U325 ( .A(\mem<13><0> ), .Y(n4684) );
  INVX1 U326 ( .A(\mem<13><1> ), .Y(n4683) );
  INVX1 U327 ( .A(\mem<13><2> ), .Y(n4682) );
  INVX1 U328 ( .A(\mem<13><3> ), .Y(n4681) );
  INVX1 U329 ( .A(\mem<13><4> ), .Y(n4680) );
  INVX1 U330 ( .A(\mem<13><5> ), .Y(n4679) );
  INVX1 U331 ( .A(\mem<13><6> ), .Y(n4678) );
  INVX1 U332 ( .A(\mem<13><7> ), .Y(n4677) );
  INVX1 U333 ( .A(\mem<12><0> ), .Y(n4676) );
  INVX1 U334 ( .A(\mem<12><1> ), .Y(n4675) );
  INVX1 U335 ( .A(\mem<12><5> ), .Y(n4671) );
  INVX1 U336 ( .A(\mem<12><6> ), .Y(n4670) );
  INVX1 U337 ( .A(\mem<12><7> ), .Y(n4669) );
  INVX1 U338 ( .A(\mem<11><0> ), .Y(n4668) );
  INVX1 U339 ( .A(\mem<11><1> ), .Y(n4667) );
  INVX1 U340 ( .A(\mem<11><2> ), .Y(n4666) );
  INVX1 U341 ( .A(\mem<11><3> ), .Y(n4665) );
  INVX1 U342 ( .A(\mem<11><4> ), .Y(n4664) );
  INVX1 U343 ( .A(\mem<11><5> ), .Y(n4663) );
  INVX1 U344 ( .A(\mem<11><6> ), .Y(n4662) );
  INVX1 U345 ( .A(\mem<11><7> ), .Y(n4661) );
  INVX1 U346 ( .A(\mem<10><0> ), .Y(n4660) );
  INVX1 U347 ( .A(\mem<10><1> ), .Y(n4659) );
  INVX1 U348 ( .A(\mem<10><5> ), .Y(n4655) );
  INVX1 U349 ( .A(\mem<10><6> ), .Y(n4654) );
  INVX1 U350 ( .A(\mem<10><7> ), .Y(n4653) );
  INVX1 U351 ( .A(\mem<9><0> ), .Y(n4652) );
  INVX1 U352 ( .A(\mem<9><1> ), .Y(n4651) );
  INVX1 U353 ( .A(\mem<9><2> ), .Y(n4650) );
  INVX1 U354 ( .A(\mem<9><3> ), .Y(n4649) );
  INVX1 U355 ( .A(\mem<9><4> ), .Y(n4648) );
  INVX1 U356 ( .A(\mem<9><5> ), .Y(n4647) );
  INVX1 U357 ( .A(\mem<9><6> ), .Y(n4646) );
  INVX1 U358 ( .A(\mem<9><7> ), .Y(n4645) );
  INVX1 U359 ( .A(\mem<8><0> ), .Y(n4644) );
  INVX1 U360 ( .A(\mem<8><1> ), .Y(n4643) );
  INVX1 U361 ( .A(\mem<8><5> ), .Y(n4639) );
  INVX1 U362 ( .A(\mem<8><6> ), .Y(n4638) );
  INVX1 U363 ( .A(\mem<8><7> ), .Y(n4637) );
  INVX1 U364 ( .A(\mem<7><0> ), .Y(n4636) );
  INVX1 U365 ( .A(\mem<7><1> ), .Y(n4635) );
  INVX1 U366 ( .A(\mem<7><2> ), .Y(n4634) );
  INVX1 U367 ( .A(\mem<7><3> ), .Y(n4633) );
  INVX1 U368 ( .A(\mem<7><4> ), .Y(n4632) );
  INVX1 U369 ( .A(\mem<7><5> ), .Y(n4631) );
  INVX1 U370 ( .A(\mem<7><6> ), .Y(n4630) );
  INVX1 U371 ( .A(\mem<7><7> ), .Y(n4629) );
  AND2X1 U372 ( .A(n456), .B(n1265), .Y(n1414) );
  INVX1 U373 ( .A(\mem<6><5> ), .Y(n4625) );
  INVX1 U374 ( .A(\mem<6><6> ), .Y(n4624) );
  INVX1 U375 ( .A(\mem<5><0> ), .Y(n4623) );
  INVX1 U376 ( .A(\mem<5><1> ), .Y(n4622) );
  INVX1 U377 ( .A(\mem<5><2> ), .Y(n4621) );
  INVX1 U378 ( .A(\mem<5><3> ), .Y(n4620) );
  INVX1 U379 ( .A(\mem<5><4> ), .Y(n4619) );
  INVX1 U380 ( .A(\mem<5><5> ), .Y(n4618) );
  INVX1 U381 ( .A(\mem<5><6> ), .Y(n4617) );
  INVX1 U382 ( .A(\mem<5><7> ), .Y(n4616) );
  AND2X1 U383 ( .A(n434), .B(n1269), .Y(n1418) );
  INVX1 U384 ( .A(\mem<4><5> ), .Y(n4611) );
  INVX1 U385 ( .A(\mem<4><6> ), .Y(n4610) );
  AND2X1 U386 ( .A(n530), .B(n1271), .Y(n1420) );
  INVX1 U387 ( .A(\mem<3><0> ), .Y(n4609) );
  INVX1 U388 ( .A(\mem<3><1> ), .Y(n4608) );
  INVX1 U389 ( .A(\mem<3><2> ), .Y(n4607) );
  INVX1 U390 ( .A(\mem<3><3> ), .Y(n4606) );
  INVX1 U391 ( .A(\mem<3><4> ), .Y(n4605) );
  INVX1 U392 ( .A(\mem<3><5> ), .Y(n4604) );
  INVX1 U393 ( .A(\mem<3><6> ), .Y(n4603) );
  INVX1 U394 ( .A(\mem<3><7> ), .Y(n4602) );
  INVX1 U395 ( .A(\mem<2><5> ), .Y(n4598) );
  INVX1 U396 ( .A(\mem<2><6> ), .Y(n4597) );
  AND2X1 U397 ( .A(n505), .B(n1275), .Y(n1424) );
  INVX1 U398 ( .A(\mem<1><5> ), .Y(n4593) );
  INVX1 U399 ( .A(\mem<1><6> ), .Y(n4592) );
  AND2X1 U400 ( .A(n467), .B(n4574), .Y(n1426) );
  AND2X1 U401 ( .A(n1294), .B(n467), .Y(n1283) );
  INVX1 U402 ( .A(n2541), .Y(n554) );
  AND2X1 U403 ( .A(n163), .B(n193), .Y(n261) );
  INVX1 U404 ( .A(n1295), .Y(n2629) );
  INVX1 U405 ( .A(n1295), .Y(n2630) );
  INVX1 U406 ( .A(n1295), .Y(n2631) );
  INVX1 U407 ( .A(n1295), .Y(n2628) );
  INVX1 U408 ( .A(n2548), .Y(n417) );
  INVX1 U409 ( .A(n2548), .Y(n519) );
  AND2X1 U410 ( .A(n620), .B(n669), .Y(n1049) );
  AND2X1 U411 ( .A(n624), .B(n673), .Y(n1051) );
  AND2X1 U412 ( .A(n629), .B(n677), .Y(n1053) );
  AND2X1 U413 ( .A(n633), .B(n681), .Y(n1055) );
  AND2X1 U414 ( .A(n637), .B(n685), .Y(n1057) );
  AND2X1 U415 ( .A(n641), .B(n689), .Y(n1059) );
  INVX1 U416 ( .A(wr), .Y(n2638) );
  AND2X1 U417 ( .A(n588), .B(n645), .Y(n1153) );
  AND2X1 U418 ( .A(n586), .B(n643), .Y(n1139) );
  OR2X1 U419 ( .A(n1036), .B(n1050), .Y(n1656) );
  AND2X1 U420 ( .A(n618), .B(n667), .Y(n1035) );
  AND2X1 U421 ( .A(n592), .B(n649), .Y(n1155) );
  AND2X1 U422 ( .A(n590), .B(n647), .Y(n1141) );
  OR2X1 U423 ( .A(n1038), .B(n1052), .Y(n1631) );
  AND2X1 U424 ( .A(n622), .B(n671), .Y(n1037) );
  AND2X1 U425 ( .A(n596), .B(n653), .Y(n1157) );
  AND2X1 U426 ( .A(n594), .B(n651), .Y(n1143) );
  OR2X1 U427 ( .A(n1040), .B(n1054), .Y(n1604) );
  AND2X1 U428 ( .A(n627), .B(n675), .Y(n1039) );
  AND2X1 U429 ( .A(n601), .B(n657), .Y(n1159) );
  AND2X1 U430 ( .A(n598), .B(n655), .Y(n1145) );
  OR2X1 U431 ( .A(n1042), .B(n1056), .Y(n1579) );
  AND2X1 U432 ( .A(n631), .B(n679), .Y(n1041) );
  AND2X1 U433 ( .A(n612), .B(n661), .Y(n1161) );
  AND2X1 U434 ( .A(n610), .B(n659), .Y(n1147) );
  OR2X1 U435 ( .A(n1044), .B(n1058), .Y(n1552) );
  AND2X1 U436 ( .A(n635), .B(n683), .Y(n1043) );
  AND2X1 U437 ( .A(n616), .B(n665), .Y(n1163) );
  AND2X1 U438 ( .A(n614), .B(n663), .Y(n1149) );
  OR2X1 U439 ( .A(n1046), .B(n1060), .Y(n1527) );
  AND2X1 U440 ( .A(n639), .B(n687), .Y(n1045) );
  INVX1 U441 ( .A(\mem<63><2> ), .Y(n5052) );
  INVX1 U442 ( .A(\mem<63><3> ), .Y(n5051) );
  INVX1 U443 ( .A(\mem<63><4> ), .Y(n5050) );
  INVX1 U444 ( .A(\mem<63><5> ), .Y(n5049) );
  INVX1 U445 ( .A(\mem<63><6> ), .Y(n5048) );
  INVX1 U446 ( .A(\data_in<0> ), .Y(n3017) );
  INVX1 U447 ( .A(n5047), .Y(n3015) );
  INVX1 U448 ( .A(\data_in<1> ), .Y(n3020) );
  INVX1 U449 ( .A(n5046), .Y(n3018) );
  INVX1 U450 ( .A(\data_in<2> ), .Y(n3023) );
  INVX1 U451 ( .A(n5045), .Y(n3021) );
  INVX1 U452 ( .A(\data_in<3> ), .Y(n3026) );
  INVX1 U453 ( .A(n5044), .Y(n3024) );
  INVX1 U454 ( .A(\data_in<4> ), .Y(n3029) );
  INVX1 U455 ( .A(n5043), .Y(n3027) );
  INVX1 U456 ( .A(\data_in<5> ), .Y(n3032) );
  INVX1 U457 ( .A(n2789), .Y(n3030) );
  INVX1 U458 ( .A(\data_in<6> ), .Y(n3035) );
  INVX1 U459 ( .A(n2831), .Y(n3033) );
  INVX1 U460 ( .A(\data_in<7> ), .Y(n3038) );
  INVX1 U461 ( .A(n5042), .Y(n3036) );
  INVX1 U462 ( .A(\data_in<0> ), .Y(n3042) );
  INVX1 U463 ( .A(n2686), .Y(n3040) );
  INVX1 U464 ( .A(\data_in<1> ), .Y(n3045) );
  INVX1 U465 ( .A(n2749), .Y(n3043) );
  INVX1 U466 ( .A(\data_in<2> ), .Y(n3048) );
  INVX1 U467 ( .A(n5041), .Y(n3046) );
  INVX1 U468 ( .A(\data_in<3> ), .Y(n3051) );
  INVX1 U469 ( .A(n5040), .Y(n3049) );
  INVX1 U470 ( .A(\data_in<4> ), .Y(n3054) );
  INVX1 U471 ( .A(n5039), .Y(n3052) );
  INVX1 U472 ( .A(\data_in<5> ), .Y(n3057) );
  INVX1 U473 ( .A(n5038), .Y(n3055) );
  INVX1 U474 ( .A(\data_in<6> ), .Y(n3060) );
  INVX1 U475 ( .A(n5037), .Y(n3058) );
  INVX1 U476 ( .A(\data_in<7> ), .Y(n3063) );
  INVX1 U477 ( .A(n2884), .Y(n3061) );
  INVX1 U478 ( .A(\data_in<0> ), .Y(n3068) );
  INVX1 U479 ( .A(n5036), .Y(n3066) );
  INVX1 U480 ( .A(\data_in<1> ), .Y(n3071) );
  INVX1 U481 ( .A(n5035), .Y(n3069) );
  INVX1 U482 ( .A(\data_in<2> ), .Y(n3074) );
  INVX1 U483 ( .A(n5034), .Y(n3072) );
  INVX1 U484 ( .A(\data_in<3> ), .Y(n3077) );
  INVX1 U485 ( .A(n5033), .Y(n3075) );
  INVX1 U486 ( .A(\data_in<4> ), .Y(n3080) );
  INVX1 U487 ( .A(n5032), .Y(n3078) );
  INVX1 U488 ( .A(\data_in<5> ), .Y(n3083) );
  INVX1 U489 ( .A(n2791), .Y(n3081) );
  INVX1 U490 ( .A(\data_in<6> ), .Y(n3086) );
  INVX1 U491 ( .A(n2833), .Y(n3084) );
  INVX1 U492 ( .A(\data_in<7> ), .Y(n3089) );
  INVX1 U493 ( .A(n5031), .Y(n3087) );
  INVX1 U494 ( .A(\data_in<0> ), .Y(n3094) );
  INVX1 U495 ( .A(n5030), .Y(n3092) );
  INVX1 U496 ( .A(\data_in<1> ), .Y(n3097) );
  INVX1 U497 ( .A(n2742), .Y(n3095) );
  INVX1 U498 ( .A(\data_in<2> ), .Y(n3100) );
  INVX1 U499 ( .A(n5029), .Y(n3098) );
  INVX1 U500 ( .A(\data_in<3> ), .Y(n3103) );
  INVX1 U501 ( .A(n5028), .Y(n3101) );
  INVX1 U502 ( .A(\data_in<4> ), .Y(n3106) );
  INVX1 U503 ( .A(n5027), .Y(n3104) );
  INVX1 U504 ( .A(\data_in<5> ), .Y(n3109) );
  INVX1 U505 ( .A(n5026), .Y(n3107) );
  INVX1 U506 ( .A(\data_in<6> ), .Y(n3112) );
  INVX1 U507 ( .A(n5025), .Y(n3110) );
  INVX1 U508 ( .A(\data_in<7> ), .Y(n3115) );
  INVX1 U509 ( .A(n2877), .Y(n3113) );
  INVX1 U510 ( .A(\data_in<0> ), .Y(n3119) );
  INVX1 U511 ( .A(n5024), .Y(n3117) );
  INVX1 U512 ( .A(\data_in<1> ), .Y(n3122) );
  INVX1 U513 ( .A(n5023), .Y(n3120) );
  INVX1 U514 ( .A(\data_in<2> ), .Y(n3125) );
  INVX1 U515 ( .A(n5022), .Y(n3123) );
  INVX1 U516 ( .A(\data_in<3> ), .Y(n3128) );
  INVX1 U517 ( .A(n5021), .Y(n3126) );
  INVX1 U518 ( .A(\data_in<4> ), .Y(n3131) );
  INVX1 U519 ( .A(n5020), .Y(n3129) );
  INVX1 U520 ( .A(\data_in<5> ), .Y(n3133) );
  INVX1 U521 ( .A(\data_in<6> ), .Y(n3136) );
  INVX1 U522 ( .A(n5019), .Y(n3134) );
  INVX1 U523 ( .A(\data_in<7> ), .Y(n3139) );
  INVX1 U524 ( .A(n5018), .Y(n3137) );
  INVX1 U525 ( .A(\data_in<0> ), .Y(n3144) );
  INVX1 U526 ( .A(n5017), .Y(n3142) );
  INVX1 U527 ( .A(\data_in<1> ), .Y(n3147) );
  INVX1 U528 ( .A(n5016), .Y(n3145) );
  INVX1 U529 ( .A(\data_in<2> ), .Y(n3150) );
  INVX1 U530 ( .A(n5015), .Y(n3148) );
  INVX1 U531 ( .A(\data_in<3> ), .Y(n3153) );
  INVX1 U532 ( .A(n5014), .Y(n3151) );
  INVX1 U533 ( .A(\data_in<4> ), .Y(n3156) );
  INVX1 U534 ( .A(n5013), .Y(n3154) );
  INVX1 U535 ( .A(\data_in<5> ), .Y(n3159) );
  INVX1 U536 ( .A(n2785), .Y(n3157) );
  INVX1 U537 ( .A(\data_in<6> ), .Y(n3162) );
  INVX1 U538 ( .A(n2827), .Y(n3160) );
  INVX1 U539 ( .A(\data_in<7> ), .Y(n3165) );
  INVX1 U540 ( .A(n5012), .Y(n3163) );
  INVX1 U541 ( .A(\data_in<0> ), .Y(n3170) );
  INVX1 U542 ( .A(n5011), .Y(n3168) );
  INVX1 U543 ( .A(\data_in<1> ), .Y(n3173) );
  INVX1 U544 ( .A(n5010), .Y(n3171) );
  INVX1 U545 ( .A(\data_in<2> ), .Y(n3176) );
  INVX1 U546 ( .A(n5009), .Y(n3174) );
  INVX1 U547 ( .A(\data_in<3> ), .Y(n3179) );
  INVX1 U548 ( .A(n5008), .Y(n3177) );
  INVX1 U549 ( .A(\data_in<4> ), .Y(n3182) );
  INVX1 U550 ( .A(n5007), .Y(n3180) );
  INVX1 U551 ( .A(\data_in<5> ), .Y(n3185) );
  INVX1 U552 ( .A(n5006), .Y(n3183) );
  INVX1 U553 ( .A(\data_in<6> ), .Y(n3188) );
  INVX1 U554 ( .A(n5005), .Y(n3186) );
  INVX1 U555 ( .A(\data_in<7> ), .Y(n3191) );
  INVX1 U556 ( .A(n5004), .Y(n3189) );
  INVX1 U557 ( .A(\data_in<0> ), .Y(n3195) );
  INVX1 U558 ( .A(n5003), .Y(n3193) );
  INVX1 U559 ( .A(\data_in<1> ), .Y(n3198) );
  INVX1 U560 ( .A(n5002), .Y(n3196) );
  INVX1 U561 ( .A(\data_in<2> ), .Y(n3201) );
  INVX1 U562 ( .A(n5001), .Y(n3199) );
  INVX1 U563 ( .A(\data_in<3> ), .Y(n3204) );
  INVX1 U564 ( .A(n5000), .Y(n3202) );
  INVX1 U565 ( .A(\data_in<4> ), .Y(n3207) );
  INVX1 U566 ( .A(n4999), .Y(n3205) );
  INVX1 U567 ( .A(\data_in<5> ), .Y(n3210) );
  INVX1 U568 ( .A(n4998), .Y(n3208) );
  INVX1 U569 ( .A(\data_in<6> ), .Y(n3213) );
  INVX1 U570 ( .A(n4997), .Y(n3211) );
  INVX1 U571 ( .A(\data_in<7> ), .Y(n3217) );
  INVX1 U572 ( .A(n4996), .Y(n3215) );
  INVX1 U573 ( .A(\data_in<0> ), .Y(n3220) );
  INVX1 U574 ( .A(n4995), .Y(n3218) );
  INVX1 U575 ( .A(\data_in<1> ), .Y(n3223) );
  INVX1 U576 ( .A(n4994), .Y(n3221) );
  INVX1 U577 ( .A(\data_in<2> ), .Y(n3226) );
  INVX1 U578 ( .A(n4993), .Y(n3224) );
  INVX1 U579 ( .A(\data_in<3> ), .Y(n3229) );
  INVX1 U580 ( .A(n4992), .Y(n3227) );
  INVX1 U581 ( .A(\data_in<4> ), .Y(n3232) );
  INVX1 U582 ( .A(n4991), .Y(n3230) );
  INVX1 U583 ( .A(\data_in<5> ), .Y(n3235) );
  INVX1 U584 ( .A(n4990), .Y(n3233) );
  INVX1 U585 ( .A(\data_in<6> ), .Y(n3238) );
  INVX1 U586 ( .A(n4989), .Y(n3236) );
  INVX1 U587 ( .A(\data_in<7> ), .Y(n3241) );
  INVX1 U588 ( .A(n4988), .Y(n3239) );
  INVX1 U589 ( .A(\data_in<0> ), .Y(n3245) );
  INVX1 U590 ( .A(n4987), .Y(n3243) );
  INVX1 U591 ( .A(\data_in<1> ), .Y(n3248) );
  INVX1 U592 ( .A(n4986), .Y(n3246) );
  INVX1 U593 ( .A(\data_in<2> ), .Y(n3251) );
  INVX1 U594 ( .A(n4985), .Y(n3249) );
  INVX1 U595 ( .A(\data_in<3> ), .Y(n3254) );
  INVX1 U596 ( .A(n4984), .Y(n3252) );
  INVX1 U597 ( .A(\data_in<4> ), .Y(n3257) );
  INVX1 U598 ( .A(n4983), .Y(n3255) );
  INVX1 U599 ( .A(\data_in<5> ), .Y(n3260) );
  INVX1 U600 ( .A(n4982), .Y(n3258) );
  INVX1 U601 ( .A(\data_in<6> ), .Y(n3263) );
  INVX1 U602 ( .A(n4981), .Y(n3261) );
  INVX1 U603 ( .A(\data_in<7> ), .Y(n3266) );
  INVX1 U604 ( .A(n4980), .Y(n3264) );
  INVX1 U605 ( .A(\data_in<0> ), .Y(n3271) );
  INVX1 U606 ( .A(n4979), .Y(n3269) );
  INVX1 U607 ( .A(\data_in<1> ), .Y(n3274) );
  INVX1 U608 ( .A(n4978), .Y(n3272) );
  INVX1 U609 ( .A(\data_in<2> ), .Y(n3277) );
  INVX1 U610 ( .A(n4977), .Y(n3275) );
  INVX1 U611 ( .A(\data_in<3> ), .Y(n3280) );
  INVX1 U612 ( .A(n4976), .Y(n3278) );
  INVX1 U613 ( .A(\data_in<4> ), .Y(n3283) );
  INVX1 U614 ( .A(n4975), .Y(n3281) );
  INVX1 U615 ( .A(\data_in<5> ), .Y(n3286) );
  INVX1 U616 ( .A(n4974), .Y(n3284) );
  INVX1 U617 ( .A(\data_in<6> ), .Y(n3289) );
  INVX1 U618 ( .A(n4973), .Y(n3287) );
  INVX1 U619 ( .A(\data_in<7> ), .Y(n3293) );
  INVX1 U620 ( .A(n4972), .Y(n3291) );
  INVX1 U621 ( .A(\data_in<0> ), .Y(n3297) );
  INVX1 U622 ( .A(n4971), .Y(n3295) );
  INVX1 U623 ( .A(\data_in<1> ), .Y(n3300) );
  INVX1 U624 ( .A(n4970), .Y(n3298) );
  INVX1 U625 ( .A(\data_in<2> ), .Y(n3303) );
  INVX1 U626 ( .A(n4969), .Y(n3301) );
  INVX1 U627 ( .A(\data_in<3> ), .Y(n3306) );
  INVX1 U628 ( .A(n4968), .Y(n3304) );
  INVX1 U629 ( .A(\data_in<4> ), .Y(n3309) );
  INVX1 U630 ( .A(n4967), .Y(n3307) );
  INVX1 U631 ( .A(\data_in<5> ), .Y(n3312) );
  INVX1 U632 ( .A(n4966), .Y(n3310) );
  INVX1 U633 ( .A(\data_in<6> ), .Y(n3315) );
  INVX1 U634 ( .A(n4965), .Y(n3313) );
  INVX1 U635 ( .A(\data_in<7> ), .Y(n3319) );
  INVX1 U636 ( .A(n4964), .Y(n3317) );
  INVX1 U637 ( .A(\data_in<0> ), .Y(n3325) );
  INVX1 U638 ( .A(n4963), .Y(n3323) );
  INVX1 U639 ( .A(\data_in<1> ), .Y(n3328) );
  INVX1 U640 ( .A(n4962), .Y(n3326) );
  INVX1 U641 ( .A(\data_in<2> ), .Y(n3331) );
  INVX1 U642 ( .A(n4961), .Y(n3329) );
  INVX1 U643 ( .A(\data_in<3> ), .Y(n3334) );
  INVX1 U644 ( .A(n4960), .Y(n3332) );
  INVX1 U645 ( .A(\data_in<4> ), .Y(n3337) );
  INVX1 U646 ( .A(n4959), .Y(n3335) );
  INVX1 U647 ( .A(\data_in<5> ), .Y(n3340) );
  INVX1 U648 ( .A(n4958), .Y(n3338) );
  INVX1 U649 ( .A(\data_in<6> ), .Y(n3343) );
  INVX1 U650 ( .A(n4957), .Y(n3341) );
  INVX1 U651 ( .A(\data_in<7> ), .Y(n3347) );
  INVX1 U652 ( .A(n4956), .Y(n3345) );
  INVX1 U653 ( .A(\data_in<0> ), .Y(n3351) );
  INVX1 U654 ( .A(n4955), .Y(n3349) );
  INVX1 U655 ( .A(\data_in<1> ), .Y(n3354) );
  INVX1 U656 ( .A(n4954), .Y(n3352) );
  INVX1 U657 ( .A(\data_in<2> ), .Y(n3357) );
  INVX1 U658 ( .A(n4953), .Y(n3355) );
  INVX1 U659 ( .A(\data_in<3> ), .Y(n3360) );
  INVX1 U660 ( .A(n4952), .Y(n3358) );
  INVX1 U661 ( .A(\data_in<4> ), .Y(n3363) );
  INVX1 U662 ( .A(n4951), .Y(n3361) );
  INVX1 U663 ( .A(\data_in<5> ), .Y(n3366) );
  INVX1 U664 ( .A(n4950), .Y(n3364) );
  INVX1 U665 ( .A(\data_in<6> ), .Y(n3369) );
  INVX1 U666 ( .A(n4949), .Y(n3367) );
  INVX1 U667 ( .A(\data_in<7> ), .Y(n3373) );
  INVX1 U668 ( .A(n4948), .Y(n3371) );
  INVX1 U669 ( .A(\data_in<0> ), .Y(n3376) );
  INVX1 U670 ( .A(n4947), .Y(n3374) );
  INVX1 U671 ( .A(\data_in<1> ), .Y(n3379) );
  INVX1 U672 ( .A(n4946), .Y(n3377) );
  INVX1 U673 ( .A(\data_in<2> ), .Y(n3382) );
  INVX1 U674 ( .A(n4945), .Y(n3380) );
  INVX1 U675 ( .A(\data_in<3> ), .Y(n3385) );
  INVX1 U676 ( .A(n4944), .Y(n3383) );
  INVX1 U677 ( .A(\data_in<4> ), .Y(n3388) );
  INVX1 U678 ( .A(n4943), .Y(n3386) );
  INVX1 U679 ( .A(\data_in<5> ), .Y(n3391) );
  INVX1 U680 ( .A(n4942), .Y(n3389) );
  INVX1 U681 ( .A(\data_in<6> ), .Y(n3394) );
  INVX1 U682 ( .A(n4941), .Y(n3392) );
  INVX1 U683 ( .A(\data_in<7> ), .Y(n3397) );
  INVX1 U684 ( .A(n4940), .Y(n3395) );
  INVX1 U685 ( .A(\data_in<0> ), .Y(n3401) );
  INVX1 U686 ( .A(n4939), .Y(n3399) );
  INVX1 U687 ( .A(\data_in<1> ), .Y(n3404) );
  INVX1 U688 ( .A(n4938), .Y(n3402) );
  INVX1 U689 ( .A(\data_in<2> ), .Y(n3407) );
  INVX1 U690 ( .A(n4937), .Y(n3405) );
  INVX1 U691 ( .A(\data_in<3> ), .Y(n3410) );
  INVX1 U692 ( .A(n4936), .Y(n3408) );
  INVX1 U693 ( .A(\data_in<4> ), .Y(n3413) );
  INVX1 U694 ( .A(n4935), .Y(n3411) );
  INVX1 U695 ( .A(\data_in<5> ), .Y(n3416) );
  INVX1 U696 ( .A(n4934), .Y(n3414) );
  INVX1 U697 ( .A(\data_in<6> ), .Y(n3419) );
  INVX1 U698 ( .A(n4933), .Y(n3417) );
  INVX1 U699 ( .A(\data_in<7> ), .Y(n3422) );
  INVX1 U700 ( .A(n4932), .Y(n3420) );
  INVX1 U701 ( .A(\data_in<0> ), .Y(n3426) );
  INVX1 U702 ( .A(n4931), .Y(n3424) );
  INVX1 U703 ( .A(\data_in<1> ), .Y(n3429) );
  INVX1 U704 ( .A(n4930), .Y(n3427) );
  INVX1 U705 ( .A(\data_in<2> ), .Y(n3432) );
  INVX1 U706 ( .A(n4929), .Y(n3430) );
  INVX1 U707 ( .A(\data_in<3> ), .Y(n3435) );
  INVX1 U708 ( .A(n4928), .Y(n3433) );
  INVX1 U709 ( .A(\data_in<4> ), .Y(n3438) );
  INVX1 U710 ( .A(n4927), .Y(n3436) );
  INVX1 U711 ( .A(\data_in<5> ), .Y(n3441) );
  INVX1 U712 ( .A(n4926), .Y(n3439) );
  INVX1 U713 ( .A(\data_in<6> ), .Y(n3444) );
  INVX1 U714 ( .A(n4925), .Y(n3442) );
  INVX1 U715 ( .A(\data_in<7> ), .Y(n3447) );
  INVX1 U716 ( .A(n4924), .Y(n3445) );
  INVX1 U717 ( .A(\data_in<0> ), .Y(n3451) );
  INVX1 U718 ( .A(n4923), .Y(n3449) );
  INVX1 U719 ( .A(\data_in<1> ), .Y(n3454) );
  INVX1 U720 ( .A(n4922), .Y(n3452) );
  INVX1 U721 ( .A(\data_in<2> ), .Y(n3457) );
  INVX1 U722 ( .A(n4921), .Y(n3455) );
  INVX1 U723 ( .A(\data_in<3> ), .Y(n3460) );
  INVX1 U724 ( .A(n4920), .Y(n3458) );
  INVX1 U725 ( .A(\data_in<4> ), .Y(n3463) );
  INVX1 U726 ( .A(n4919), .Y(n3461) );
  INVX1 U727 ( .A(\data_in<5> ), .Y(n3466) );
  INVX1 U728 ( .A(n4918), .Y(n3464) );
  INVX1 U729 ( .A(\data_in<6> ), .Y(n3469) );
  INVX1 U730 ( .A(n4917), .Y(n3467) );
  INVX1 U731 ( .A(\data_in<7> ), .Y(n3472) );
  INVX1 U732 ( .A(n4916), .Y(n3470) );
  INVX1 U733 ( .A(\data_in<0> ), .Y(n3476) );
  INVX1 U734 ( .A(n4915), .Y(n3474) );
  INVX1 U735 ( .A(\data_in<1> ), .Y(n3479) );
  INVX1 U736 ( .A(n4914), .Y(n3477) );
  INVX1 U737 ( .A(\data_in<2> ), .Y(n3482) );
  INVX1 U738 ( .A(n4913), .Y(n3480) );
  INVX1 U739 ( .A(\data_in<3> ), .Y(n3485) );
  INVX1 U740 ( .A(n4912), .Y(n3483) );
  INVX1 U741 ( .A(\data_in<4> ), .Y(n3488) );
  INVX1 U742 ( .A(n4911), .Y(n3486) );
  INVX1 U743 ( .A(\data_in<5> ), .Y(n3491) );
  INVX1 U744 ( .A(n4910), .Y(n3489) );
  INVX1 U745 ( .A(\data_in<6> ), .Y(n3494) );
  INVX1 U746 ( .A(n4909), .Y(n3492) );
  INVX1 U747 ( .A(\data_in<7> ), .Y(n3497) );
  INVX1 U748 ( .A(n4908), .Y(n3495) );
  INVX1 U749 ( .A(\data_in<0> ), .Y(n3500) );
  INVX1 U750 ( .A(n4907), .Y(n3498) );
  INVX1 U751 ( .A(\data_in<1> ), .Y(n3503) );
  INVX1 U752 ( .A(n4906), .Y(n3501) );
  INVX1 U753 ( .A(\data_in<2> ), .Y(n3506) );
  INVX1 U754 ( .A(n4905), .Y(n3504) );
  INVX1 U755 ( .A(\data_in<3> ), .Y(n3509) );
  INVX1 U756 ( .A(n4904), .Y(n3507) );
  INVX1 U757 ( .A(\data_in<4> ), .Y(n3512) );
  INVX1 U758 ( .A(n4903), .Y(n3510) );
  INVX1 U759 ( .A(\data_in<5> ), .Y(n3515) );
  INVX1 U760 ( .A(n4902), .Y(n3513) );
  INVX1 U761 ( .A(\data_in<6> ), .Y(n3518) );
  INVX1 U762 ( .A(n4901), .Y(n3516) );
  INVX1 U763 ( .A(\data_in<7> ), .Y(n3521) );
  INVX1 U764 ( .A(n4900), .Y(n3519) );
  INVX1 U765 ( .A(\data_in<0> ), .Y(n3525) );
  INVX1 U766 ( .A(n4899), .Y(n3523) );
  INVX1 U767 ( .A(\data_in<1> ), .Y(n3528) );
  INVX1 U768 ( .A(n4898), .Y(n3526) );
  INVX1 U769 ( .A(\data_in<2> ), .Y(n3531) );
  INVX1 U770 ( .A(n4897), .Y(n3529) );
  INVX1 U771 ( .A(\data_in<3> ), .Y(n3534) );
  INVX1 U772 ( .A(n4896), .Y(n3532) );
  INVX1 U773 ( .A(\data_in<4> ), .Y(n3537) );
  INVX1 U774 ( .A(n4895), .Y(n3535) );
  INVX1 U775 ( .A(\data_in<5> ), .Y(n3540) );
  INVX1 U776 ( .A(n4894), .Y(n3538) );
  INVX1 U777 ( .A(\data_in<6> ), .Y(n3543) );
  INVX1 U778 ( .A(n4893), .Y(n3541) );
  INVX1 U779 ( .A(\data_in<7> ), .Y(n3546) );
  INVX1 U780 ( .A(n4892), .Y(n3544) );
  INVX1 U781 ( .A(\data_in<0> ), .Y(n3550) );
  INVX1 U782 ( .A(n4891), .Y(n3548) );
  INVX1 U783 ( .A(\data_in<1> ), .Y(n3553) );
  INVX1 U784 ( .A(n4890), .Y(n3551) );
  INVX1 U785 ( .A(\data_in<2> ), .Y(n3556) );
  INVX1 U786 ( .A(n4889), .Y(n3554) );
  INVX1 U787 ( .A(\data_in<3> ), .Y(n3559) );
  INVX1 U788 ( .A(n4888), .Y(n3557) );
  INVX1 U789 ( .A(\data_in<4> ), .Y(n3562) );
  INVX1 U790 ( .A(n4887), .Y(n3560) );
  INVX1 U791 ( .A(\data_in<5> ), .Y(n3565) );
  INVX1 U792 ( .A(n4886), .Y(n3563) );
  INVX1 U793 ( .A(\data_in<6> ), .Y(n3568) );
  INVX1 U794 ( .A(n4885), .Y(n3566) );
  INVX1 U795 ( .A(\data_in<7> ), .Y(n3571) );
  INVX1 U796 ( .A(n4884), .Y(n3569) );
  INVX1 U797 ( .A(\data_in<0> ), .Y(n3575) );
  INVX1 U798 ( .A(n4883), .Y(n3573) );
  INVX1 U799 ( .A(\data_in<1> ), .Y(n3578) );
  INVX1 U800 ( .A(n4882), .Y(n3576) );
  INVX1 U801 ( .A(\data_in<2> ), .Y(n3581) );
  INVX1 U802 ( .A(n4881), .Y(n3579) );
  INVX1 U803 ( .A(\data_in<3> ), .Y(n3584) );
  INVX1 U804 ( .A(n4880), .Y(n3582) );
  INVX1 U805 ( .A(\data_in<4> ), .Y(n3587) );
  INVX1 U806 ( .A(n4879), .Y(n3585) );
  INVX1 U807 ( .A(\data_in<5> ), .Y(n3590) );
  INVX1 U808 ( .A(n4878), .Y(n3588) );
  INVX1 U809 ( .A(\data_in<6> ), .Y(n3593) );
  INVX1 U810 ( .A(n4877), .Y(n3591) );
  INVX1 U811 ( .A(\data_in<7> ), .Y(n3596) );
  INVX1 U812 ( .A(n4876), .Y(n3594) );
  INVX1 U813 ( .A(\data_in<0> ), .Y(n3600) );
  INVX1 U814 ( .A(n4875), .Y(n3598) );
  INVX1 U815 ( .A(\data_in<1> ), .Y(n3603) );
  INVX1 U816 ( .A(n4874), .Y(n3601) );
  INVX1 U818 ( .A(\data_in<2> ), .Y(n3606) );
  INVX1 U820 ( .A(n4873), .Y(n3604) );
  INVX1 U822 ( .A(\data_in<3> ), .Y(n3609) );
  INVX1 U824 ( .A(n557), .Y(n3607) );
  INVX1 U826 ( .A(\data_in<4> ), .Y(n3612) );
  INVX1 U828 ( .A(n4872), .Y(n3610) );
  INVX1 U830 ( .A(\data_in<5> ), .Y(n3615) );
  INVX1 U832 ( .A(n4871), .Y(n3613) );
  INVX1 U833 ( .A(\data_in<6> ), .Y(n3618) );
  INVX1 U834 ( .A(n4870), .Y(n3616) );
  INVX1 U835 ( .A(\data_in<7> ), .Y(n3621) );
  INVX1 U836 ( .A(n4869), .Y(n3619) );
  INVX1 U837 ( .A(\data_in<0> ), .Y(n3624) );
  INVX1 U838 ( .A(n4868), .Y(n3622) );
  INVX1 U839 ( .A(\data_in<1> ), .Y(n3627) );
  INVX1 U840 ( .A(n4867), .Y(n3625) );
  INVX1 U841 ( .A(\data_in<2> ), .Y(n3630) );
  INVX1 U842 ( .A(n4866), .Y(n3628) );
  INVX1 U843 ( .A(\data_in<3> ), .Y(n3633) );
  INVX1 U844 ( .A(n556), .Y(n3631) );
  INVX1 U845 ( .A(\data_in<4> ), .Y(n3636) );
  INVX1 U846 ( .A(n4865), .Y(n3634) );
  INVX1 U847 ( .A(\data_in<5> ), .Y(n3639) );
  INVX1 U848 ( .A(n4864), .Y(n3637) );
  INVX1 U849 ( .A(\data_in<6> ), .Y(n3642) );
  INVX1 U850 ( .A(n4863), .Y(n3640) );
  INVX1 U851 ( .A(\data_in<7> ), .Y(n3645) );
  INVX1 U852 ( .A(n4862), .Y(n3643) );
  INVX1 U853 ( .A(\data_in<0> ), .Y(n3649) );
  INVX1 U854 ( .A(n4861), .Y(n3647) );
  INVX1 U855 ( .A(\data_in<1> ), .Y(n3652) );
  INVX1 U856 ( .A(n4860), .Y(n3650) );
  INVX1 U857 ( .A(\data_in<2> ), .Y(n3655) );
  INVX1 U858 ( .A(n4859), .Y(n3653) );
  INVX1 U859 ( .A(\data_in<3> ), .Y(n3658) );
  INVX1 U860 ( .A(n4858), .Y(n3656) );
  INVX1 U861 ( .A(\data_in<4> ), .Y(n3661) );
  INVX1 U862 ( .A(n4857), .Y(n3659) );
  INVX1 U863 ( .A(\data_in<5> ), .Y(n3664) );
  INVX1 U864 ( .A(n4856), .Y(n3662) );
  INVX1 U865 ( .A(\data_in<6> ), .Y(n3667) );
  INVX1 U866 ( .A(n4855), .Y(n3665) );
  INVX1 U867 ( .A(\data_in<7> ), .Y(n3670) );
  INVX1 U868 ( .A(n4854), .Y(n3668) );
  INVX1 U869 ( .A(\data_in<0> ), .Y(n3674) );
  INVX1 U870 ( .A(n4853), .Y(n3672) );
  INVX1 U871 ( .A(\data_in<1> ), .Y(n3677) );
  INVX1 U872 ( .A(n4852), .Y(n3675) );
  INVX1 U873 ( .A(\data_in<2> ), .Y(n3680) );
  INVX1 U874 ( .A(n4851), .Y(n3678) );
  INVX1 U875 ( .A(\data_in<3> ), .Y(n3683) );
  INVX1 U876 ( .A(n4850), .Y(n3681) );
  INVX1 U877 ( .A(\data_in<4> ), .Y(n3686) );
  INVX1 U878 ( .A(n4849), .Y(n3684) );
  INVX1 U879 ( .A(\data_in<5> ), .Y(n3689) );
  INVX1 U880 ( .A(n4848), .Y(n3687) );
  INVX1 U881 ( .A(\data_in<6> ), .Y(n3692) );
  INVX1 U882 ( .A(n4847), .Y(n3690) );
  INVX1 U883 ( .A(\data_in<7> ), .Y(n3695) );
  INVX1 U884 ( .A(n4846), .Y(n3693) );
  INVX1 U885 ( .A(\data_in<0> ), .Y(n3699) );
  INVX1 U886 ( .A(n4845), .Y(n3697) );
  INVX1 U887 ( .A(\data_in<1> ), .Y(n3702) );
  INVX1 U888 ( .A(n4844), .Y(n3700) );
  INVX1 U889 ( .A(\data_in<2> ), .Y(n3705) );
  INVX1 U890 ( .A(n4843), .Y(n3703) );
  INVX1 U891 ( .A(\data_in<3> ), .Y(n3708) );
  INVX1 U892 ( .A(n4842), .Y(n3706) );
  INVX1 U893 ( .A(\data_in<4> ), .Y(n3711) );
  INVX1 U894 ( .A(n4841), .Y(n3709) );
  INVX1 U895 ( .A(\data_in<5> ), .Y(n3714) );
  INVX1 U896 ( .A(n4840), .Y(n3712) );
  INVX1 U897 ( .A(\data_in<6> ), .Y(n3717) );
  INVX1 U898 ( .A(n4839), .Y(n3715) );
  INVX1 U899 ( .A(\data_in<7> ), .Y(n3720) );
  INVX1 U900 ( .A(n4838), .Y(n3718) );
  INVX1 U901 ( .A(\data_in<0> ), .Y(n3724) );
  INVX1 U902 ( .A(n4837), .Y(n3722) );
  INVX1 U903 ( .A(\data_in<1> ), .Y(n3727) );
  INVX1 U904 ( .A(n4836), .Y(n3725) );
  INVX1 U905 ( .A(\data_in<2> ), .Y(n3730) );
  INVX1 U906 ( .A(n4835), .Y(n3728) );
  INVX1 U907 ( .A(\data_in<3> ), .Y(n3733) );
  INVX1 U908 ( .A(n4834), .Y(n3731) );
  INVX1 U909 ( .A(\data_in<4> ), .Y(n3736) );
  INVX1 U910 ( .A(n4833), .Y(n3734) );
  INVX1 U911 ( .A(\data_in<5> ), .Y(n3739) );
  INVX1 U912 ( .A(n4832), .Y(n3737) );
  INVX1 U913 ( .A(\data_in<6> ), .Y(n3742) );
  INVX1 U914 ( .A(n4831), .Y(n3740) );
  INVX1 U915 ( .A(\data_in<7> ), .Y(n3745) );
  INVX1 U916 ( .A(n4830), .Y(n3743) );
  INVX1 U917 ( .A(\data_in<0> ), .Y(n3750) );
  INVX1 U918 ( .A(n4829), .Y(n3748) );
  INVX1 U919 ( .A(\data_in<1> ), .Y(n3753) );
  INVX1 U920 ( .A(n4828), .Y(n3751) );
  INVX1 U921 ( .A(\data_in<2> ), .Y(n3756) );
  INVX1 U922 ( .A(n4827), .Y(n3754) );
  INVX1 U923 ( .A(\data_in<3> ), .Y(n3759) );
  INVX1 U924 ( .A(n4826), .Y(n3757) );
  INVX1 U925 ( .A(\data_in<4> ), .Y(n3762) );
  INVX1 U926 ( .A(n4825), .Y(n3760) );
  INVX1 U927 ( .A(\data_in<5> ), .Y(n3765) );
  INVX1 U928 ( .A(n4824), .Y(n3763) );
  INVX1 U929 ( .A(\data_in<6> ), .Y(n3768) );
  INVX1 U930 ( .A(n4823), .Y(n3766) );
  INVX1 U931 ( .A(\data_in<7> ), .Y(n3771) );
  INVX1 U932 ( .A(n4822), .Y(n3769) );
  INVX1 U933 ( .A(\data_in<0> ), .Y(n3775) );
  INVX1 U934 ( .A(n2679), .Y(n3773) );
  INVX1 U935 ( .A(\data_in<1> ), .Y(n3778) );
  INVX1 U936 ( .A(n2743), .Y(n3776) );
  INVX1 U937 ( .A(\data_in<2> ), .Y(n3781) );
  INVX1 U938 ( .A(n4821), .Y(n3779) );
  INVX1 U939 ( .A(\data_in<3> ), .Y(n3784) );
  INVX1 U940 ( .A(n4820), .Y(n3782) );
  INVX1 U941 ( .A(\data_in<4> ), .Y(n3787) );
  INVX1 U942 ( .A(n4819), .Y(n3785) );
  INVX1 U943 ( .A(\data_in<5> ), .Y(n3790) );
  INVX1 U944 ( .A(n4818), .Y(n3788) );
  INVX1 U945 ( .A(\data_in<6> ), .Y(n3793) );
  INVX1 U946 ( .A(n4817), .Y(n3791) );
  INVX1 U947 ( .A(\data_in<7> ), .Y(n3796) );
  INVX1 U948 ( .A(n2878), .Y(n3794) );
  INVX1 U949 ( .A(\data_in<0> ), .Y(n3801) );
  INVX1 U950 ( .A(n4816), .Y(n3799) );
  INVX1 U951 ( .A(\data_in<1> ), .Y(n3804) );
  INVX1 U952 ( .A(n4815), .Y(n3802) );
  INVX1 U953 ( .A(\data_in<2> ), .Y(n3807) );
  INVX1 U954 ( .A(n4814), .Y(n3805) );
  INVX1 U955 ( .A(\data_in<3> ), .Y(n3810) );
  INVX1 U956 ( .A(n4813), .Y(n3808) );
  INVX1 U957 ( .A(\data_in<4> ), .Y(n3813) );
  INVX1 U958 ( .A(n4812), .Y(n3811) );
  INVX1 U959 ( .A(\data_in<5> ), .Y(n3816) );
  INVX1 U960 ( .A(n4811), .Y(n3814) );
  INVX1 U961 ( .A(\data_in<6> ), .Y(n3819) );
  INVX1 U962 ( .A(n4810), .Y(n3817) );
  INVX1 U963 ( .A(\data_in<7> ), .Y(n3822) );
  INVX1 U964 ( .A(n4809), .Y(n3820) );
  INVX1 U965 ( .A(\data_in<0> ), .Y(n3826) );
  INVX1 U966 ( .A(n4808), .Y(n3824) );
  INVX1 U967 ( .A(\data_in<1> ), .Y(n3829) );
  INVX1 U968 ( .A(n4807), .Y(n3827) );
  INVX1 U969 ( .A(\data_in<2> ), .Y(n3832) );
  INVX1 U970 ( .A(n4806), .Y(n3830) );
  INVX1 U971 ( .A(\data_in<3> ), .Y(n3835) );
  INVX1 U972 ( .A(n4805), .Y(n3833) );
  INVX1 U973 ( .A(\data_in<4> ), .Y(n3838) );
  INVX1 U974 ( .A(n4804), .Y(n3836) );
  INVX1 U975 ( .A(\data_in<5> ), .Y(n3841) );
  INVX1 U976 ( .A(n4803), .Y(n3839) );
  INVX1 U977 ( .A(\data_in<6> ), .Y(n3844) );
  INVX1 U978 ( .A(n4802), .Y(n3842) );
  INVX1 U979 ( .A(\data_in<7> ), .Y(n3847) );
  INVX1 U980 ( .A(n4801), .Y(n3845) );
  INVX1 U981 ( .A(\data_in<0> ), .Y(n3852) );
  INVX1 U982 ( .A(n4800), .Y(n3850) );
  INVX1 U983 ( .A(\data_in<1> ), .Y(n3855) );
  INVX1 U984 ( .A(n4799), .Y(n3853) );
  INVX1 U985 ( .A(\data_in<2> ), .Y(n3858) );
  INVX1 U986 ( .A(n4798), .Y(n3856) );
  INVX1 U987 ( .A(\data_in<3> ), .Y(n3861) );
  INVX1 U988 ( .A(n4797), .Y(n3859) );
  INVX1 U989 ( .A(\data_in<4> ), .Y(n3864) );
  INVX1 U990 ( .A(n4796), .Y(n3862) );
  INVX1 U991 ( .A(\data_in<5> ), .Y(n3867) );
  INVX1 U992 ( .A(n2795), .Y(n3865) );
  INVX1 U993 ( .A(\data_in<6> ), .Y(n3870) );
  INVX1 U994 ( .A(n2837), .Y(n3868) );
  INVX1 U995 ( .A(\data_in<7> ), .Y(n3873) );
  INVX1 U996 ( .A(n4795), .Y(n3871) );
  INVX1 U997 ( .A(\data_in<0> ), .Y(n3878) );
  INVX1 U998 ( .A(n2702), .Y(n3876) );
  INVX1 U999 ( .A(\data_in<1> ), .Y(n3881) );
  INVX1 U1000 ( .A(\data_in<2> ), .Y(n3884) );
  INVX1 U1001 ( .A(n4793), .Y(n3882) );
  INVX1 U1002 ( .A(\data_in<3> ), .Y(n3887) );
  INVX1 U1003 ( .A(n4792), .Y(n3885) );
  INVX1 U1004 ( .A(\data_in<4> ), .Y(n3890) );
  INVX1 U1005 ( .A(n4791), .Y(n3888) );
  INVX1 U1006 ( .A(\data_in<5> ), .Y(n3893) );
  INVX1 U1007 ( .A(n4790), .Y(n3891) );
  INVX1 U1008 ( .A(\data_in<6> ), .Y(n3896) );
  INVX1 U1009 ( .A(n4789), .Y(n3894) );
  INVX1 U1010 ( .A(\data_in<7> ), .Y(n3899) );
  INVX1 U1011 ( .A(n2896), .Y(n3897) );
  INVX1 U1012 ( .A(\data_in<0> ), .Y(n3904) );
  INVX1 U1013 ( .A(n4788), .Y(n3902) );
  INVX1 U1014 ( .A(\data_in<1> ), .Y(n3907) );
  INVX1 U1015 ( .A(n4787), .Y(n3905) );
  INVX1 U1016 ( .A(\data_in<2> ), .Y(n3910) );
  INVX1 U1017 ( .A(n4786), .Y(n3908) );
  INVX1 U1018 ( .A(\data_in<3> ), .Y(n3913) );
  INVX1 U1019 ( .A(n4785), .Y(n3911) );
  INVX1 U1020 ( .A(\data_in<4> ), .Y(n3916) );
  INVX1 U1021 ( .A(n4784), .Y(n3914) );
  INVX1 U1022 ( .A(\data_in<5> ), .Y(n3919) );
  INVX1 U1023 ( .A(n2797), .Y(n3917) );
  INVX1 U1024 ( .A(\data_in<6> ), .Y(n3922) );
  INVX1 U1025 ( .A(n2839), .Y(n3920) );
  INVX1 U1026 ( .A(\data_in<7> ), .Y(n3925) );
  INVX1 U1027 ( .A(n4783), .Y(n3923) );
  INVX1 U1028 ( .A(\data_in<0> ), .Y(n3930) );
  INVX1 U1029 ( .A(n2690), .Y(n3928) );
  INVX1 U1030 ( .A(\data_in<1> ), .Y(n3933) );
  INVX1 U1031 ( .A(n2753), .Y(n3931) );
  INVX1 U1032 ( .A(\data_in<2> ), .Y(n3936) );
  INVX1 U1033 ( .A(n4782), .Y(n3934) );
  INVX1 U1034 ( .A(\data_in<3> ), .Y(n3939) );
  INVX1 U1035 ( .A(n4781), .Y(n3937) );
  INVX1 U1036 ( .A(\data_in<4> ), .Y(n3942) );
  INVX1 U1037 ( .A(n4780), .Y(n3940) );
  INVX1 U1038 ( .A(\data_in<5> ), .Y(n3945) );
  INVX1 U1039 ( .A(n4779), .Y(n3943) );
  INVX1 U1040 ( .A(\data_in<6> ), .Y(n3948) );
  INVX1 U1041 ( .A(n4778), .Y(n3946) );
  INVX1 U1042 ( .A(\data_in<7> ), .Y(n3951) );
  INVX1 U1043 ( .A(n2888), .Y(n3949) );
  INVX1 U1044 ( .A(\data_in<0> ), .Y(n3956) );
  INVX1 U1045 ( .A(n2691), .Y(n3954) );
  INVX1 U1046 ( .A(\data_in<1> ), .Y(n3959) );
  INVX1 U1047 ( .A(n2754), .Y(n3957) );
  INVX1 U1048 ( .A(\data_in<2> ), .Y(n3962) );
  INVX1 U1049 ( .A(n4777), .Y(n3960) );
  INVX1 U1050 ( .A(\data_in<3> ), .Y(n3965) );
  INVX1 U1051 ( .A(n4776), .Y(n3963) );
  INVX1 U1052 ( .A(\data_in<4> ), .Y(n3968) );
  INVX1 U1053 ( .A(n4775), .Y(n3966) );
  INVX1 U1054 ( .A(\data_in<5> ), .Y(n3971) );
  INVX1 U1055 ( .A(n4774), .Y(n3969) );
  INVX1 U1056 ( .A(\data_in<6> ), .Y(n3974) );
  INVX1 U1057 ( .A(n4773), .Y(n3972) );
  INVX1 U1058 ( .A(\data_in<7> ), .Y(n3977) );
  INVX1 U1059 ( .A(n2890), .Y(n3975) );
  INVX1 U1060 ( .A(\data_in<0> ), .Y(n3981) );
  INVX1 U1061 ( .A(n4772), .Y(n3979) );
  INVX1 U1062 ( .A(\data_in<1> ), .Y(n3984) );
  INVX1 U1063 ( .A(n4771), .Y(n3982) );
  INVX1 U1064 ( .A(\data_in<2> ), .Y(n3987) );
  INVX1 U1065 ( .A(n4770), .Y(n3985) );
  INVX1 U1066 ( .A(\data_in<3> ), .Y(n3990) );
  INVX1 U1067 ( .A(n4769), .Y(n3988) );
  INVX1 U1068 ( .A(\data_in<4> ), .Y(n3993) );
  INVX1 U1069 ( .A(n4768), .Y(n3991) );
  INVX1 U1070 ( .A(\data_in<5> ), .Y(n3996) );
  INVX1 U1071 ( .A(n4767), .Y(n3994) );
  INVX1 U1072 ( .A(\data_in<6> ), .Y(n3999) );
  INVX1 U1073 ( .A(n4766), .Y(n3997) );
  INVX1 U1074 ( .A(\data_in<7> ), .Y(n4002) );
  INVX1 U1075 ( .A(n4765), .Y(n4000) );
  INVX1 U1076 ( .A(\data_in<0> ), .Y(n4006) );
  INVX1 U1077 ( .A(n4764), .Y(n4004) );
  INVX1 U1078 ( .A(\data_in<1> ), .Y(n4009) );
  INVX1 U1079 ( .A(n4763), .Y(n4007) );
  INVX1 U1080 ( .A(\data_in<2> ), .Y(n4012) );
  INVX1 U1081 ( .A(n4762), .Y(n4010) );
  INVX1 U1082 ( .A(\data_in<3> ), .Y(n4015) );
  INVX1 U1083 ( .A(n4761), .Y(n4013) );
  INVX1 U1084 ( .A(\data_in<4> ), .Y(n4018) );
  INVX1 U1085 ( .A(n4760), .Y(n4016) );
  INVX1 U1086 ( .A(\data_in<5> ), .Y(n4021) );
  INVX1 U1087 ( .A(n4759), .Y(n4019) );
  INVX1 U1088 ( .A(\data_in<6> ), .Y(n4024) );
  INVX1 U1089 ( .A(n4758), .Y(n4022) );
  INVX1 U1090 ( .A(\data_in<7> ), .Y(n4027) );
  INVX1 U1091 ( .A(n4757), .Y(n4025) );
  INVX1 U1092 ( .A(\data_in<0> ), .Y(n4031) );
  INVX1 U1093 ( .A(n4756), .Y(n4029) );
  INVX1 U1094 ( .A(\data_in<1> ), .Y(n4034) );
  INVX1 U1095 ( .A(n4755), .Y(n4032) );
  INVX1 U1096 ( .A(\data_in<2> ), .Y(n4037) );
  INVX1 U1097 ( .A(n4754), .Y(n4035) );
  INVX1 U1098 ( .A(\data_in<3> ), .Y(n4040) );
  INVX1 U1099 ( .A(n4753), .Y(n4038) );
  INVX1 U1100 ( .A(\data_in<4> ), .Y(n4043) );
  INVX1 U1101 ( .A(n4752), .Y(n4041) );
  INVX1 U1102 ( .A(\data_in<5> ), .Y(n4046) );
  INVX1 U1103 ( .A(n4751), .Y(n4044) );
  INVX1 U1104 ( .A(\data_in<6> ), .Y(n4049) );
  INVX1 U1105 ( .A(n4750), .Y(n4047) );
  INVX1 U1106 ( .A(\data_in<7> ), .Y(n4052) );
  INVX1 U1107 ( .A(n4749), .Y(n4050) );
  INVX1 U1108 ( .A(\data_in<0> ), .Y(n4056) );
  INVX1 U1109 ( .A(n4748), .Y(n4054) );
  INVX1 U1110 ( .A(\data_in<1> ), .Y(n4059) );
  INVX1 U1111 ( .A(n4747), .Y(n4057) );
  INVX1 U1112 ( .A(\data_in<2> ), .Y(n4062) );
  INVX1 U1113 ( .A(n4746), .Y(n4060) );
  INVX1 U1114 ( .A(\data_in<3> ), .Y(n4065) );
  INVX1 U1115 ( .A(n4745), .Y(n4063) );
  INVX1 U1116 ( .A(\data_in<4> ), .Y(n4068) );
  INVX1 U1117 ( .A(n4744), .Y(n4066) );
  INVX1 U1118 ( .A(\data_in<5> ), .Y(n4071) );
  INVX1 U1119 ( .A(n4743), .Y(n4069) );
  INVX1 U1120 ( .A(\data_in<6> ), .Y(n4074) );
  INVX1 U1121 ( .A(n4742), .Y(n4072) );
  INVX1 U1122 ( .A(\data_in<7> ), .Y(n4077) );
  INVX1 U1123 ( .A(n4741), .Y(n4075) );
  INVX1 U1124 ( .A(\data_in<0> ), .Y(n4081) );
  INVX1 U1125 ( .A(n4740), .Y(n4079) );
  INVX1 U1126 ( .A(\data_in<1> ), .Y(n4084) );
  INVX1 U1127 ( .A(n4739), .Y(n4082) );
  INVX1 U1128 ( .A(\data_in<2> ), .Y(n4087) );
  INVX1 U1129 ( .A(n4738), .Y(n4085) );
  INVX1 U1130 ( .A(\data_in<3> ), .Y(n4090) );
  INVX1 U1131 ( .A(n4737), .Y(n4088) );
  INVX1 U1132 ( .A(\data_in<4> ), .Y(n4093) );
  INVX1 U1133 ( .A(n4736), .Y(n4091) );
  INVX1 U1134 ( .A(\data_in<5> ), .Y(n4096) );
  INVX1 U1135 ( .A(n4735), .Y(n4094) );
  INVX1 U1136 ( .A(\data_in<6> ), .Y(n4099) );
  INVX1 U1137 ( .A(n4734), .Y(n4097) );
  INVX1 U1138 ( .A(\data_in<7> ), .Y(n4102) );
  INVX1 U1139 ( .A(n4733), .Y(n4100) );
  INVX1 U1140 ( .A(\data_in<0> ), .Y(n4106) );
  INVX1 U1141 ( .A(n4732), .Y(n4104) );
  INVX1 U1142 ( .A(\data_in<1> ), .Y(n4109) );
  INVX1 U1143 ( .A(n4731), .Y(n4107) );
  INVX1 U1144 ( .A(\data_in<2> ), .Y(n4112) );
  INVX1 U1145 ( .A(n4730), .Y(n4110) );
  INVX1 U1146 ( .A(\data_in<3> ), .Y(n4115) );
  INVX1 U1147 ( .A(n4729), .Y(n4113) );
  INVX1 U1148 ( .A(\data_in<4> ), .Y(n4118) );
  INVX1 U1149 ( .A(n4728), .Y(n4116) );
  INVX1 U1150 ( .A(\data_in<5> ), .Y(n4121) );
  INVX1 U1151 ( .A(n4727), .Y(n4119) );
  INVX1 U1152 ( .A(\data_in<6> ), .Y(n4124) );
  INVX1 U1153 ( .A(n4726), .Y(n4122) );
  INVX1 U1154 ( .A(\data_in<7> ), .Y(n4127) );
  INVX1 U1155 ( .A(n4725), .Y(n4125) );
  INVX1 U1156 ( .A(\data_in<0> ), .Y(n4131) );
  INVX1 U1157 ( .A(n4724), .Y(n4129) );
  INVX1 U1158 ( .A(\data_in<1> ), .Y(n4134) );
  INVX1 U1159 ( .A(n4723), .Y(n4132) );
  INVX1 U1160 ( .A(\data_in<2> ), .Y(n4137) );
  INVX1 U1161 ( .A(n4722), .Y(n4135) );
  INVX1 U1162 ( .A(\data_in<3> ), .Y(n4140) );
  INVX1 U1163 ( .A(n4721), .Y(n4138) );
  INVX1 U1164 ( .A(\data_in<4> ), .Y(n4143) );
  INVX1 U1165 ( .A(n4720), .Y(n4141) );
  INVX1 U1166 ( .A(\data_in<5> ), .Y(n4146) );
  INVX1 U1167 ( .A(n4719), .Y(n4144) );
  INVX1 U1168 ( .A(\data_in<6> ), .Y(n4149) );
  INVX1 U1169 ( .A(n4718), .Y(n4147) );
  INVX1 U1170 ( .A(\data_in<7> ), .Y(n4152) );
  INVX1 U1171 ( .A(n4717), .Y(n4150) );
  INVX1 U1172 ( .A(\data_in<0> ), .Y(n4156) );
  INVX1 U1173 ( .A(n4716), .Y(n4154) );
  INVX1 U1174 ( .A(\data_in<1> ), .Y(n4159) );
  INVX1 U1175 ( .A(n4715), .Y(n4157) );
  INVX1 U1176 ( .A(\data_in<2> ), .Y(n4162) );
  INVX1 U1177 ( .A(n4714), .Y(n4160) );
  INVX1 U1178 ( .A(\data_in<3> ), .Y(n4165) );
  INVX1 U1179 ( .A(n4713), .Y(n4163) );
  INVX1 U1180 ( .A(\data_in<4> ), .Y(n4168) );
  INVX1 U1181 ( .A(n4712), .Y(n4166) );
  INVX1 U1182 ( .A(\data_in<5> ), .Y(n4171) );
  INVX1 U1183 ( .A(n4711), .Y(n4169) );
  INVX1 U1184 ( .A(\data_in<6> ), .Y(n4174) );
  INVX1 U1185 ( .A(n4710), .Y(n4172) );
  INVX1 U1186 ( .A(\data_in<7> ), .Y(n4177) );
  INVX1 U1187 ( .A(n4709), .Y(n4175) );
  INVX1 U1188 ( .A(\data_in<0> ), .Y(n4180) );
  INVX1 U1189 ( .A(n4708), .Y(n4178) );
  INVX1 U1190 ( .A(\data_in<1> ), .Y(n4183) );
  INVX1 U1191 ( .A(n4707), .Y(n4181) );
  INVX1 U1192 ( .A(\data_in<2> ), .Y(n4186) );
  INVX1 U1193 ( .A(n4706), .Y(n4184) );
  INVX1 U1194 ( .A(\data_in<3> ), .Y(n4189) );
  INVX1 U1195 ( .A(n4705), .Y(n4187) );
  INVX1 U1196 ( .A(\data_in<4> ), .Y(n4192) );
  INVX1 U1197 ( .A(n4704), .Y(n4190) );
  INVX1 U1198 ( .A(\data_in<5> ), .Y(n4195) );
  INVX1 U1199 ( .A(n4703), .Y(n4193) );
  INVX1 U1200 ( .A(\data_in<6> ), .Y(n4198) );
  INVX1 U1201 ( .A(n4702), .Y(n4196) );
  INVX1 U1202 ( .A(\data_in<7> ), .Y(n4201) );
  INVX1 U1203 ( .A(n4701), .Y(n4199) );
  INVX1 U1204 ( .A(\data_in<0> ), .Y(n4206) );
  INVX1 U1205 ( .A(n4700), .Y(n4204) );
  INVX1 U1206 ( .A(\data_in<1> ), .Y(n4209) );
  INVX1 U1207 ( .A(n4699), .Y(n4207) );
  INVX1 U1208 ( .A(\data_in<2> ), .Y(n4212) );
  INVX1 U1209 ( .A(n4698), .Y(n4210) );
  INVX1 U1210 ( .A(\data_in<3> ), .Y(n4215) );
  INVX1 U1211 ( .A(n4697), .Y(n4213) );
  INVX1 U1212 ( .A(\data_in<4> ), .Y(n4218) );
  INVX1 U1213 ( .A(n4696), .Y(n4216) );
  INVX1 U1214 ( .A(\data_in<5> ), .Y(n4221) );
  INVX1 U1215 ( .A(n4695), .Y(n4219) );
  INVX1 U1216 ( .A(\data_in<6> ), .Y(n4224) );
  INVX1 U1217 ( .A(n4694), .Y(n4222) );
  INVX1 U1218 ( .A(\data_in<7> ), .Y(n4227) );
  INVX1 U1219 ( .A(n4693), .Y(n4225) );
  INVX1 U1220 ( .A(\data_in<0> ), .Y(n4230) );
  INVX1 U1221 ( .A(n4692), .Y(n4228) );
  INVX1 U1222 ( .A(\data_in<1> ), .Y(n4233) );
  INVX1 U1223 ( .A(n4691), .Y(n4231) );
  INVX1 U1224 ( .A(\data_in<2> ), .Y(n4236) );
  INVX1 U1225 ( .A(n4690), .Y(n4234) );
  INVX1 U1226 ( .A(\data_in<3> ), .Y(n4239) );
  INVX1 U1227 ( .A(n4689), .Y(n4237) );
  INVX1 U1228 ( .A(\data_in<4> ), .Y(n4242) );
  INVX1 U1229 ( .A(n4688), .Y(n4240) );
  INVX1 U1230 ( .A(\data_in<5> ), .Y(n4245) );
  INVX1 U1231 ( .A(n4687), .Y(n4243) );
  INVX1 U1232 ( .A(\data_in<6> ), .Y(n4248) );
  INVX1 U1233 ( .A(n4686), .Y(n4246) );
  INVX1 U1234 ( .A(\data_in<7> ), .Y(n4251) );
  INVX1 U1235 ( .A(n4685), .Y(n4249) );
  INVX1 U1236 ( .A(\data_in<0> ), .Y(n4255) );
  INVX1 U1237 ( .A(n4684), .Y(n4253) );
  INVX1 U1238 ( .A(\data_in<1> ), .Y(n4258) );
  INVX1 U1239 ( .A(n4683), .Y(n4256) );
  INVX1 U1240 ( .A(\data_in<2> ), .Y(n4261) );
  INVX1 U1241 ( .A(n4682), .Y(n4259) );
  INVX1 U1242 ( .A(\data_in<3> ), .Y(n4264) );
  INVX1 U1243 ( .A(n4681), .Y(n4262) );
  INVX1 U1244 ( .A(\data_in<4> ), .Y(n4267) );
  INVX1 U1245 ( .A(n4680), .Y(n4265) );
  INVX1 U1246 ( .A(\data_in<5> ), .Y(n4270) );
  INVX1 U1247 ( .A(n4679), .Y(n4268) );
  INVX1 U1248 ( .A(\data_in<6> ), .Y(n4273) );
  INVX1 U1249 ( .A(n4678), .Y(n4271) );
  INVX1 U1250 ( .A(\data_in<7> ), .Y(n4276) );
  INVX1 U1251 ( .A(n4677), .Y(n4274) );
  INVX1 U1252 ( .A(\data_in<0> ), .Y(n4280) );
  INVX1 U1253 ( .A(n4676), .Y(n4278) );
  INVX1 U1254 ( .A(\data_in<1> ), .Y(n4283) );
  INVX1 U1255 ( .A(n4675), .Y(n4281) );
  INVX1 U1256 ( .A(\data_in<2> ), .Y(n4286) );
  INVX1 U1257 ( .A(n4674), .Y(n4284) );
  INVX1 U1258 ( .A(\data_in<3> ), .Y(n4289) );
  INVX1 U1259 ( .A(n4673), .Y(n4287) );
  INVX1 U1260 ( .A(\data_in<4> ), .Y(n4292) );
  INVX1 U1261 ( .A(n4672), .Y(n4290) );
  INVX1 U1262 ( .A(\data_in<5> ), .Y(n4295) );
  INVX1 U1263 ( .A(n4671), .Y(n4293) );
  INVX1 U1264 ( .A(\data_in<6> ), .Y(n4298) );
  INVX1 U1265 ( .A(n4670), .Y(n4296) );
  INVX1 U1266 ( .A(\data_in<7> ), .Y(n4301) );
  INVX1 U1267 ( .A(n4669), .Y(n4299) );
  INVX1 U1268 ( .A(\data_in<0> ), .Y(n4305) );
  INVX1 U1269 ( .A(n4668), .Y(n4303) );
  INVX1 U1270 ( .A(\data_in<1> ), .Y(n4308) );
  INVX1 U1271 ( .A(n4667), .Y(n4306) );
  INVX1 U1272 ( .A(\data_in<2> ), .Y(n4311) );
  INVX1 U1273 ( .A(n4666), .Y(n4309) );
  INVX1 U1274 ( .A(\data_in<3> ), .Y(n4314) );
  INVX1 U1275 ( .A(n4665), .Y(n4312) );
  INVX1 U1276 ( .A(\data_in<4> ), .Y(n4317) );
  INVX1 U1277 ( .A(n4664), .Y(n4315) );
  INVX1 U1278 ( .A(\data_in<5> ), .Y(n4320) );
  INVX1 U1279 ( .A(n4663), .Y(n4318) );
  INVX1 U1280 ( .A(\data_in<6> ), .Y(n4323) );
  INVX1 U1281 ( .A(n4662), .Y(n4321) );
  INVX1 U1282 ( .A(\data_in<7> ), .Y(n4326) );
  INVX1 U1283 ( .A(n4661), .Y(n4324) );
  INVX1 U1284 ( .A(\data_in<0> ), .Y(n4330) );
  INVX1 U1285 ( .A(n4660), .Y(n4328) );
  INVX1 U1286 ( .A(\data_in<1> ), .Y(n4333) );
  INVX1 U1287 ( .A(n4659), .Y(n4331) );
  INVX1 U1288 ( .A(\data_in<2> ), .Y(n4336) );
  INVX1 U1289 ( .A(n4658), .Y(n4334) );
  INVX1 U1290 ( .A(\data_in<3> ), .Y(n4339) );
  INVX1 U1291 ( .A(n4657), .Y(n4337) );
  INVX1 U1292 ( .A(\data_in<4> ), .Y(n4342) );
  INVX1 U1293 ( .A(n4656), .Y(n4340) );
  INVX1 U1294 ( .A(\data_in<5> ), .Y(n4345) );
  INVX1 U1295 ( .A(n4655), .Y(n4343) );
  INVX1 U1296 ( .A(\data_in<6> ), .Y(n4348) );
  INVX1 U1297 ( .A(n4654), .Y(n4346) );
  INVX1 U1298 ( .A(\data_in<7> ), .Y(n4351) );
  INVX1 U1299 ( .A(n4653), .Y(n4349) );
  INVX1 U1300 ( .A(\data_in<0> ), .Y(n4355) );
  INVX1 U1301 ( .A(n4652), .Y(n4353) );
  INVX1 U1302 ( .A(\data_in<1> ), .Y(n4358) );
  INVX1 U1303 ( .A(n4651), .Y(n4356) );
  INVX1 U1304 ( .A(\data_in<2> ), .Y(n4361) );
  INVX1 U1305 ( .A(n4650), .Y(n4359) );
  INVX1 U1306 ( .A(\data_in<3> ), .Y(n4364) );
  INVX1 U1307 ( .A(n4649), .Y(n4362) );
  INVX1 U1308 ( .A(\data_in<4> ), .Y(n4367) );
  INVX1 U1309 ( .A(n4648), .Y(n4365) );
  INVX1 U1310 ( .A(\data_in<5> ), .Y(n4370) );
  INVX1 U1311 ( .A(n4647), .Y(n4368) );
  INVX1 U1312 ( .A(\data_in<6> ), .Y(n4373) );
  INVX1 U1313 ( .A(n4646), .Y(n4371) );
  INVX1 U1314 ( .A(\data_in<7> ), .Y(n4376) );
  INVX1 U1315 ( .A(n4645), .Y(n4374) );
  INVX1 U1316 ( .A(\data_in<0> ), .Y(n4380) );
  INVX1 U1317 ( .A(n4644), .Y(n4378) );
  INVX1 U1318 ( .A(\data_in<1> ), .Y(n4383) );
  INVX1 U1319 ( .A(n4643), .Y(n4381) );
  INVX1 U1320 ( .A(\data_in<2> ), .Y(n4386) );
  INVX1 U1321 ( .A(n4642), .Y(n4384) );
  INVX1 U1322 ( .A(\data_in<3> ), .Y(n4389) );
  INVX1 U1323 ( .A(n4641), .Y(n4387) );
  INVX1 U1324 ( .A(\data_in<4> ), .Y(n4392) );
  INVX1 U1325 ( .A(n4640), .Y(n4390) );
  INVX1 U1326 ( .A(\data_in<5> ), .Y(n4395) );
  INVX1 U1327 ( .A(n4639), .Y(n4393) );
  INVX1 U1328 ( .A(\data_in<6> ), .Y(n4398) );
  INVX1 U1329 ( .A(n4638), .Y(n4396) );
  INVX1 U1330 ( .A(\data_in<7> ), .Y(n4401) );
  INVX1 U1331 ( .A(n4637), .Y(n4399) );
  INVX1 U1332 ( .A(\data_in<0> ), .Y(n4405) );
  INVX1 U1333 ( .A(n4636), .Y(n4403) );
  INVX1 U1334 ( .A(\data_in<1> ), .Y(n4408) );
  INVX1 U1335 ( .A(n4635), .Y(n4406) );
  INVX1 U1336 ( .A(\data_in<2> ), .Y(n4411) );
  INVX1 U1337 ( .A(n4634), .Y(n4409) );
  INVX1 U1338 ( .A(\data_in<3> ), .Y(n4414) );
  INVX1 U1339 ( .A(n4633), .Y(n4412) );
  INVX1 U1340 ( .A(\data_in<4> ), .Y(n4417) );
  INVX1 U1341 ( .A(n4632), .Y(n4415) );
  INVX1 U1342 ( .A(\data_in<5> ), .Y(n4420) );
  INVX1 U1343 ( .A(n4631), .Y(n4418) );
  INVX1 U1344 ( .A(\data_in<6> ), .Y(n4423) );
  INVX1 U1345 ( .A(n4630), .Y(n4421) );
  INVX1 U1346 ( .A(\data_in<7> ), .Y(n4426) );
  INVX1 U1347 ( .A(n4629), .Y(n4424) );
  INVX1 U1348 ( .A(\data_in<0> ), .Y(n4429) );
  INVX1 U1349 ( .A(n2709), .Y(n4427) );
  INVX1 U1350 ( .A(\data_in<1> ), .Y(n4432) );
  INVX1 U1351 ( .A(n2764), .Y(n4430) );
  INVX1 U1352 ( .A(\data_in<2> ), .Y(n4435) );
  INVX1 U1353 ( .A(n4628), .Y(n4433) );
  INVX1 U1354 ( .A(\data_in<3> ), .Y(n4438) );
  INVX1 U1355 ( .A(n4627), .Y(n4436) );
  INVX1 U1356 ( .A(\data_in<4> ), .Y(n4441) );
  INVX1 U1357 ( .A(n4626), .Y(n4439) );
  INVX1 U1358 ( .A(\data_in<5> ), .Y(n4444) );
  INVX1 U1359 ( .A(n4625), .Y(n4442) );
  INVX1 U1360 ( .A(\data_in<6> ), .Y(n4447) );
  INVX1 U1361 ( .A(n4624), .Y(n4445) );
  INVX1 U1362 ( .A(\data_in<7> ), .Y(n4450) );
  INVX1 U1363 ( .A(n2901), .Y(n4448) );
  INVX1 U1364 ( .A(\data_in<0> ), .Y(n4454) );
  INVX1 U1365 ( .A(n4623), .Y(n4452) );
  INVX1 U1366 ( .A(\data_in<1> ), .Y(n4457) );
  INVX1 U1367 ( .A(n4622), .Y(n4455) );
  INVX1 U1368 ( .A(\data_in<2> ), .Y(n4460) );
  INVX1 U1369 ( .A(n4621), .Y(n4458) );
  INVX1 U1370 ( .A(\data_in<3> ), .Y(n4463) );
  INVX1 U1371 ( .A(n4620), .Y(n4461) );
  INVX1 U1372 ( .A(\data_in<4> ), .Y(n4466) );
  INVX1 U1373 ( .A(n4619), .Y(n4464) );
  INVX1 U1374 ( .A(\data_in<5> ), .Y(n4469) );
  INVX1 U1375 ( .A(n4618), .Y(n4467) );
  INVX1 U1376 ( .A(\data_in<6> ), .Y(n4472) );
  INVX1 U1377 ( .A(n4617), .Y(n4470) );
  INVX1 U1378 ( .A(\data_in<7> ), .Y(n4475) );
  INVX1 U1379 ( .A(n4616), .Y(n4473) );
  INVX1 U1380 ( .A(\data_in<0> ), .Y(n4479) );
  INVX1 U1381 ( .A(n4615), .Y(n4477) );
  INVX1 U1382 ( .A(\data_in<1> ), .Y(n4482) );
  INVX1 U1383 ( .A(n2763), .Y(n4480) );
  INVX1 U1384 ( .A(\data_in<2> ), .Y(n4485) );
  INVX1 U1385 ( .A(n4614), .Y(n4483) );
  INVX1 U1386 ( .A(\data_in<3> ), .Y(n4488) );
  INVX1 U1387 ( .A(n4613), .Y(n4486) );
  INVX1 U1388 ( .A(\data_in<4> ), .Y(n4491) );
  INVX1 U1389 ( .A(n4612), .Y(n4489) );
  INVX1 U1390 ( .A(\data_in<5> ), .Y(n4494) );
  INVX1 U1391 ( .A(n4611), .Y(n4492) );
  INVX1 U1392 ( .A(\data_in<6> ), .Y(n4497) );
  INVX1 U1393 ( .A(n4610), .Y(n4495) );
  INVX1 U1394 ( .A(\data_in<7> ), .Y(n4500) );
  INVX1 U1395 ( .A(n2900), .Y(n4498) );
  INVX1 U1396 ( .A(\data_in<0> ), .Y(n4504) );
  INVX1 U1397 ( .A(n4609), .Y(n4502) );
  INVX1 U1398 ( .A(\data_in<1> ), .Y(n4507) );
  INVX1 U1399 ( .A(n4608), .Y(n4505) );
  INVX1 U1400 ( .A(\data_in<2> ), .Y(n4510) );
  INVX1 U1401 ( .A(n4607), .Y(n4508) );
  INVX1 U1402 ( .A(\data_in<3> ), .Y(n4513) );
  INVX1 U1403 ( .A(n4606), .Y(n4511) );
  INVX1 U1404 ( .A(\data_in<4> ), .Y(n4516) );
  INVX1 U1405 ( .A(n4605), .Y(n4514) );
  INVX1 U1406 ( .A(\data_in<5> ), .Y(n4519) );
  INVX1 U1407 ( .A(n4604), .Y(n4517) );
  INVX1 U1408 ( .A(\data_in<6> ), .Y(n4522) );
  INVX1 U1409 ( .A(n4603), .Y(n4520) );
  INVX1 U1410 ( .A(\data_in<7> ), .Y(n4525) );
  INVX1 U1411 ( .A(n4602), .Y(n4523) );
  INVX1 U1412 ( .A(\data_in<0> ), .Y(n4529) );
  INVX1 U1413 ( .A(n2712), .Y(n4527) );
  INVX1 U1414 ( .A(\data_in<1> ), .Y(n4532) );
  INVX1 U1415 ( .A(n2769), .Y(n4530) );
  INVX1 U1416 ( .A(\data_in<2> ), .Y(n4535) );
  INVX1 U1417 ( .A(n4601), .Y(n4533) );
  INVX1 U1418 ( .A(\data_in<3> ), .Y(n4538) );
  INVX1 U1419 ( .A(n4600), .Y(n4536) );
  INVX1 U1420 ( .A(\data_in<4> ), .Y(n4541) );
  INVX1 U1421 ( .A(n4599), .Y(n4539) );
  INVX1 U1422 ( .A(\data_in<5> ), .Y(n4544) );
  INVX1 U1423 ( .A(n4598), .Y(n4542) );
  INVX1 U1424 ( .A(\data_in<6> ), .Y(n4547) );
  INVX1 U1425 ( .A(n4597), .Y(n4545) );
  INVX1 U1426 ( .A(\data_in<7> ), .Y(n4550) );
  INVX1 U1427 ( .A(n2906), .Y(n4548) );
  INVX1 U1428 ( .A(\data_in<0> ), .Y(n4555) );
  INVX1 U1429 ( .A(\data_in<1> ), .Y(n4558) );
  INVX1 U1430 ( .A(\data_in<2> ), .Y(n4561) );
  INVX1 U1431 ( .A(\data_in<3> ), .Y(n4564) );
  INVX1 U1432 ( .A(\data_in<4> ), .Y(n4567) );
  INVX1 U1433 ( .A(\data_in<5> ), .Y(n4570) );
  INVX1 U1434 ( .A(\data_in<6> ), .Y(n4573) );
  INVX1 U1435 ( .A(\data_in<7> ), .Y(n4577) );
  INVX1 U1436 ( .A(\data_in<8> ), .Y(n4578) );
  INVX1 U1437 ( .A(\data_in<9> ), .Y(n4579) );
  INVX1 U1438 ( .A(\data_in<10> ), .Y(n4580) );
  INVX1 U1439 ( .A(\mem<0><2> ), .Y(n4591) );
  INVX1 U1440 ( .A(\data_in<11> ), .Y(n4581) );
  INVX1 U1441 ( .A(\mem<0><3> ), .Y(n4590) );
  INVX1 U1442 ( .A(\data_in<12> ), .Y(n4582) );
  INVX1 U1443 ( .A(\mem<0><4> ), .Y(n4589) );
  INVX1 U1444 ( .A(\data_in<13> ), .Y(n4583) );
  INVX1 U1445 ( .A(\mem<0><5> ), .Y(n4588) );
  INVX1 U1446 ( .A(\data_in<14> ), .Y(n4584) );
  INVX1 U1447 ( .A(\mem<0><6> ), .Y(n4587) );
  INVX1 U1448 ( .A(\data_in<15> ), .Y(n4585) );
  INVX4 U1449 ( .A(n2545), .Y(n2548) );
  INVX8 U1450 ( .A(n2545), .Y(n2546) );
  INVX4 U1451 ( .A(n451), .Y(n2549) );
  INVX1 U1452 ( .A(n451), .Y(n2560) );
  AND2X1 U1453 ( .A(n2626), .B(n1169), .Y(n1072) );
  AND2X1 U1454 ( .A(n444), .B(n1175), .Y(n1075) );
  AND2X1 U1455 ( .A(n2630), .B(n739), .Y(n1213) );
  INVX1 U1456 ( .A(n2544), .Y(n1455) );
  INVX1 U1457 ( .A(n2542), .Y(n478) );
  INVX1 U1458 ( .A(n2546), .Y(n513) );
  AND2X2 U1459 ( .A(n1465), .B(n545), .Y(n3) );
  INVX1 U1460 ( .A(n2546), .Y(n452) );
  AND2X1 U1461 ( .A(n2629), .B(n721), .Y(n1195) );
  AND2X1 U1462 ( .A(n2629), .B(n735), .Y(n1209) );
  AND2X1 U1463 ( .A(n2629), .B(n737), .Y(n1211) );
  AND2X1 U1464 ( .A(n1294), .B(n785), .Y(n1259) );
  AND2X1 U1465 ( .A(n2631), .B(n787), .Y(n1261) );
  AND2X1 U1466 ( .A(n2630), .B(n691), .Y(n1165) );
  AND2X1 U1467 ( .A(n2628), .B(n693), .Y(n1167) );
  AND2X1 U1468 ( .A(n2628), .B(n697), .Y(n1171) );
  AND2X1 U1469 ( .A(n2628), .B(n699), .Y(n1173) );
  AND2X1 U1470 ( .A(n2628), .B(n705), .Y(n1179) );
  AND2X1 U1471 ( .A(n2628), .B(n707), .Y(n1181) );
  AND2X1 U1472 ( .A(n2629), .B(n717), .Y(n1191) );
  AND2X1 U1473 ( .A(n2629), .B(n723), .Y(n1197) );
  AND2X1 U1474 ( .A(n2629), .B(n725), .Y(n1199) );
  AND2X1 U1475 ( .A(n2629), .B(n729), .Y(n1203) );
  AND2X1 U1476 ( .A(n2629), .B(n731), .Y(n1205) );
  AND2X1 U1477 ( .A(n2629), .B(n733), .Y(n1207) );
  AND2X1 U1478 ( .A(n2630), .B(n741), .Y(n1215) );
  AND2X1 U1479 ( .A(n2630), .B(n745), .Y(n1219) );
  AND2X1 U1480 ( .A(n2630), .B(n747), .Y(n1221) );
  AND2X1 U1481 ( .A(n2630), .B(n749), .Y(n1223) );
  AND2X1 U1482 ( .A(n2630), .B(n753), .Y(n1227) );
  AND2X1 U1483 ( .A(n2630), .B(n755), .Y(n1229) );
  AND2X1 U1484 ( .A(n2630), .B(n757), .Y(n1231) );
  AND2X1 U1485 ( .A(n2630), .B(n759), .Y(n1233) );
  AND2X1 U1486 ( .A(n2631), .B(n761), .Y(n1235) );
  AND2X1 U1487 ( .A(n2631), .B(n763), .Y(n1237) );
  AND2X1 U1488 ( .A(n2631), .B(n765), .Y(n1239) );
  AND2X1 U1489 ( .A(n2631), .B(n767), .Y(n1241) );
  AND2X1 U1490 ( .A(n2631), .B(n769), .Y(n1243) );
  AND2X1 U1491 ( .A(n2631), .B(n773), .Y(n1247) );
  AND2X1 U1492 ( .A(n2631), .B(n781), .Y(n1255) );
  AND2X1 U1493 ( .A(n1294), .B(n783), .Y(n1257) );
  AND2X1 U1494 ( .A(n1294), .B(n789), .Y(n1263) );
  AND2X1 U1495 ( .A(n1294), .B(n795), .Y(n1269) );
  AND2X1 U1496 ( .A(n1294), .B(n799), .Y(n1273) );
  AND2X1 U1497 ( .A(n2630), .B(n743), .Y(n1217) );
  AND2X1 U1498 ( .A(n2631), .B(n771), .Y(n1245) );
  AND2X1 U1499 ( .A(n1294), .B(n791), .Y(n1265) );
  AND2X1 U1500 ( .A(n2628), .B(n711), .Y(n1185) );
  AND2X1 U1501 ( .A(n2628), .B(n695), .Y(n1169) );
  AND2X1 U1502 ( .A(n2628), .B(n701), .Y(n1175) );
  AND2X1 U1503 ( .A(n2630), .B(n751), .Y(n1225) );
  AND2X1 U1504 ( .A(n1294), .B(n793), .Y(n1267) );
  AND2X1 U1505 ( .A(n1294), .B(n797), .Y(n1271) );
  AND2X1 U1506 ( .A(n2628), .B(n801), .Y(n1275) );
  INVX1 U1507 ( .A(\mem<38><3> ), .Y(n556) );
  BUFX2 U1508 ( .A(n394), .Y(n2623) );
  INVX4 U1509 ( .A(n2540), .Y(n2541) );
  INVX1 U1510 ( .A(n1512), .Y(n78) );
  INVX1 U1511 ( .A(\mem<4><0> ), .Y(n4615) );
  AND2X1 U1512 ( .A(n3268), .B(n3267), .Y(n1080) );
  INVX1 U1513 ( .A(\mem<63><7> ), .Y(n2882) );
  INVX1 U1514 ( .A(\mem<63><1> ), .Y(n2747) );
  INVX1 U1515 ( .A(\mem<63><0> ), .Y(n2684) );
  INVX1 U1516 ( .A(\mem<0><0> ), .Y(n2700) );
  INVX1 U1517 ( .A(\mem<0><1> ), .Y(n2758) );
  INVX1 U1518 ( .A(\mem<0><7> ), .Y(n2894) );
  INVX1 U1519 ( .A(\mem<28><0> ), .Y(n2702) );
  INVX1 U1520 ( .A(\mem<26><0> ), .Y(n2690) );
  INVX1 U1521 ( .A(\mem<62><5> ), .Y(n2789) );
  INVX1 U1522 ( .A(\mem<62><6> ), .Y(n2831) );
  INVX1 U1523 ( .A(\mem<61><0> ), .Y(n2686) );
  INVX1 U1524 ( .A(\mem<60><5> ), .Y(n2791) );
  INVX1 U1525 ( .A(\mem<60><6> ), .Y(n2833) );
  INVX1 U1526 ( .A(n2783), .Y(n536) );
  INVX1 U1527 ( .A(\mem<32><0> ), .Y(n2679) );
  INVX1 U1528 ( .A(\mem<32><1> ), .Y(n2743) );
  INVX1 U1529 ( .A(\mem<32><7> ), .Y(n2878) );
  INVX1 U1530 ( .A(\mem<28><7> ), .Y(n2896) );
  INVX1 U1531 ( .A(\mem<26><7> ), .Y(n2888) );
  INVX1 U1532 ( .A(\mem<6><1> ), .Y(n2764) );
  INVX1 U1533 ( .A(\mem<6><7> ), .Y(n2901) );
  INVX1 U1534 ( .A(\mem<4><1> ), .Y(n2763) );
  INVX1 U1535 ( .A(\mem<4><7> ), .Y(n2900) );
  INVX1 U1536 ( .A(\mem<2><0> ), .Y(n2712) );
  INVX1 U1537 ( .A(\mem<2><7> ), .Y(n2906) );
  INVX1 U1538 ( .A(\mem<1><1> ), .Y(n2768) );
  INVX1 U1539 ( .A(\mem<1><7> ), .Y(n2905) );
  INVX1 U1540 ( .A(\mem<1><0> ), .Y(n2711) );
  INVX1 U1541 ( .A(\mem<39><3> ), .Y(n557) );
  INVX1 U1542 ( .A(\mem<61><7> ), .Y(n2884) );
  INVX1 U1543 ( .A(\mem<59><1> ), .Y(n2742) );
  INVX1 U1544 ( .A(\mem<59><7> ), .Y(n2877) );
  INVX1 U1545 ( .A(\mem<57><5> ), .Y(n2785) );
  INVX1 U1546 ( .A(\mem<57><6> ), .Y(n2827) );
  INVX1 U1547 ( .A(\mem<29><5> ), .Y(n2795) );
  INVX1 U1548 ( .A(\mem<29><6> ), .Y(n2837) );
  INVX1 U1549 ( .A(\mem<27><5> ), .Y(n2797) );
  INVX1 U1550 ( .A(\mem<27><6> ), .Y(n2839) );
  INVX1 U1551 ( .A(\mem<26><1> ), .Y(n2753) );
  INVX1 U1552 ( .A(\mem<25><7> ), .Y(n2890) );
  INVX1 U1553 ( .A(\mem<6><0> ), .Y(n2709) );
  INVX1 U1554 ( .A(\mem<2><1> ), .Y(n2769) );
  INVX1 U1555 ( .A(\mem<61><1> ), .Y(n2749) );
  INVX1 U1556 ( .A(\mem<25><0> ), .Y(n2691) );
  INVX1 U1557 ( .A(\mem<25><1> ), .Y(n2754) );
  INVX1 U1558 ( .A(\mem<1><2> ), .Y(n4596) );
  INVX1 U1559 ( .A(\mem<57><2> ), .Y(n5015) );
  INVX1 U1560 ( .A(\mem<1><3> ), .Y(n4595) );
  INVX1 U1561 ( .A(\mem<57><3> ), .Y(n5014) );
  INVX1 U1562 ( .A(\mem<1><4> ), .Y(n4594) );
  INVX1 U1563 ( .A(\mem<57><4> ), .Y(n5013) );
  INVX1 U1564 ( .A(\mem<52><4> ), .Y(n4975) );
  INVX1 U1565 ( .A(\mem<25><2> ), .Y(n4777) );
  INVX1 U1566 ( .A(\mem<41><2> ), .Y(n4889) );
  INVX1 U1567 ( .A(\mem<30><3> ), .Y(n4805) );
  INVX1 U1568 ( .A(\mem<25><3> ), .Y(n4776) );
  INVX1 U1569 ( .A(\mem<41><3> ), .Y(n4888) );
  INVX1 U1570 ( .A(\mem<32><3> ), .Y(n4820) );
  INVX1 U1571 ( .A(\mem<25><4> ), .Y(n4775) );
  INVX1 U1572 ( .A(\mem<22><4> ), .Y(n4752) );
  INVX1 U1573 ( .A(\mem<41><4> ), .Y(n4887) );
  INVX1 U1574 ( .A(\mem<12><2> ), .Y(n4674) );
  INVX1 U1575 ( .A(\mem<14><2> ), .Y(n4690) );
  INVX1 U1576 ( .A(\mem<8><2> ), .Y(n4642) );
  INVX1 U1577 ( .A(\mem<10><2> ), .Y(n4658) );
  INVX1 U1578 ( .A(\mem<4><2> ), .Y(n4614) );
  INVX1 U1579 ( .A(\mem<6><2> ), .Y(n4628) );
  INVX1 U1580 ( .A(\mem<2><2> ), .Y(n4601) );
  INVX1 U1581 ( .A(\mem<60><2> ), .Y(n5034) );
  INVX1 U1582 ( .A(\mem<62><2> ), .Y(n5045) );
  INVX1 U1583 ( .A(\mem<58><2> ), .Y(n5022) );
  INVX1 U1584 ( .A(\mem<52><2> ), .Y(n4977) );
  INVX1 U1585 ( .A(\mem<54><2> ), .Y(n4993) );
  INVX1 U1586 ( .A(\mem<48><2> ), .Y(n4945) );
  INVX1 U1587 ( .A(\mem<50><2> ), .Y(n4961) );
  INVX1 U1588 ( .A(\mem<12><3> ), .Y(n4673) );
  INVX1 U1589 ( .A(\mem<14><3> ), .Y(n4689) );
  INVX1 U1590 ( .A(\mem<8><3> ), .Y(n4641) );
  INVX1 U1591 ( .A(\mem<10><3> ), .Y(n4657) );
  INVX1 U1592 ( .A(\mem<4><3> ), .Y(n4613) );
  INVX1 U1593 ( .A(\mem<6><3> ), .Y(n4627) );
  INVX1 U1594 ( .A(\mem<2><3> ), .Y(n4600) );
  INVX1 U1595 ( .A(\mem<60><3> ), .Y(n5033) );
  INVX1 U1596 ( .A(\mem<62><3> ), .Y(n5044) );
  INVX1 U1597 ( .A(\mem<58><3> ), .Y(n5021) );
  INVX1 U1598 ( .A(\mem<52><3> ), .Y(n4976) );
  INVX1 U1599 ( .A(\mem<54><3> ), .Y(n4992) );
  INVX1 U1600 ( .A(\mem<48><3> ), .Y(n4944) );
  INVX1 U1601 ( .A(\mem<50><3> ), .Y(n4960) );
  INVX1 U1602 ( .A(\mem<12><4> ), .Y(n4672) );
  INVX1 U1603 ( .A(\mem<14><4> ), .Y(n4688) );
  INVX1 U1604 ( .A(\mem<8><4> ), .Y(n4640) );
  INVX1 U1605 ( .A(\mem<10><4> ), .Y(n4656) );
  INVX1 U1606 ( .A(\mem<4><4> ), .Y(n4612) );
  INVX1 U1607 ( .A(\mem<6><4> ), .Y(n4626) );
  INVX1 U1608 ( .A(\mem<2><4> ), .Y(n4599) );
  INVX1 U1609 ( .A(\mem<60><4> ), .Y(n5032) );
  INVX1 U1610 ( .A(\mem<62><4> ), .Y(n5043) );
  INVX1 U1611 ( .A(\mem<58><4> ), .Y(n5020) );
  INVX1 U1612 ( .A(\mem<54><4> ), .Y(n4991) );
  INVX1 U1613 ( .A(\mem<48><4> ), .Y(n4943) );
  INVX1 U1614 ( .A(\mem<50><4> ), .Y(n4959) );
  INVX1 U1615 ( .A(\mem<28><2> ), .Y(n4793) );
  INVX1 U1616 ( .A(\mem<30><2> ), .Y(n4806) );
  INVX1 U1617 ( .A(\mem<26><2> ), .Y(n4782) );
  INVX1 U1618 ( .A(\mem<20><2> ), .Y(n4738) );
  INVX1 U1619 ( .A(\mem<22><2> ), .Y(n4754) );
  INVX1 U1620 ( .A(\mem<16><2> ), .Y(n4706) );
  INVX1 U1621 ( .A(\mem<18><2> ), .Y(n4722) );
  INVX1 U1622 ( .A(\mem<44><2> ), .Y(n4913) );
  INVX1 U1623 ( .A(\mem<46><2> ), .Y(n4929) );
  INVX1 U1624 ( .A(\mem<42><2> ), .Y(n4897) );
  INVX1 U1625 ( .A(\mem<36><2> ), .Y(n4851) );
  INVX1 U1626 ( .A(\mem<38><2> ), .Y(n4866) );
  INVX1 U1627 ( .A(\mem<32><2> ), .Y(n4821) );
  INVX1 U1628 ( .A(\mem<34><2> ), .Y(n4835) );
  INVX1 U1629 ( .A(\mem<28><3> ), .Y(n4792) );
  INVX1 U1630 ( .A(\mem<26><3> ), .Y(n4781) );
  INVX1 U1631 ( .A(\mem<20><3> ), .Y(n4737) );
  INVX1 U1632 ( .A(\mem<22><3> ), .Y(n4753) );
  INVX1 U1633 ( .A(\mem<16><3> ), .Y(n4705) );
  INVX1 U1634 ( .A(\mem<18><3> ), .Y(n4721) );
  INVX1 U1635 ( .A(\mem<44><3> ), .Y(n4912) );
  INVX1 U1636 ( .A(\mem<46><3> ), .Y(n4928) );
  INVX1 U1637 ( .A(\mem<42><3> ), .Y(n4896) );
  INVX1 U1638 ( .A(\mem<36><3> ), .Y(n4850) );
  INVX1 U1639 ( .A(\mem<34><3> ), .Y(n4834) );
  INVX1 U1640 ( .A(\mem<28><4> ), .Y(n4791) );
  INVX1 U1641 ( .A(\mem<30><4> ), .Y(n4804) );
  INVX1 U1642 ( .A(\mem<26><4> ), .Y(n4780) );
  INVX1 U1643 ( .A(\mem<20><4> ), .Y(n4736) );
  INVX1 U1644 ( .A(\mem<16><4> ), .Y(n4704) );
  INVX1 U1645 ( .A(\mem<18><4> ), .Y(n4720) );
  INVX1 U1646 ( .A(\mem<44><4> ), .Y(n4911) );
  INVX1 U1647 ( .A(\mem<46><4> ), .Y(n4927) );
  INVX1 U1648 ( .A(\mem<42><4> ), .Y(n4895) );
  INVX1 U1649 ( .A(\mem<36><4> ), .Y(n4849) );
  INVX1 U1650 ( .A(\mem<38><4> ), .Y(n4865) );
  INVX1 U1651 ( .A(\mem<32><4> ), .Y(n4819) );
  INVX1 U1652 ( .A(\mem<34><4> ), .Y(n4833) );
  INVX1 U1653 ( .A(n430), .Y(n4) );
  INVX1 U1654 ( .A(n4), .Y(n5) );
  AND2X2 U1655 ( .A(n2962), .B(n2610), .Y(n6) );
  INVX1 U1656 ( .A(n3572), .Y(n7) );
  NOR3X1 U1657 ( .A(n347), .B(n360), .C(n110), .Y(n8) );
  INVX2 U1658 ( .A(n8), .Y(n2726) );
  INVX4 U1659 ( .A(n370), .Y(n435) );
  AND2X2 U1660 ( .A(n282), .B(n272), .Y(n59) );
  INVX1 U1661 ( .A(n576), .Y(n9) );
  AND2X2 U1662 ( .A(n3875), .B(n3879), .Y(n2760) );
  INVX2 U1663 ( .A(n395), .Y(n3875) );
  INVX1 U1664 ( .A(n4794), .Y(n3879) );
  INVX1 U1665 ( .A(n2698), .Y(n10) );
  INVX1 U1666 ( .A(n10), .Y(n11) );
  INVX1 U1667 ( .A(n367), .Y(n12) );
  AND2X2 U1668 ( .A(n231), .B(n309), .Y(n13) );
  AND2X2 U1669 ( .A(\mem<9><1> ), .B(n438), .Y(n14) );
  INVX1 U1670 ( .A(\addr<6> ), .Y(n15) );
  INVX1 U1671 ( .A(n399), .Y(n16) );
  INVX1 U1672 ( .A(n3522), .Y(n17) );
  INVX1 U1673 ( .A(n1515), .Y(n18) );
  INVX1 U1674 ( .A(n18), .Y(n19) );
  INVX1 U1675 ( .A(N181), .Y(n20) );
  INVX1 U1676 ( .A(n1437), .Y(n21) );
  INVX4 U1677 ( .A(n564), .Y(n534) );
  INVX1 U1678 ( .A(N180), .Y(n1466) );
  OR2X2 U1679 ( .A(n33), .B(n50), .Y(n22) );
  INVX1 U1680 ( .A(n1504), .Y(n23) );
  INVX1 U1681 ( .A(n23), .Y(n24) );
  INVX1 U1682 ( .A(n70), .Y(n25) );
  INVX1 U1683 ( .A(\addr<8> ), .Y(n2715) );
  INVX1 U1684 ( .A(N181), .Y(n26) );
  INVX1 U1685 ( .A(n26), .Y(n27) );
  INVX1 U1686 ( .A(n35), .Y(n28) );
  INVX4 U1687 ( .A(n455), .Y(n1471) );
  INVX1 U1688 ( .A(n15), .Y(n29) );
  INVX1 U1689 ( .A(n1431), .Y(n30) );
  INVX1 U1690 ( .A(n2652), .Y(n31) );
  INVX1 U1691 ( .A(n1439), .Y(n32) );
  INVX1 U1692 ( .A(n463), .Y(n33) );
  INVX1 U1693 ( .A(n42), .Y(n34) );
  INVX1 U1694 ( .A(N182), .Y(n35) );
  INVX1 U1695 ( .A(n35), .Y(n36) );
  INVX1 U1696 ( .A(\addr<11> ), .Y(n37) );
  INVX1 U1697 ( .A(n37), .Y(n38) );
  INVX1 U1698 ( .A(\addr<6> ), .Y(n39) );
  INVX1 U1699 ( .A(n39), .Y(n40) );
  INVX1 U1700 ( .A(n384), .Y(n41) );
  INVX1 U1701 ( .A(N180), .Y(n42) );
  INVX1 U1702 ( .A(n42), .Y(n43) );
  AND2X2 U1703 ( .A(n1454), .B(n45), .Y(n44) );
  AND2X2 U1704 ( .A(n1465), .B(n545), .Y(n45) );
  INVX4 U1705 ( .A(n2617), .Y(n46) );
  INVX1 U1706 ( .A(n2617), .Y(n4501) );
  OR2X2 U1707 ( .A(n1473), .B(n29), .Y(n47) );
  AND2X2 U1708 ( .A(n41), .B(n1454), .Y(n48) );
  INVX1 U1709 ( .A(\addr<12> ), .Y(n49) );
  INVX1 U1710 ( .A(n49), .Y(n50) );
  AND2X2 U1711 ( .A(n62), .B(n1509), .Y(n2663) );
  AND2X2 U1712 ( .A(n392), .B(n581), .Y(n51) );
  BUFX2 U1713 ( .A(n1466), .Y(n448) );
  OR2X2 U1714 ( .A(n2565), .B(n579), .Y(n52) );
  OR2X2 U1715 ( .A(n2585), .B(n2877), .Y(n53) );
  INVX1 U1716 ( .A(n53), .Y(n54) );
  INVX1 U1717 ( .A(n22), .Y(n55) );
  INVX1 U1718 ( .A(n1502), .Y(n56) );
  OR2X2 U1719 ( .A(N182), .B(n88), .Y(n57) );
  AND2X2 U1720 ( .A(n271), .B(n71), .Y(n58) );
  INVX1 U1721 ( .A(n2632), .Y(n475) );
  INVX4 U1722 ( .A(n2560), .Y(n2561) );
  AND2X2 U1723 ( .A(n61), .B(n527), .Y(n60) );
  INVX1 U1724 ( .A(n60), .Y(n109) );
  INVX1 U1725 ( .A(n2708), .Y(n61) );
  INVX1 U1726 ( .A(n411), .Y(n2613) );
  INVX1 U1727 ( .A(\addr<6> ), .Y(n62) );
  AND2X2 U1728 ( .A(n1445), .B(\mem<35><5> ), .Y(n1470) );
  INVX1 U1729 ( .A(n399), .Y(n63) );
  INVX1 U1730 ( .A(n382), .Y(n64) );
  INVX4 U1731 ( .A(n408), .Y(n439) );
  AND2X2 U1732 ( .A(n2698), .B(n72), .Y(n65) );
  INVX1 U1733 ( .A(n78), .Y(n66) );
  INVX1 U1734 ( .A(n78), .Y(n67) );
  INVX1 U1735 ( .A(n1513), .Y(n503) );
  AND2X2 U1736 ( .A(N179), .B(N178), .Y(n68) );
  INVX4 U1737 ( .A(N179), .Y(n2635) );
  INVX1 U1738 ( .A(N178), .Y(n564) );
  INVX1 U1739 ( .A(n1287), .Y(n433) );
  AND2X2 U1740 ( .A(n212), .B(n298), .Y(n69) );
  OR2X2 U1741 ( .A(n373), .B(n52), .Y(n70) );
  INVX1 U1742 ( .A(n70), .Y(n1449) );
  NOR3X1 U1743 ( .A(n348), .B(n361), .C(n119), .Y(n71) );
  INVX4 U1744 ( .A(n402), .Y(n436) );
  INVX1 U1745 ( .A(n1285), .Y(n72) );
  AND2X2 U1746 ( .A(n104), .B(n291), .Y(n84) );
  AND2X2 U1747 ( .A(n283), .B(n273), .Y(n73) );
  OR2X2 U1748 ( .A(n4501), .B(n4615), .Y(n450) );
  AND2X2 U1749 ( .A(n43), .B(n20), .Y(n74) );
  AND2X2 U1750 ( .A(n2584), .B(\mem<59><0> ), .Y(n75) );
  AND2X2 U1751 ( .A(n275), .B(n285), .Y(n76) );
  INVX1 U1752 ( .A(n109), .Y(n1498) );
  INVX1 U1753 ( .A(n1292), .Y(n77) );
  INVX1 U1754 ( .A(n78), .Y(n79) );
  AND2X1 U1755 ( .A(n2587), .B(n2723), .Y(n1484) );
  INVX1 U1756 ( .A(n528), .Y(n80) );
  INVX1 U1757 ( .A(n561), .Y(n81) );
  INVX1 U1758 ( .A(n81), .Y(n82) );
  AND2X2 U1759 ( .A(n2699), .B(n65), .Y(n561) );
  AND2X2 U1760 ( .A(n244), .B(n324), .Y(n83) );
  AND2X2 U1761 ( .A(n155), .B(n185), .Y(n274) );
  INVX1 U1762 ( .A(n34), .Y(n2636) );
  OR2X2 U1763 ( .A(n57), .B(n90), .Y(n85) );
  INVX1 U1764 ( .A(n1279), .Y(n2723) );
  AND2X2 U1765 ( .A(n274), .B(n284), .Y(n86) );
  INVX1 U1766 ( .A(n47), .Y(n87) );
  INVX1 U1767 ( .A(N181), .Y(n88) );
  INVX1 U1768 ( .A(n2718), .Y(n89) );
  INVX1 U1769 ( .A(n1466), .Y(n90) );
  OR2X2 U1770 ( .A(n201), .B(n92), .Y(n91) );
  OR2X2 U1771 ( .A(n200), .B(n1136), .Y(n92) );
  OR2X2 U1772 ( .A(n471), .B(n94), .Y(n93) );
  OR2X2 U1773 ( .A(n365), .B(n364), .Y(n94) );
  AND2X2 U1774 ( .A(n199), .B(n2802), .Y(n95) );
  AND2X2 U1775 ( .A(n499), .B(n500), .Y(n96) );
  OR2X2 U1776 ( .A(n2683), .B(n2696), .Y(n97) );
  INVX1 U1777 ( .A(\addr<9> ), .Y(n2716) );
  AND2X2 U1778 ( .A(n2658), .B(n2657), .Y(n98) );
  INVX1 U1779 ( .A(n98), .Y(n99) );
  OR2X2 U1780 ( .A(n99), .B(n290), .Y(n100) );
  INVX1 U1781 ( .A(n100), .Y(n101) );
  AND2X2 U1782 ( .A(n2673), .B(n2672), .Y(n102) );
  INVX1 U1783 ( .A(n102), .Y(n103) );
  AND2X2 U1784 ( .A(n197), .B(n195), .Y(n104) );
  AND2X2 U1785 ( .A(n36), .B(n1479), .Y(n105) );
  AND2X2 U1786 ( .A(n2682), .B(n2681), .Y(n106) );
  OR2X2 U1787 ( .A(n1030), .B(n293), .Y(n107) );
  AND2X2 U1788 ( .A(n2705), .B(n2704), .Y(n108) );
  OR2X2 U1789 ( .A(n211), .B(n295), .Y(n110) );
  AND2X2 U1790 ( .A(n2730), .B(n2731), .Y(n111) );
  INVX1 U1791 ( .A(n111), .Y(n112) );
  OR2X2 U1792 ( .A(n112), .B(n297), .Y(n113) );
  INVX1 U1793 ( .A(n113), .Y(n114) );
  AND2X2 U1794 ( .A(n2741), .B(n2740), .Y(n115) );
  INVX1 U1795 ( .A(n115), .Y(n116) );
  AND2X2 U1796 ( .A(n2762), .B(n2761), .Y(n117) );
  INVX1 U1797 ( .A(n117), .Y(n118) );
  OR2X2 U1798 ( .A(n222), .B(n302), .Y(n119) );
  OR2X2 U1799 ( .A(n252), .B(n332), .Y(n120) );
  INVX1 U1800 ( .A(n120), .Y(n121) );
  OR2X2 U1801 ( .A(n256), .B(n427), .Y(n122) );
  INVX1 U1802 ( .A(n122), .Y(n123) );
  OR2X2 U1803 ( .A(n258), .B(n334), .Y(n124) );
  INVX1 U1804 ( .A(n124), .Y(n125) );
  OR2X2 U1805 ( .A(n254), .B(n336), .Y(n126) );
  INVX1 U1806 ( .A(n126), .Y(n127) );
  AND2X2 U1807 ( .A(n2881), .B(n2880), .Y(n128) );
  INVX1 U1808 ( .A(n128), .Y(n129) );
  AND2X2 U1809 ( .A(n2899), .B(n2898), .Y(n130) );
  INVX1 U1810 ( .A(n130), .Y(n131) );
  OR2X2 U1811 ( .A(n264), .B(n340), .Y(n132) );
  INVX1 U1812 ( .A(n132), .Y(n133) );
  OR2X2 U1813 ( .A(n262), .B(n286), .Y(n134) );
  INVX1 U1814 ( .A(n134), .Y(n135) );
  OR2X2 U1815 ( .A(n563), .B(n562), .Y(n136) );
  INVX1 U1816 ( .A(n136), .Y(n137) );
  INVX1 U1817 ( .A(n138), .Y(n139) );
  OR2X2 U1818 ( .A(n1029), .B(n1062), .Y(n140) );
  INVX1 U1819 ( .A(n140), .Y(n141) );
  OR2X2 U1820 ( .A(n203), .B(n1065), .Y(n142) );
  INVX1 U1821 ( .A(n142), .Y(n143) );
  OR2X2 U1822 ( .A(n214), .B(n425), .Y(n144) );
  INVX1 U1823 ( .A(n144), .Y(n145) );
  OR2X2 U1824 ( .A(n218), .B(n300), .Y(n146) );
  INVX1 U1825 ( .A(n146), .Y(n147) );
  OR2X2 U1826 ( .A(n224), .B(n304), .Y(n148) );
  INVX1 U1827 ( .A(n148), .Y(n149) );
  OR2X2 U1828 ( .A(n230), .B(n288), .Y(n150) );
  INVX1 U1829 ( .A(n150), .Y(n151) );
  OR2X2 U1830 ( .A(n235), .B(n313), .Y(n152) );
  INVX1 U1831 ( .A(n152), .Y(n153) );
  OR2X2 U1832 ( .A(n317), .B(n239), .Y(n154) );
  INVX1 U1833 ( .A(n154), .Y(n155) );
  OR2X2 U1834 ( .A(n243), .B(n321), .Y(n156) );
  INVX1 U1835 ( .A(n156), .Y(n157) );
  OR2X2 U1836 ( .A(n248), .B(n328), .Y(n158) );
  INVX1 U1837 ( .A(n158), .Y(n159) );
  OR2X2 U1838 ( .A(n1032), .B(n1067), .Y(n160) );
  INVX1 U1839 ( .A(n160), .Y(n161) );
  OR2X2 U1840 ( .A(n129), .B(n338), .Y(n162) );
  INVX1 U1841 ( .A(n162), .Y(n163) );
  OR2X2 U1842 ( .A(n453), .B(n454), .Y(n164) );
  INVX1 U1843 ( .A(n164), .Y(n165) );
  OR2X2 U1844 ( .A(n1469), .B(n1470), .Y(n166) );
  INVX1 U1845 ( .A(n166), .Y(n167) );
  AND2X2 U1846 ( .A(\mem<34><6> ), .B(n2586), .Y(n168) );
  INVX1 U1847 ( .A(n168), .Y(n169) );
  OR2X2 U1848 ( .A(n209), .B(n1063), .Y(n170) );
  INVX1 U1849 ( .A(n170), .Y(n171) );
  OR2X2 U1850 ( .A(n216), .B(n116), .Y(n172) );
  INVX1 U1851 ( .A(n172), .Y(n173) );
  OR2X2 U1852 ( .A(n220), .B(n118), .Y(n174) );
  INVX1 U1853 ( .A(n174), .Y(n175) );
  OR2X2 U1854 ( .A(n226), .B(n306), .Y(n176) );
  INVX1 U1855 ( .A(n176), .Y(n177) );
  OR2X2 U1856 ( .A(n228), .B(n308), .Y(n178) );
  INVX1 U1857 ( .A(n178), .Y(n179) );
  OR2X2 U1858 ( .A(n233), .B(n311), .Y(n180) );
  INVX1 U1859 ( .A(n180), .Y(n181) );
  OR2X2 U1860 ( .A(n237), .B(n315), .Y(n182) );
  INVX1 U1861 ( .A(n182), .Y(n183) );
  OR2X2 U1862 ( .A(n241), .B(n319), .Y(n184) );
  INVX1 U1863 ( .A(n184), .Y(n185) );
  OR2X2 U1864 ( .A(n91), .B(n323), .Y(n186) );
  INVX1 U1865 ( .A(n186), .Y(n187) );
  OR2X2 U1866 ( .A(n246), .B(n326), .Y(n188) );
  INVX1 U1867 ( .A(n188), .Y(n189) );
  OR2X2 U1868 ( .A(n250), .B(n330), .Y(n190) );
  INVX1 U1869 ( .A(n190), .Y(n191) );
  OR2X2 U1870 ( .A(n260), .B(n131), .Y(n192) );
  INVX1 U1871 ( .A(n192), .Y(n193) );
  OR2X2 U1872 ( .A(n207), .B(n103), .Y(n194) );
  INVX1 U1873 ( .A(n194), .Y(n195) );
  OR2X2 U1874 ( .A(n205), .B(n423), .Y(n196) );
  INVX1 U1875 ( .A(n196), .Y(n197) );
  AND2X2 U1876 ( .A(n3798), .B(\mem<31><5> ), .Y(n198) );
  INVX1 U1877 ( .A(n198), .Y(n199) );
  INVX1 U1878 ( .A(n2843), .Y(n200) );
  INVX1 U1879 ( .A(n2844), .Y(n201) );
  AND2X2 U1880 ( .A(n2727), .B(n165), .Y(n202) );
  INVX1 U1881 ( .A(n202), .Y(n203) );
  AND2X2 U1882 ( .A(n2666), .B(n2665), .Y(n204) );
  INVX1 U1883 ( .A(n204), .Y(n205) );
  AND2X2 U1884 ( .A(n2671), .B(n2670), .Y(n206) );
  INVX1 U1885 ( .A(n206), .Y(n207) );
  AND2X2 U1886 ( .A(n2694), .B(n2693), .Y(n208) );
  INVX1 U1887 ( .A(n208), .Y(n209) );
  AND2X2 U1888 ( .A(n2720), .B(n2721), .Y(n210) );
  INVX1 U1889 ( .A(n210), .Y(n211) );
  AND2X2 U1890 ( .A(n143), .B(n114), .Y(n212) );
  AND2X2 U1891 ( .A(n2735), .B(n2734), .Y(n213) );
  INVX1 U1892 ( .A(n213), .Y(n214) );
  AND2X2 U1893 ( .A(n2739), .B(n2738), .Y(n215) );
  INVX1 U1894 ( .A(n215), .Y(n216) );
  AND2X2 U1895 ( .A(n2746), .B(n2745), .Y(n217) );
  INVX1 U1896 ( .A(n217), .Y(n218) );
  AND2X2 U1897 ( .A(n2757), .B(n2756), .Y(n219) );
  INVX1 U1898 ( .A(n219), .Y(n220) );
  AND2X2 U1899 ( .A(n2773), .B(n2772), .Y(n221) );
  INVX1 U1900 ( .A(n221), .Y(n222) );
  AND2X2 U1901 ( .A(n137), .B(n2776), .Y(n223) );
  INVX1 U1902 ( .A(n223), .Y(n224) );
  AND2X2 U1903 ( .A(n2782), .B(n2781), .Y(n225) );
  INVX1 U1904 ( .A(n225), .Y(n226) );
  AND2X2 U1906 ( .A(n2788), .B(n2787), .Y(n227) );
  INVX1 U1907 ( .A(n227), .Y(n228) );
  AND2X2 U1908 ( .A(n2800), .B(n2799), .Y(n229) );
  INVX1 U1909 ( .A(n229), .Y(n230) );
  AND2X2 U1910 ( .A(n2803), .B(n167), .Y(n231) );
  AND2X2 U1911 ( .A(n2806), .B(n2807), .Y(n232) );
  INVX1 U1912 ( .A(n232), .Y(n233) );
  AND2X2 U1913 ( .A(n2810), .B(n2811), .Y(n234) );
  INVX1 U1914 ( .A(n234), .Y(n235) );
  AND2X2 U1915 ( .A(n2816), .B(n2817), .Y(n236) );
  INVX1 U1916 ( .A(n236), .Y(n237) );
  AND2X2 U1917 ( .A(n2821), .B(n2820), .Y(n238) );
  INVX1 U1918 ( .A(n238), .Y(n239) );
  AND2X2 U1919 ( .A(n2825), .B(n2824), .Y(n240) );
  INVX1 U1920 ( .A(n240), .Y(n241) );
  AND2X2 U1921 ( .A(n2836), .B(n2835), .Y(n242) );
  INVX1 U1922 ( .A(n242), .Y(n243) );
  AND2X2 U1923 ( .A(n2848), .B(n2847), .Y(n244) );
  AND2X2 U1924 ( .A(n2852), .B(n2851), .Y(n245) );
  INVX1 U1925 ( .A(n245), .Y(n246) );
  AND2X2 U1926 ( .A(n2854), .B(n2853), .Y(n247) );
  INVX1 U1927 ( .A(n247), .Y(n248) );
  AND2X2 U1928 ( .A(n2860), .B(n2859), .Y(n249) );
  INVX1 U1929 ( .A(n249), .Y(n250) );
  AND2X2 U1930 ( .A(n2866), .B(n2865), .Y(n251) );
  INVX1 U1931 ( .A(n251), .Y(n252) );
  AND2X2 U1932 ( .A(n161), .B(n121), .Y(n253) );
  INVX1 U1933 ( .A(n253), .Y(n254) );
  AND2X2 U1934 ( .A(n2870), .B(n2869), .Y(n255) );
  INVX1 U1935 ( .A(n255), .Y(n256) );
  AND2X2 U1936 ( .A(n2874), .B(n2873), .Y(n257) );
  INVX1 U1937 ( .A(n257), .Y(n258) );
  AND2X2 U1938 ( .A(n2893), .B(n2892), .Y(n259) );
  INVX1 U1939 ( .A(n259), .Y(n260) );
  INVX1 U1940 ( .A(n261), .Y(n262) );
  AND2X2 U1941 ( .A(n2910), .B(n2909), .Y(n263) );
  INVX1 U1942 ( .A(n263), .Y(n264) );
  AND2X2 U1943 ( .A(n450), .B(n819), .Y(n265) );
  INVX1 U1944 ( .A(n265), .Y(n266) );
  AND2X2 U1945 ( .A(n40), .B(N182), .Y(n267) );
  INVX1 U1946 ( .A(n267), .Y(n268) );
  AND2X2 U1947 ( .A(n575), .B(n171), .Y(n269) );
  INVX1 U1948 ( .A(n269), .Y(n270) );
  AND2X2 U1949 ( .A(n147), .B(n175), .Y(n271) );
  AND2X2 U1950 ( .A(n151), .B(n179), .Y(n272) );
  AND2X2 U1951 ( .A(n153), .B(n183), .Y(n273) );
  AND2X2 U1952 ( .A(n159), .B(n191), .Y(n275) );
  AND2X2 U1953 ( .A(n2655), .B(n2654), .Y(n276) );
  INVX1 U1954 ( .A(n276), .Y(n277) );
  AND2X2 U1955 ( .A(n1493), .B(n2663), .Y(n278) );
  INVX1 U1956 ( .A(n278), .Y(n279) );
  AND2X2 U1957 ( .A(n74), .B(n2669), .Y(n280) );
  INVX1 U1958 ( .A(n280), .Y(n281) );
  AND2X2 U1959 ( .A(n149), .B(n177), .Y(n282) );
  AND2X2 U1960 ( .A(n13), .B(n181), .Y(n283) );
  AND2X2 U1961 ( .A(n157), .B(n187), .Y(n284) );
  AND2X2 U1962 ( .A(n83), .B(n189), .Y(n285) );
  BUFX2 U1963 ( .A(n2913), .Y(n286) );
  AND2X2 U1964 ( .A(n2801), .B(n95), .Y(n287) );
  INVX1 U1965 ( .A(n287), .Y(n288) );
  AND2X2 U1966 ( .A(n2660), .B(n2659), .Y(n289) );
  INVX1 U1967 ( .A(n289), .Y(n290) );
  AND2X2 U1968 ( .A(n141), .B(n101), .Y(n291) );
  AND2X2 U1969 ( .A(n2689), .B(n2688), .Y(n292) );
  INVX1 U1970 ( .A(n292), .Y(n293) );
  AND2X2 U1971 ( .A(n2724), .B(n2725), .Y(n294) );
  INVX1 U1972 ( .A(n294), .Y(n295) );
  AND2X2 U1973 ( .A(n2733), .B(n2732), .Y(n296) );
  INVX1 U1974 ( .A(n296), .Y(n297) );
  AND2X2 U1975 ( .A(n145), .B(n173), .Y(n298) );
  AND2X2 U1976 ( .A(n2752), .B(n2751), .Y(n299) );
  INVX1 U1977 ( .A(n299), .Y(n300) );
  AND2X2 U1978 ( .A(n2775), .B(n2774), .Y(n301) );
  INVX1 U1979 ( .A(n301), .Y(n302) );
  AND2X2 U1980 ( .A(n2778), .B(n2777), .Y(n303) );
  INVX1 U1981 ( .A(n303), .Y(n304) );
  AND2X2 U1982 ( .A(n2780), .B(n2779), .Y(n305) );
  INVX1 U1983 ( .A(n305), .Y(n306) );
  AND2X2 U1984 ( .A(n2794), .B(n2793), .Y(n307) );
  INVX1 U1985 ( .A(n307), .Y(n308) );
  AND2X2 U1986 ( .A(n2805), .B(n2804), .Y(n309) );
  AND2X2 U1987 ( .A(n2809), .B(n2808), .Y(n310) );
  INVX1 U1988 ( .A(n310), .Y(n311) );
  AND2X2 U1989 ( .A(n2813), .B(n2812), .Y(n312) );
  INVX1 U1990 ( .A(n312), .Y(n313) );
  AND2X2 U1991 ( .A(n2814), .B(n2815), .Y(n314) );
  INVX1 U1992 ( .A(n314), .Y(n315) );
  AND2X2 U1993 ( .A(n2819), .B(n2818), .Y(n316) );
  INVX1 U1994 ( .A(n316), .Y(n317) );
  AND2X2 U1995 ( .A(n2822), .B(n2823), .Y(n318) );
  INVX1 U1996 ( .A(n318), .Y(n319) );
  AND2X2 U1997 ( .A(n2829), .B(n2830), .Y(n320) );
  INVX1 U1998 ( .A(n320), .Y(n321) );
  AND2X2 U1999 ( .A(n2841), .B(n2842), .Y(n322) );
  INVX1 U2000 ( .A(n322), .Y(n323) );
  AND2X2 U2001 ( .A(n2846), .B(n2845), .Y(n324) );
  AND2X2 U2002 ( .A(n2849), .B(n2850), .Y(n325) );
  INVX1 U2003 ( .A(n325), .Y(n326) );
  AND2X2 U2004 ( .A(n2856), .B(n2855), .Y(n327) );
  INVX1 U2005 ( .A(n327), .Y(n328) );
  AND2X2 U2006 ( .A(n2857), .B(n2858), .Y(n329) );
  INVX1 U2007 ( .A(n329), .Y(n330) );
  AND2X2 U2008 ( .A(n2868), .B(n2867), .Y(n331) );
  INVX1 U2009 ( .A(n331), .Y(n332) );
  AND2X2 U2010 ( .A(n2876), .B(n2875), .Y(n333) );
  INVX1 U2011 ( .A(n333), .Y(n334) );
  AND2X2 U2012 ( .A(n123), .B(n125), .Y(n335) );
  INVX1 U2013 ( .A(n335), .Y(n336) );
  AND2X2 U2014 ( .A(n2887), .B(n2886), .Y(n337) );
  INVX1 U2015 ( .A(n337), .Y(n338) );
  AND2X2 U2016 ( .A(n2912), .B(n2911), .Y(n339) );
  INVX1 U2017 ( .A(n339), .Y(n340) );
  OR2X2 U2018 ( .A(n397), .B(n2690), .Y(n341) );
  INVX1 U2019 ( .A(n341), .Y(n342) );
  OR2X2 U2020 ( .A(n93), .B(n2742), .Y(n343) );
  INVX1 U2021 ( .A(n343), .Y(n344) );
  OR2X2 U2022 ( .A(n542), .B(n2753), .Y(n345) );
  INVX1 U2023 ( .A(n345), .Y(n346) );
  OR2X2 U2024 ( .A(n266), .B(n2710), .Y(n347) );
  OR2X1 U2025 ( .A(n2766), .B(n2765), .Y(n348) );
  OR2X1 U2026 ( .A(n2903), .B(n2902), .Y(n349) );
  INVX1 U2027 ( .A(n349), .Y(n350) );
  BUFX2 U2028 ( .A(n2645), .Y(n351) );
  INVX1 U2029 ( .A(n351), .Y(n352) );
  INVX1 U2030 ( .A(n351), .Y(n353) );
  BUFX2 U2031 ( .A(n2648), .Y(n354) );
  INVX1 U2032 ( .A(n354), .Y(n355) );
  INVX1 U2033 ( .A(n354), .Y(n356) );
  AND2X2 U2034 ( .A(n568), .B(n1497), .Y(n357) );
  OR2X2 U2037 ( .A(n270), .B(n2726), .Y(n358) );
  INVX1 U2038 ( .A(n358), .Y(n359) );
  OR2X2 U2039 ( .A(n2714), .B(n2713), .Y(n360) );
  OR2X2 U2040 ( .A(n2770), .B(n2771), .Y(n361) );
  OR2X2 U2041 ( .A(n2908), .B(n2907), .Y(n362) );
  INVX1 U2042 ( .A(n362), .Y(n363) );
  INVX1 U2043 ( .A(n45), .Y(n364) );
  INVX1 U2044 ( .A(n1476), .Y(n365) );
  AND2X2 U2045 ( .A(n485), .B(n2594), .Y(n366) );
  INVX1 U2046 ( .A(n366), .Y(n367) );
  INVX1 U2047 ( .A(n366), .Y(n368) );
  AND2X2 U2048 ( .A(n2723), .B(n48), .Y(n369) );
  INVX1 U2049 ( .A(n369), .Y(n370) );
  INVX1 U2050 ( .A(n369), .Y(n371) );
  AND2X2 U2051 ( .A(n391), .B(n581), .Y(n372) );
  INVX1 U2052 ( .A(n372), .Y(n373) );
  AND2X2 U2053 ( .A(n2661), .B(n2662), .Y(n374) );
  OR2X2 U2054 ( .A(n2643), .B(n2644), .Y(n375) );
  INVX1 U2055 ( .A(n375), .Y(n376) );
  AND2X2 U2056 ( .A(n356), .B(n2611), .Y(n377) );
  INVX1 U2058 ( .A(n377), .Y(n378) );
  AND2X2 U2059 ( .A(n355), .B(n48), .Y(n379) );
  AND2X2 U2060 ( .A(n51), .B(n3), .Y(n380) );
  INVX1 U2061 ( .A(n380), .Y(n381) );
  INVX1 U2062 ( .A(n380), .Y(n382) );
  AND2X2 U2063 ( .A(n356), .B(n1498), .Y(n383) );
  OR2X2 U2064 ( .A(n2656), .B(n277), .Y(n384) );
  INVX1 U2065 ( .A(n384), .Y(n385) );
  INVX1 U2066 ( .A(n384), .Y(n386) );
  OR2X2 U2067 ( .A(n2706), .B(n281), .Y(n387) );
  INVX1 U2068 ( .A(n387), .Y(n388) );
  INVX1 U2069 ( .A(n387), .Y(n389) );
  OR2X2 U2070 ( .A(n2664), .B(n279), .Y(n390) );
  INVX1 U2071 ( .A(n390), .Y(n391) );
  INVX1 U2072 ( .A(n390), .Y(n392) );
  AND2X1 U2073 ( .A(enable), .B(n2638), .Y(n393) );
  INVX1 U2074 ( .A(n393), .Y(n394) );
  BUFX2 U2075 ( .A(n3900), .Y(n395) );
  BUFX2 U2076 ( .A(n3013), .Y(n396) );
  BUFX2 U2077 ( .A(n3952), .Y(n397) );
  BUFX2 U2080 ( .A(n3848), .Y(n398) );
  BUFX2 U2081 ( .A(n3823), .Y(n399) );
  AND2X2 U2082 ( .A(n353), .B(n51), .Y(n400) );
  INVX1 U2083 ( .A(n400), .Y(n401) );
  INVX1 U2084 ( .A(n400), .Y(n402) );
  AND2X2 U2085 ( .A(n355), .B(n2587), .Y(n403) );
  INVX1 U2086 ( .A(n403), .Y(n404) );
  AND2X2 U2087 ( .A(n569), .B(n2611), .Y(n405) );
  AND2X2 U2088 ( .A(n438), .B(n48), .Y(n406) );
  INVX1 U2089 ( .A(n406), .Y(n407) );
  INVX1 U2090 ( .A(n406), .Y(n408) );
  BUFX2 U2091 ( .A(n1450), .Y(n409) );
  AND2X2 U2092 ( .A(n2723), .B(n540), .Y(n410) );
  INVX1 U2093 ( .A(n410), .Y(n411) );
  AND2X2 U2094 ( .A(n2962), .B(n2594), .Y(n412) );
  AND2X2 U2095 ( .A(n2722), .B(n2962), .Y(n413) );
  AND2X2 U2096 ( .A(n438), .B(n2587), .Y(n414) );
  BUFX2 U2097 ( .A(n3166), .Y(n415) );
  BUFX2 U2098 ( .A(n3874), .Y(n416) );
  MUX2X1 U2099 ( .B(n1590), .A(n1593), .S(n417), .Y(n1605) );
  MUX2X1 U2101 ( .B(n1524), .A(n1521), .S(n2548), .Y(n1538) );
  INVX1 U2102 ( .A(n559), .Y(n418) );
  INVX4 U2103 ( .A(n547), .Y(n2569) );
  AND2X2 U2104 ( .A(n489), .B(n545), .Y(n419) );
  AND2X2 U2105 ( .A(\mem<8><0> ), .B(n490), .Y(n420) );
  INVX1 U2106 ( .A(n420), .Y(n421) );
  INVX2 U2107 ( .A(n550), .Y(n3901) );
  AND2X2 U2108 ( .A(n2668), .B(n2667), .Y(n422) );
  INVX1 U2109 ( .A(n422), .Y(n423) );
  AND2X2 U2110 ( .A(n2736), .B(n2737), .Y(n424) );
  INVX1 U2111 ( .A(n424), .Y(n425) );
  AND2X2 U2112 ( .A(n2872), .B(n2871), .Y(n426) );
  INVX1 U2113 ( .A(n426), .Y(n427) );
  INVX1 U2114 ( .A(n2599), .Y(n428) );
  INVX1 U2115 ( .A(n3064), .Y(n2597) );
  AND2X2 U2116 ( .A(n376), .B(n438), .Y(n429) );
  AND2X2 U2117 ( .A(n558), .B(n438), .Y(n430) );
  AND2X2 U2118 ( .A(n1465), .B(n68), .Y(n431) );
  INVX1 U2119 ( .A(n398), .Y(n432) );
  INVX2 U2120 ( .A(n398), .Y(n2600) );
  INVX1 U2123 ( .A(n399), .Y(n3798) );
  INVX1 U2124 ( .A(n4476), .Y(n434) );
  INVX1 U2125 ( .A(n371), .Y(n2593) );
  INVX1 U2126 ( .A(n401), .Y(n1520) );
  INVX1 U2127 ( .A(n404), .Y(n437) );
  AND2X2 U2128 ( .A(n1465), .B(n511), .Y(n438) );
  INVX1 U2129 ( .A(n407), .Y(n3747) );
  INVX1 U2130 ( .A(n1289), .Y(n440) );
  INVX1 U2131 ( .A(n3090), .Y(n441) );
  INVX1 U2132 ( .A(n441), .Y(n442) );
  INVX1 U2133 ( .A(n441), .Y(n443) );
  INVX1 U2134 ( .A(n3141), .Y(n444) );
  INVX1 U2135 ( .A(n3978), .Y(n445) );
  INVX1 U2136 ( .A(n445), .Y(n446) );
  INVX1 U2137 ( .A(n445), .Y(n447) );
  MUX2X1 U2138 ( .B(n2358), .A(n2355), .S(n2547), .Y(n2369) );
  INVX4 U2139 ( .A(n492), .Y(n493) );
  INVX1 U2140 ( .A(n3926), .Y(n1483) );
  INVX1 U2141 ( .A(n522), .Y(n449) );
  INVX1 U2142 ( .A(n555), .Y(n1742) );
  BUFX2 U2144 ( .A(N178), .Y(n451) );
  INVX1 U2145 ( .A(N178), .Y(n2633) );
  MUX2X1 U2146 ( .B(n1772), .A(n1771), .S(n2551), .Y(n1770) );
  MUX2X1 U2147 ( .B(\mem<21><5> ), .A(\mem<20><5> ), .S(n1465), .Y(n2391) );
  MUX2X1 U2148 ( .B(\mem<45><1> ), .A(\mem<44><1> ), .S(n578), .Y(n1607) );
  MUX2X1 U2149 ( .B(\mem<25><1> ), .A(\mem<24><1> ), .S(n493), .Y(n1625) );
  MUX2X1 U2150 ( .B(n2467), .A(n2470), .S(n452), .Y(n2474) );
  MUX2X1 U2151 ( .B(\mem<51><0> ), .A(\mem<50><0> ), .S(n2564), .Y(n1535) );
  MUX2X1 U2152 ( .B(\mem<9><0> ), .A(\mem<8><0> ), .S(n494), .Y(n1574) );
  AND2X2 U2153 ( .A(\mem<16><1> ), .B(n1513), .Y(n453) );
  AND2X2 U2154 ( .A(n376), .B(n14), .Y(n454) );
  MUX2X1 U2155 ( .B(\mem<11><0> ), .A(\mem<10><0> ), .S(n1471), .Y(n1575) );
  INVX1 U2156 ( .A(n368), .Y(n543) );
  INVX2 U2157 ( .A(n1434), .Y(n455) );
  INVX2 U2158 ( .A(n1434), .Y(n2582) );
  INVX1 U2159 ( .A(n1291), .Y(n456) );
  AND2X2 U2160 ( .A(n558), .B(n485), .Y(n457) );
  AND2X2 U2161 ( .A(n2612), .B(n485), .Y(n458) );
  INVX1 U2162 ( .A(n492), .Y(n459) );
  INVX1 U2163 ( .A(n487), .Y(n460) );
  INVX1 U2164 ( .A(n4078), .Y(n461) );
  INVX1 U2165 ( .A(n2605), .Y(n462) );
  MUX2X1 U2166 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n2567), .Y(n1557) );
  MUX2X1 U2167 ( .B(n2407), .A(n2406), .S(n2550), .Y(n2405) );
  MUX2X1 U2168 ( .B(n1574), .A(n1575), .S(n2557), .Y(n1573) );
  INVX4 U2169 ( .A(n475), .Y(n2557) );
  INVX1 U2170 ( .A(\addr<13> ), .Y(n463) );
  INVX1 U2171 ( .A(n463), .Y(n464) );
  INVX1 U2172 ( .A(n4003), .Y(n465) );
  MUX2X1 U2173 ( .B(n2466), .A(n2465), .S(n1447), .Y(n2464) );
  INVX2 U2174 ( .A(n479), .Y(n466) );
  MUX2X1 U2175 ( .B(n1560), .A(n1559), .S(n475), .Y(n1558) );
  INVX1 U2176 ( .A(n4552), .Y(n467) );
  MUX2X1 U2177 ( .B(n1735), .A(n1736), .S(n2554), .Y(n1734) );
  INVX1 U2178 ( .A(n1507), .Y(n468) );
  INVX1 U2179 ( .A(n468), .Y(n469) );
  INVX1 U2180 ( .A(n468), .Y(n470) );
  INVX1 U2181 ( .A(n105), .Y(n471) );
  INVX1 U2182 ( .A(n471), .Y(n472) );
  INVX1 U2183 ( .A(n2696), .Y(n473) );
  INVX1 U2184 ( .A(n502), .Y(n474) );
  INVX1 U2185 ( .A(n1302), .Y(n476) );
  INVX1 U2186 ( .A(n2633), .Y(n477) );
  INVX1 U2187 ( .A(n2633), .Y(n2632) );
  MUX2X1 U2188 ( .B(n2475), .A(n2474), .S(n478), .Y(n2473) );
  INVX1 U2189 ( .A(n2588), .Y(n479) );
  INVX1 U2190 ( .A(n479), .Y(n480) );
  INVX1 U2191 ( .A(n1511), .Y(n481) );
  MUX2X1 U2192 ( .B(n1531), .A(n1532), .S(n2557), .Y(n1530) );
  INVX1 U2193 ( .A(n1290), .Y(n482) );
  INVX1 U2194 ( .A(n3597), .Y(n483) );
  AND2X2 U2195 ( .A(n2634), .B(n564), .Y(n484) );
  AND2X2 U2196 ( .A(n560), .B(n1488), .Y(n485) );
  MUX2X1 U2197 ( .B(\mem<45><0> ), .A(\mem<44><0> ), .S(n459), .Y(n1540) );
  MUX2X1 U2198 ( .B(\mem<13><1> ), .A(\mem<12><1> ), .S(n493), .Y(n1640) );
  MUX2X1 U2199 ( .B(n1582), .A(n1576), .S(n2548), .Y(n1586) );
  INVX1 U2200 ( .A(n532), .Y(n486) );
  INVX1 U2201 ( .A(n2586), .Y(n487) );
  INVX1 U2202 ( .A(n487), .Y(n488) );
  INVX1 U2203 ( .A(n2583), .Y(n489) );
  MUX2X1 U2204 ( .B(\mem<25><0> ), .A(\mem<24><0> ), .S(n1471), .Y(n1559) );
  AND2X2 U2205 ( .A(n60), .B(n2962), .Y(n490) );
  INVX1 U2206 ( .A(n2588), .Y(n491) );
  INVX1 U2207 ( .A(n2583), .Y(n492) );
  MUX2X1 U2208 ( .B(n2403), .A(n2404), .S(n2561), .Y(n2402) );
  INVX2 U2209 ( .A(n2596), .Y(n4552) );
  MUX2X1 U2210 ( .B(\mem<47><5> ), .A(\mem<46><5> ), .S(n560), .Y(n2372) );
  INVX1 U2211 ( .A(n378), .Y(n4203) );
  MUX2X1 U2212 ( .B(n1565), .A(n1566), .S(n510), .Y(n1564) );
  INVX1 U2213 ( .A(n559), .Y(n494) );
  INVX1 U2214 ( .A(n2609), .Y(n495) );
  INVX1 U2215 ( .A(n495), .Y(n496) );
  MUX2X1 U2216 ( .B(n2357), .A(n2356), .S(n2549), .Y(n2355) );
  INVX2 U2217 ( .A(n2565), .Y(n2571) );
  INVX1 U2218 ( .A(n2555), .Y(n546) );
  INVX1 U2219 ( .A(n2569), .Y(n497) );
  INVX1 U2220 ( .A(N182), .Y(n2718) );
  MUX2X1 U2221 ( .B(\mem<31><3> ), .A(\mem<30><3> ), .S(n498), .Y(n1751) );
  INVX1 U2222 ( .A(n1444), .Y(n1435) );
  MUX2X1 U2223 ( .B(n1595), .A(n1594), .S(n523), .Y(n1593) );
  INVX1 U2224 ( .A(n2569), .Y(n498) );
  MUX2X1 U2225 ( .B(n2408), .A(n2405), .S(n2547), .Y(n2412) );
  NAND2X1 U2226 ( .A(\mem<40><5> ), .B(n497), .Y(n499) );
  NAND2X1 U2227 ( .A(\mem<41><5> ), .B(n2574), .Y(n500) );
  AND2X2 U2228 ( .A(n538), .B(n2612), .Y(n501) );
  MUX2X1 U2229 ( .B(\mem<9><5> ), .A(\mem<8><5> ), .S(n497), .Y(n2403) );
  INVX1 U2230 ( .A(n1484), .Y(n502) );
  INVX1 U2231 ( .A(n503), .Y(n504) );
  INVX1 U2232 ( .A(n4551), .Y(n505) );
  MUX2X1 U2233 ( .B(n1608), .A(n1607), .S(n523), .Y(n1606) );
  INVX4 U2234 ( .A(n534), .Y(n523) );
  MUX2X1 U2235 ( .B(n2374), .A(n96), .S(n2549), .Y(n2373) );
  INVX1 U2236 ( .A(n3268), .Y(n506) );
  INVX1 U2237 ( .A(n2567), .Y(n507) );
  INVX1 U2238 ( .A(n2605), .Y(n2566) );
  INVX8 U2239 ( .A(n2605), .Y(n547) );
  INVX1 U2240 ( .A(n2614), .Y(n508) );
  INVX1 U2241 ( .A(n508), .Y(n509) );
  AND2X2 U2242 ( .A(n2636), .B(n528), .Y(n2707) );
  INVX1 U2243 ( .A(n515), .Y(n510) );
  INVX1 U2244 ( .A(n3140), .Y(n1296) );
  MUX2X1 U2245 ( .B(n2372), .A(n2371), .S(n2549), .Y(n2370) );
  MUX2X1 U2246 ( .B(n2369), .A(n2368), .S(n448), .Y(n2367) );
  MUX2X1 U2247 ( .B(n1562), .A(n1563), .S(n2561), .Y(n1561) );
  AND2X2 U2248 ( .A(n576), .B(n2635), .Y(n511) );
  INVX1 U2249 ( .A(n517), .Y(n512) );
  INVX1 U2250 ( .A(n534), .Y(n517) );
  MUX2X1 U2251 ( .B(n1748), .A(n1747), .S(n478), .Y(n1746) );
  MUX2X1 U2252 ( .B(n1725), .A(n1728), .S(n513), .Y(n1732) );
  INVX1 U2253 ( .A(n534), .Y(n515) );
  INVX1 U2254 ( .A(n3242), .Y(n514) );
  INVX4 U2255 ( .A(n1465), .Y(n1452) );
  MUX2X1 U2256 ( .B(n1623), .A(n1622), .S(n515), .Y(n1621) );
  MUX2X1 U2257 ( .B(\mem<61><1> ), .A(\mem<60><1> ), .S(n516), .Y(n1591) );
  INVX1 U2258 ( .A(n559), .Y(n516) );
  INVX2 U2259 ( .A(n2566), .Y(n2567) );
  MUX2X1 U2260 ( .B(\mem<27><0> ), .A(\mem<26><0> ), .S(n462), .Y(n1560) );
  MUX2X1 U2261 ( .B(n1650), .A(n1649), .S(n517), .Y(n1648) );
  INVX1 U2262 ( .A(n367), .Y(n518) );
  MUX2X1 U2263 ( .B(n1645), .A(n1648), .S(n519), .Y(n1652) );
  AND2X2 U2264 ( .A(n558), .B(n355), .Y(n520) );
  AND2X2 U2265 ( .A(n2612), .B(n356), .Y(n521) );
  MUX2X1 U2266 ( .B(\mem<57><0> ), .A(\mem<56><0> ), .S(n462), .Y(n1528) );
  INVX1 U2267 ( .A(\addr<14> ), .Y(n2655) );
  MUX2X1 U2268 ( .B(\mem<49><0> ), .A(\mem<48><0> ), .S(n1471), .Y(n1534) );
  INVX1 U2269 ( .A(n479), .Y(n522) );
  MUX2X1 U2270 ( .B(n1535), .A(n1534), .S(n523), .Y(n1533) );
  MUX2X1 U2271 ( .B(\mem<37><0> ), .A(\mem<36><0> ), .S(n1471), .Y(n1546) );
  INVX1 U2272 ( .A(n2557), .Y(n1447) );
  INVX1 U2273 ( .A(n2557), .Y(n1462) );
  MUX2X1 U2274 ( .B(n1809), .A(n1810), .S(n2542), .Y(n1808) );
  INVX1 U2275 ( .A(n382), .Y(n524) );
  INVX1 U2276 ( .A(n2652), .Y(n525) );
  INVX1 U2277 ( .A(n381), .Y(n3320) );
  BUFX2 U2278 ( .A(n442), .Y(n2626) );
  INVX1 U2279 ( .A(\addr<13> ), .Y(n2675) );
  MUX2X1 U2280 ( .B(\mem<11><5> ), .A(\mem<10><5> ), .S(n560), .Y(n2404) );
  MUX2X1 U2281 ( .B(\mem<47><0> ), .A(\mem<46><0> ), .S(n449), .Y(n1541) );
  INVX1 U2282 ( .A(n81), .Y(n526) );
  INVX1 U2283 ( .A(n2603), .Y(n527) );
  INVX1 U2284 ( .A(N181), .Y(n528) );
  INVX1 U2285 ( .A(n26), .Y(n529) );
  INVX1 U2286 ( .A(n443), .Y(n3065) );
  MUX2X1 U2287 ( .B(n1651), .A(n1636), .S(n2541), .Y(n1654) );
  MUX2X1 U2288 ( .B(n1732), .A(n1733), .S(n2543), .Y(n1731) );
  INVX1 U2289 ( .A(n46), .Y(n530) );
  INVX1 U2290 ( .A(n49), .Y(n531) );
  INVX1 U2291 ( .A(n1514), .Y(n532) );
  INVX1 U2292 ( .A(n532), .Y(n533) );
  MUX2X1 U2293 ( .B(n1605), .A(n1603), .S(n448), .Y(n1602) );
  INVX4 U2294 ( .A(n448), .Y(n2544) );
  MUX2X1 U2295 ( .B(n1544), .A(n1543), .S(n2551), .Y(n1542) );
  INVX2 U2296 ( .A(n2551), .Y(n2553) );
  INVX1 U2297 ( .A(n481), .Y(n535) );
  INVX1 U2298 ( .A(n571), .Y(n574) );
  BUFX2 U2299 ( .A(n395), .Y(n2627) );
  AND2X2 U2300 ( .A(n1296), .B(n536), .Y(n2784) );
  AND2X2 U2301 ( .A(n480), .B(n484), .Y(n537) );
  AND2X2 U2302 ( .A(n480), .B(n484), .Y(n538) );
  INVX1 U2303 ( .A(n1518), .Y(n539) );
  INVX1 U2304 ( .A(n1302), .Y(n3772) );
  AND2X2 U2305 ( .A(n388), .B(n1454), .Y(n540) );
  MUX2X1 U2306 ( .B(n1814), .A(n1811), .S(n2547), .Y(n2337) );
  INVX1 U2307 ( .A(n2614), .Y(n541) );
  MUX2X1 U2308 ( .B(\mem<35><5> ), .A(\mem<34><5> ), .S(n516), .Y(n2380) );
  INVX1 U2309 ( .A(n3927), .Y(n542) );
  INVX2 U2310 ( .A(n397), .Y(n3927) );
  AND2X2 U2311 ( .A(n2594), .B(n485), .Y(n544) );
  AND2X2 U2312 ( .A(n2635), .B(n477), .Y(n545) );
  INVX1 U2313 ( .A(n93), .Y(n2584) );
  MUX2X1 U2314 ( .B(n1553), .A(n1554), .S(n2543), .Y(n1551) );
  MUX2X1 U2315 ( .B(n1766), .A(n1765), .S(n546), .Y(n1764) );
  NOR2X1 U2316 ( .A(\addr<10> ), .B(\addr<9> ), .Y(n548) );
  AND2X2 U2317 ( .A(n1296), .B(\mem<58><6> ), .Y(n2826) );
  INVX1 U2318 ( .A(n1483), .Y(n549) );
  INVX1 U2319 ( .A(n1483), .Y(n550) );
  INVX1 U2320 ( .A(n70), .Y(n551) );
  INVX1 U2321 ( .A(n567), .Y(n552) );
  INVX1 U2322 ( .A(n552), .Y(n553) );
  INVX1 U2323 ( .A(n373), .Y(n2612) );
  MUX2X1 U2324 ( .B(n2338), .A(n2341), .S(n452), .Y(n2352) );
  MUX2X1 U2325 ( .B(n1793), .A(n1808), .S(n554), .Y(n2354) );
  MUX2X1 U2326 ( .B(n557), .A(n556), .S(n2565), .Y(n555) );
  AND2X2 U2327 ( .A(n392), .B(n581), .Y(n558) );
  INVX2 U2328 ( .A(n1464), .Y(n559) );
  INVX8 U2329 ( .A(n559), .Y(n560) );
  INVX2 U2330 ( .A(n396), .Y(n2964) );
  NOR2X1 U2331 ( .A(n1465), .B(n97), .Y(n2699) );
  AND2X2 U2332 ( .A(\mem<18><5> ), .B(n1514), .Y(n562) );
  AND2X2 U2333 ( .A(\mem<20><5> ), .B(n1484), .Y(n563) );
  NOR2X1 U2334 ( .A(\addr<15> ), .B(\addr<14> ), .Y(n565) );
  INVX2 U2335 ( .A(n2621), .Y(n4551) );
  MUX2X1 U2336 ( .B(\mem<29><0> ), .A(\mem<28><0> ), .S(n1465), .Y(n1556) );
  INVX1 U2337 ( .A(n4128), .Y(n566) );
  AND2X2 U2338 ( .A(n2722), .B(n3), .Y(n567) );
  INVX1 U2339 ( .A(n93), .Y(n3091) );
  AND2X2 U2340 ( .A(N182), .B(n15), .Y(n2669) );
  MUX2X1 U2341 ( .B(n1581), .A(n1580), .S(n2551), .Y(n1576) );
  INVX1 U2342 ( .A(n1467), .Y(n3268) );
  MUX2X1 U2343 ( .B(n1556), .A(n1557), .S(n9), .Y(n1555) );
  INVX4 U2344 ( .A(n2634), .Y(n2545) );
  AND2X2 U2345 ( .A(n560), .B(n1488), .Y(n568) );
  AND2X2 U2346 ( .A(n560), .B(n1488), .Y(n569) );
  INVX1 U2347 ( .A(n1448), .Y(n2377) );
  AND2X2 U2348 ( .A(n1454), .B(n389), .Y(n570) );
  INVX4 U2349 ( .A(n52), .Y(n2962) );
  INVX1 U2350 ( .A(n1511), .Y(n571) );
  INVX1 U2351 ( .A(n481), .Y(n572) );
  INVX1 U2352 ( .A(n481), .Y(n573) );
  INVX1 U2353 ( .A(n107), .Y(n575) );
  INVX1 U2354 ( .A(n2632), .Y(n576) );
  INVX1 U2355 ( .A(n2634), .Y(n577) );
  INVX1 U2356 ( .A(n492), .Y(n578) );
  NOR2X1 U2357 ( .A(n576), .B(n577), .Y(n580) );
  INVX1 U2358 ( .A(n580), .Y(n579) );
  INVX1 U2359 ( .A(n582), .Y(n581) );
  INVX1 U2360 ( .A(n374), .Y(n582) );
  INVX1 U2361 ( .A(n374), .Y(n583) );
  INVX1 U2362 ( .A(rst), .Y(n2637) );
  AND2X2 U2363 ( .A(n511), .B(n489), .Y(n584) );
  OR2X1 U2364 ( .A(n2915), .B(n2914), .Y(n585) );
  INVX1 U2365 ( .A(n585), .Y(n586) );
  OR2X1 U2366 ( .A(n2919), .B(n2918), .Y(n587) );
  INVX1 U2367 ( .A(n587), .Y(n588) );
  OR2X1 U2368 ( .A(n2923), .B(n2922), .Y(n589) );
  INVX1 U2369 ( .A(n589), .Y(n590) );
  OR2X1 U2370 ( .A(n2927), .B(n2926), .Y(n591) );
  INVX1 U2371 ( .A(n591), .Y(n592) );
  OR2X1 U2372 ( .A(n2931), .B(n2930), .Y(n593) );
  INVX1 U2373 ( .A(n593), .Y(n594) );
  OR2X1 U2374 ( .A(n2935), .B(n2934), .Y(n595) );
  INVX1 U2375 ( .A(n595), .Y(n596) );
  OR2X1 U2376 ( .A(n2939), .B(n2938), .Y(n597) );
  INVX1 U2377 ( .A(n597), .Y(n598) );
  OR2X1 U2378 ( .A(n2943), .B(n2942), .Y(n600) );
  INVX1 U2379 ( .A(n600), .Y(n601) );
  OR2X1 U2380 ( .A(n2947), .B(n2946), .Y(n609) );
  INVX1 U2381 ( .A(n609), .Y(n610) );
  OR2X1 U2382 ( .A(n2951), .B(n2950), .Y(n611) );
  INVX1 U2383 ( .A(n611), .Y(n612) );
  OR2X1 U2384 ( .A(n2955), .B(n2954), .Y(n613) );
  INVX1 U2385 ( .A(n613), .Y(n614) );
  OR2X1 U2386 ( .A(n2959), .B(n2958), .Y(n615) );
  INVX1 U2387 ( .A(n615), .Y(n616) );
  OR2X1 U2388 ( .A(n2966), .B(n2965), .Y(n617) );
  INVX1 U2389 ( .A(n617), .Y(n618) );
  OR2X1 U2390 ( .A(n2970), .B(n2969), .Y(n619) );
  INVX1 U2391 ( .A(n619), .Y(n620) );
  OR2X1 U2392 ( .A(n2974), .B(n2973), .Y(n621) );
  INVX1 U2393 ( .A(n621), .Y(n622) );
  OR2X1 U2394 ( .A(n2978), .B(n2977), .Y(n623) );
  INVX1 U2395 ( .A(n623), .Y(n624) );
  OR2X1 U2396 ( .A(n2982), .B(n2981), .Y(n626) );
  INVX1 U2397 ( .A(n626), .Y(n627) );
  OR2X1 U2398 ( .A(n2986), .B(n2985), .Y(n628) );
  INVX1 U2399 ( .A(n628), .Y(n629) );
  OR2X1 U2400 ( .A(n2990), .B(n2989), .Y(n630) );
  INVX1 U2401 ( .A(n630), .Y(n631) );
  OR2X1 U2402 ( .A(n2994), .B(n2993), .Y(n632) );
  INVX1 U2403 ( .A(n632), .Y(n633) );
  OR2X1 U2404 ( .A(n2998), .B(n2997), .Y(n634) );
  INVX1 U2405 ( .A(n634), .Y(n635) );
  OR2X1 U2406 ( .A(n3002), .B(n3001), .Y(n636) );
  INVX1 U2407 ( .A(n636), .Y(n637) );
  OR2X1 U2408 ( .A(n3006), .B(n3005), .Y(n638) );
  INVX1 U2409 ( .A(n638), .Y(n639) );
  OR2X1 U2410 ( .A(n3010), .B(n3009), .Y(n640) );
  INVX1 U2411 ( .A(n640), .Y(n641) );
  OR2X1 U2412 ( .A(n2917), .B(n2916), .Y(n642) );
  INVX1 U2413 ( .A(n642), .Y(n643) );
  OR2X1 U2414 ( .A(n2921), .B(n2920), .Y(n644) );
  INVX1 U2415 ( .A(n644), .Y(n645) );
  OR2X1 U2416 ( .A(n2925), .B(n2924), .Y(n646) );
  INVX1 U2417 ( .A(n646), .Y(n647) );
  OR2X1 U2418 ( .A(n2929), .B(n2928), .Y(n648) );
  INVX1 U2419 ( .A(n648), .Y(n649) );
  OR2X1 U2420 ( .A(n2933), .B(n2932), .Y(n650) );
  INVX1 U2421 ( .A(n650), .Y(n651) );
  OR2X1 U2422 ( .A(n2937), .B(n2936), .Y(n652) );
  INVX1 U2423 ( .A(n652), .Y(n653) );
  OR2X1 U2424 ( .A(n2941), .B(n2940), .Y(n654) );
  INVX1 U2425 ( .A(n654), .Y(n655) );
  OR2X1 U2426 ( .A(n2945), .B(n2944), .Y(n656) );
  INVX1 U2427 ( .A(n656), .Y(n657) );
  OR2X1 U2428 ( .A(n2949), .B(n2948), .Y(n658) );
  INVX1 U2429 ( .A(n658), .Y(n659) );
  OR2X1 U2430 ( .A(n2953), .B(n2952), .Y(n660) );
  INVX1 U2431 ( .A(n660), .Y(n661) );
  OR2X1 U2432 ( .A(n2957), .B(n2956), .Y(n662) );
  INVX1 U2433 ( .A(n662), .Y(n663) );
  OR2X1 U2434 ( .A(n2961), .B(n2960), .Y(n664) );
  INVX1 U2435 ( .A(n664), .Y(n665) );
  OR2X1 U2436 ( .A(n2968), .B(n2967), .Y(n666) );
  INVX1 U2437 ( .A(n666), .Y(n667) );
  OR2X1 U2438 ( .A(n2972), .B(n2971), .Y(n668) );
  INVX1 U2439 ( .A(n668), .Y(n669) );
  OR2X1 U2440 ( .A(n2976), .B(n2975), .Y(n670) );
  INVX1 U2441 ( .A(n670), .Y(n671) );
  OR2X1 U2442 ( .A(n2980), .B(n2979), .Y(n672) );
  INVX1 U2443 ( .A(n672), .Y(n673) );
  OR2X1 U2444 ( .A(n2984), .B(n2983), .Y(n674) );
  INVX1 U2445 ( .A(n674), .Y(n675) );
  OR2X1 U2446 ( .A(n2988), .B(n2987), .Y(n676) );
  INVX1 U2447 ( .A(n676), .Y(n677) );
  OR2X1 U2448 ( .A(n2992), .B(n2991), .Y(n678) );
  INVX1 U2449 ( .A(n678), .Y(n679) );
  OR2X1 U2450 ( .A(n2996), .B(n2995), .Y(n680) );
  INVX1 U2451 ( .A(n680), .Y(n681) );
  OR2X1 U2452 ( .A(n3000), .B(n2999), .Y(n682) );
  INVX1 U2453 ( .A(n682), .Y(n683) );
  OR2X1 U2454 ( .A(n3004), .B(n3003), .Y(n684) );
  INVX1 U2455 ( .A(n684), .Y(n685) );
  OR2X1 U2456 ( .A(n3008), .B(n3007), .Y(n686) );
  INVX1 U2457 ( .A(n686), .Y(n687) );
  OR2X1 U2458 ( .A(n3012), .B(n3011), .Y(n688) );
  INVX1 U2459 ( .A(n688), .Y(n689) );
  AND2X2 U2460 ( .A(n2625), .B(n1500), .Y(n690) );
  INVX1 U2461 ( .A(n690), .Y(n691) );
  AND2X2 U2462 ( .A(n2625), .B(n2599), .Y(n692) );
  INVX1 U2463 ( .A(n692), .Y(n693) );
  AND2X2 U2464 ( .A(n2626), .B(n2599), .Y(n694) );
  INVX1 U2465 ( .A(n694), .Y(n695) );
  AND2X2 U2466 ( .A(n2626), .B(n2585), .Y(n696) );
  INVX1 U2467 ( .A(n696), .Y(n697) );
  AND2X2 U2468 ( .A(n2624), .B(n2585), .Y(n698) );
  INVX1 U2469 ( .A(n698), .Y(n699) );
  INVX1 U2470 ( .A(n700), .Y(n701) );
  INVX1 U2471 ( .A(n702), .Y(n703) );
  AND2X1 U2472 ( .A(n3242), .B(n1478), .Y(n704) );
  INVX1 U2473 ( .A(n704), .Y(n705) );
  AND2X1 U2474 ( .A(n3242), .B(n1290), .Y(n706) );
  INVX1 U2475 ( .A(n706), .Y(n707) );
  AND2X1 U2476 ( .A(n1289), .B(n3398), .Y(n708) );
  INVX1 U2477 ( .A(n708), .Y(n709) );
  AND2X1 U2478 ( .A(n3398), .B(n3423), .Y(n710) );
  INVX1 U2479 ( .A(n710), .Y(n711) );
  AND2X1 U2480 ( .A(n3448), .B(n3423), .Y(n712) );
  INVX1 U2481 ( .A(n712), .Y(n713) );
  AND2X1 U2482 ( .A(n3448), .B(n3473), .Y(n714) );
  INVX1 U2483 ( .A(n714), .Y(n715) );
  AND2X1 U2484 ( .A(n411), .B(n3473), .Y(n716) );
  INVX1 U2485 ( .A(n716), .Y(n717) );
  AND2X1 U2486 ( .A(n411), .B(n3522), .Y(n718) );
  INVX1 U2487 ( .A(n718), .Y(n719) );
  AND2X1 U2488 ( .A(n3547), .B(n3522), .Y(n720) );
  INVX1 U2489 ( .A(n720), .Y(n721) );
  AND2X1 U2490 ( .A(n3547), .B(n3572), .Y(n722) );
  INVX1 U2491 ( .A(n722), .Y(n723) );
  AND2X1 U2492 ( .A(n3572), .B(n3597), .Y(n724) );
  INVX1 U2493 ( .A(n724), .Y(n725) );
  AND2X1 U2494 ( .A(n3597), .B(n1277), .Y(n726) );
  INVX1 U2495 ( .A(n726), .Y(n727) );
  AND2X1 U2496 ( .A(n3646), .B(n1277), .Y(n728) );
  INVX1 U2497 ( .A(n728), .Y(n729) );
  AND2X1 U2498 ( .A(n3646), .B(n3671), .Y(n730) );
  INVX1 U2499 ( .A(n730), .Y(n731) );
  AND2X1 U2500 ( .A(n3696), .B(n3671), .Y(n732) );
  INVX1 U2501 ( .A(n732), .Y(n733) );
  AND2X1 U2502 ( .A(n3696), .B(n3721), .Y(n734) );
  INVX1 U2503 ( .A(n734), .Y(n735) );
  AND2X1 U2504 ( .A(n3746), .B(n3721), .Y(n736) );
  INVX1 U2505 ( .A(n736), .Y(n737) );
  AND2X1 U2506 ( .A(n3746), .B(n1288), .Y(n738) );
  INVX1 U2507 ( .A(n738), .Y(n739) );
  AND2X1 U2508 ( .A(n1288), .B(n1518), .Y(n740) );
  INVX1 U2509 ( .A(n740), .Y(n741) );
  AND2X1 U2510 ( .A(n1518), .B(n1287), .Y(n742) );
  INVX1 U2511 ( .A(n742), .Y(n743) );
  AND2X1 U2512 ( .A(n2601), .B(n1287), .Y(n744) );
  INVX1 U2513 ( .A(n744), .Y(n745) );
  AND2X1 U2514 ( .A(n2601), .B(n1453), .Y(n746) );
  INVX1 U2515 ( .A(n746), .Y(n747) );
  AND2X1 U2516 ( .A(n1480), .B(n1453), .Y(n748) );
  INVX1 U2517 ( .A(n748), .Y(n749) );
  AND2X2 U2518 ( .A(n1480), .B(n550), .Y(n750) );
  INVX1 U2519 ( .A(n750), .Y(n751) );
  AND2X2 U2520 ( .A(n2591), .B(n549), .Y(n752) );
  INVX1 U2521 ( .A(n752), .Y(n753) );
  AND2X1 U2522 ( .A(n2591), .B(n1485), .Y(n754) );
  INVX1 U2523 ( .A(n754), .Y(n755) );
  AND2X1 U2524 ( .A(n4003), .B(n1485), .Y(n756) );
  INVX1 U2525 ( .A(n756), .Y(n757) );
  AND2X1 U2526 ( .A(n4028), .B(n4003), .Y(n758) );
  INVX1 U2527 ( .A(n758), .Y(n759) );
  AND2X1 U2528 ( .A(n4053), .B(n4028), .Y(n760) );
  INVX1 U2529 ( .A(n760), .Y(n761) );
  AND2X1 U2530 ( .A(n4053), .B(n4078), .Y(n762) );
  INVX1 U2531 ( .A(n762), .Y(n763) );
  AND2X1 U2532 ( .A(n4103), .B(n4078), .Y(n764) );
  INVX1 U2533 ( .A(n764), .Y(n765) );
  AND2X1 U2534 ( .A(n4103), .B(n4128), .Y(n766) );
  INVX1 U2535 ( .A(n766), .Y(n767) );
  AND2X1 U2536 ( .A(n4153), .B(n4128), .Y(n768) );
  INVX1 U2537 ( .A(n768), .Y(n769) );
  AND2X1 U2538 ( .A(n4153), .B(n1292), .Y(n770) );
  INVX1 U2539 ( .A(n770), .Y(n771) );
  AND2X1 U2540 ( .A(n4202), .B(n1292), .Y(n772) );
  INVX1 U2541 ( .A(n772), .Y(n773) );
  AND2X1 U2542 ( .A(n1456), .B(n4202), .Y(n774) );
  INVX1 U2543 ( .A(n774), .Y(n775) );
  AND2X1 U2544 ( .A(n4252), .B(n1456), .Y(n776) );
  INVX1 U2545 ( .A(n776), .Y(n777) );
  AND2X1 U2546 ( .A(n4252), .B(n4277), .Y(n778) );
  INVX1 U2547 ( .A(n778), .Y(n779) );
  AND2X1 U2548 ( .A(n4302), .B(n4277), .Y(n780) );
  INVX1 U2549 ( .A(n780), .Y(n781) );
  AND2X1 U2550 ( .A(n4302), .B(n4327), .Y(n782) );
  INVX1 U2551 ( .A(n782), .Y(n783) );
  AND2X1 U2552 ( .A(n4352), .B(n4327), .Y(n784) );
  INVX1 U2553 ( .A(n784), .Y(n785) );
  AND2X1 U2554 ( .A(n4352), .B(n4377), .Y(n786) );
  INVX1 U2555 ( .A(n786), .Y(n787) );
  AND2X1 U2556 ( .A(n4377), .B(n4402), .Y(n788) );
  INVX1 U2557 ( .A(n788), .Y(n789) );
  AND2X1 U2558 ( .A(n1291), .B(n4402), .Y(n790) );
  INVX1 U2559 ( .A(n790), .Y(n791) );
  AND2X2 U2560 ( .A(n4451), .B(n1291), .Y(n792) );
  INVX1 U2561 ( .A(n792), .Y(n793) );
  AND2X2 U2562 ( .A(n4451), .B(n4476), .Y(n794) );
  INVX1 U2563 ( .A(n794), .Y(n795) );
  AND2X2 U2564 ( .A(n46), .B(n4476), .Y(n796) );
  INVX1 U2565 ( .A(n796), .Y(n797) );
  AND2X2 U2566 ( .A(n46), .B(n4526), .Y(n798) );
  INVX1 U2567 ( .A(n798), .Y(n799) );
  AND2X2 U2568 ( .A(n4551), .B(n4526), .Y(n800) );
  INVX1 U2569 ( .A(n800), .Y(n801) );
  BUFX2 U2570 ( .A(n608), .Y(n802) );
  BUFX2 U2571 ( .A(n607), .Y(n803) );
  BUFX2 U2572 ( .A(n606), .Y(n804) );
  BUFX2 U2573 ( .A(n605), .Y(n805) );
  BUFX2 U2574 ( .A(n604), .Y(n806) );
  BUFX2 U2575 ( .A(n603), .Y(n807) );
  BUFX2 U2576 ( .A(n602), .Y(n808) );
  BUFX2 U2577 ( .A(n599), .Y(n809) );
  BUFX2 U2578 ( .A(n4554), .Y(n810) );
  BUFX2 U2579 ( .A(n4557), .Y(n811) );
  BUFX2 U2580 ( .A(n4560), .Y(n812) );
  BUFX2 U2581 ( .A(n4563), .Y(n813) );
  BUFX2 U2582 ( .A(n4566), .Y(n814) );
  BUFX2 U2583 ( .A(n4569), .Y(n815) );
  BUFX2 U2584 ( .A(n4572), .Y(n816) );
  BUFX2 U2585 ( .A(n4576), .Y(n817) );
  AND2X2 U2586 ( .A(\mem<5><0> ), .B(n357), .Y(n818) );
  INVX1 U2587 ( .A(n818), .Y(n819) );
  AND2X2 U2588 ( .A(\mem<7><0> ), .B(n383), .Y(n820) );
  INVX1 U2589 ( .A(n820), .Y(n821) );
  AND2X2 U2590 ( .A(\mem<3><0> ), .B(n572), .Y(n822) );
  INVX1 U2591 ( .A(n822), .Y(n823) );
  AND2X2 U2592 ( .A(\mem<5><1> ), .B(n357), .Y(n824) );
  INVX1 U2593 ( .A(n824), .Y(n825) );
  AND2X2 U2594 ( .A(\mem<7><1> ), .B(n383), .Y(n826) );
  INVX1 U2595 ( .A(n826), .Y(n827) );
  AND2X2 U2596 ( .A(\mem<3><1> ), .B(n573), .Y(n828) );
  INVX1 U2597 ( .A(n828), .Y(n829) );
  AND2X2 U2598 ( .A(\mem<5><7> ), .B(n357), .Y(n830) );
  INVX1 U2599 ( .A(n830), .Y(n831) );
  AND2X2 U2600 ( .A(\mem<7><7> ), .B(n383), .Y(n832) );
  INVX1 U2601 ( .A(n832), .Y(n833) );
  AND2X2 U2602 ( .A(\mem<3><7> ), .B(n535), .Y(n834) );
  INVX1 U2603 ( .A(n834), .Y(n835) );
  AND2X2 U2604 ( .A(\mem<13><2> ), .B(n1436), .Y(n836) );
  INVX1 U2605 ( .A(n836), .Y(n837) );
  AND2X2 U2606 ( .A(\mem<15><2> ), .B(n1442), .Y(n838) );
  INVX1 U2607 ( .A(n838), .Y(n839) );
  AND2X2 U2608 ( .A(\mem<9><2> ), .B(n1457), .Y(n840) );
  INVX1 U2609 ( .A(n840), .Y(n841) );
  AND2X2 U2610 ( .A(\mem<11><2> ), .B(n1489), .Y(n842) );
  INVX1 U2611 ( .A(n842), .Y(n843) );
  AND2X2 U2612 ( .A(\mem<5><2> ), .B(n434), .Y(n844) );
  INVX1 U2613 ( .A(n844), .Y(n845) );
  AND2X2 U2614 ( .A(\mem<7><2> ), .B(n456), .Y(n846) );
  INVX1 U2615 ( .A(n846), .Y(n847) );
  AND2X2 U2616 ( .A(\mem<0><2> ), .B(n526), .Y(n848) );
  INVX1 U2617 ( .A(n848), .Y(n849) );
  AND2X2 U2618 ( .A(\mem<3><2> ), .B(n573), .Y(n850) );
  INVX1 U2619 ( .A(n850), .Y(n851) );
  AND2X2 U2620 ( .A(\mem<61><2> ), .B(n428), .Y(n852) );
  INVX1 U2621 ( .A(n852), .Y(n853) );
  AND2X2 U2622 ( .A(\mem<63><2> ), .B(n2964), .Y(n854) );
  INVX1 U2623 ( .A(n854), .Y(n855) );
  AND2X2 U2624 ( .A(\mem<56><2> ), .B(n1487), .Y(n856) );
  INVX1 U2625 ( .A(n856), .Y(n857) );
  AND2X2 U2626 ( .A(\mem<59><2> ), .B(n2602), .Y(n858) );
  INVX1 U2627 ( .A(n858), .Y(n859) );
  AND2X2 U2628 ( .A(\mem<53><2> ), .B(n482), .Y(n860) );
  INVX1 U2629 ( .A(n860), .Y(n861) );
  AND2X2 U2630 ( .A(\mem<55><2> ), .B(n1477), .Y(n862) );
  INVX1 U2631 ( .A(n862), .Y(n863) );
  AND2X2 U2632 ( .A(\mem<49><2> ), .B(n440), .Y(n864) );
  INVX1 U2633 ( .A(n864), .Y(n865) );
  AND2X2 U2634 ( .A(\mem<51><2> ), .B(n1491), .Y(n866) );
  INVX1 U2635 ( .A(n866), .Y(n867) );
  AND2X2 U2636 ( .A(\mem<13><3> ), .B(n1436), .Y(n868) );
  INVX1 U2637 ( .A(n868), .Y(n869) );
  AND2X2 U2638 ( .A(\mem<15><3> ), .B(n1442), .Y(n870) );
  INVX1 U2639 ( .A(n870), .Y(n871) );
  AND2X2 U2640 ( .A(\mem<9><3> ), .B(n1457), .Y(n872) );
  INVX1 U2641 ( .A(n872), .Y(n873) );
  AND2X2 U2642 ( .A(\mem<11><3> ), .B(n1489), .Y(n874) );
  INVX1 U2643 ( .A(n874), .Y(n875) );
  AND2X2 U2644 ( .A(\mem<5><3> ), .B(n434), .Y(n876) );
  INVX1 U2645 ( .A(n876), .Y(n877) );
  AND2X2 U2646 ( .A(\mem<7><3> ), .B(n456), .Y(n878) );
  INVX1 U2647 ( .A(n878), .Y(n879) );
  AND2X2 U2648 ( .A(\mem<0><3> ), .B(n526), .Y(n880) );
  INVX1 U2649 ( .A(n880), .Y(n881) );
  AND2X2 U2650 ( .A(\mem<3><3> ), .B(n573), .Y(n882) );
  INVX1 U2651 ( .A(n882), .Y(n883) );
  AND2X2 U2652 ( .A(\mem<61><3> ), .B(n428), .Y(n884) );
  INVX1 U2653 ( .A(n884), .Y(n885) );
  AND2X2 U2654 ( .A(\mem<63><3> ), .B(n2964), .Y(n886) );
  INVX1 U2655 ( .A(n886), .Y(n887) );
  AND2X2 U2656 ( .A(\mem<56><3> ), .B(n1487), .Y(n888) );
  INVX1 U2657 ( .A(n888), .Y(n889) );
  AND2X2 U2658 ( .A(\mem<59><3> ), .B(n2602), .Y(n890) );
  INVX1 U2659 ( .A(n890), .Y(n891) );
  AND2X2 U2660 ( .A(\mem<53><3> ), .B(n482), .Y(n892) );
  INVX1 U2661 ( .A(n892), .Y(n893) );
  AND2X2 U2662 ( .A(\mem<55><3> ), .B(n1477), .Y(n894) );
  INVX1 U2663 ( .A(n894), .Y(n895) );
  AND2X2 U2664 ( .A(\mem<49><3> ), .B(n440), .Y(n896) );
  INVX1 U2665 ( .A(n896), .Y(n897) );
  AND2X2 U2666 ( .A(\mem<51><3> ), .B(n1491), .Y(n898) );
  INVX1 U2667 ( .A(n898), .Y(n899) );
  AND2X2 U2668 ( .A(\mem<13><4> ), .B(n1436), .Y(n900) );
  INVX1 U2669 ( .A(n900), .Y(n901) );
  AND2X2 U2670 ( .A(\mem<15><4> ), .B(n1442), .Y(n902) );
  INVX1 U2671 ( .A(n902), .Y(n903) );
  AND2X2 U2672 ( .A(\mem<9><4> ), .B(n1457), .Y(n904) );
  INVX1 U2673 ( .A(n904), .Y(n905) );
  AND2X2 U2674 ( .A(\mem<11><4> ), .B(n1489), .Y(n906) );
  INVX1 U2675 ( .A(n906), .Y(n907) );
  AND2X2 U2676 ( .A(\mem<5><4> ), .B(n434), .Y(n908) );
  INVX1 U2677 ( .A(n908), .Y(n909) );
  AND2X2 U2678 ( .A(\mem<7><4> ), .B(n456), .Y(n910) );
  INVX1 U2679 ( .A(n910), .Y(n911) );
  AND2X2 U2680 ( .A(\mem<0><4> ), .B(n526), .Y(n912) );
  INVX1 U2681 ( .A(n912), .Y(n913) );
  AND2X2 U2682 ( .A(\mem<3><4> ), .B(n573), .Y(n914) );
  INVX1 U2683 ( .A(n914), .Y(n915) );
  AND2X2 U2684 ( .A(\mem<61><4> ), .B(n428), .Y(n916) );
  INVX1 U2685 ( .A(n916), .Y(n917) );
  AND2X2 U2686 ( .A(\mem<63><4> ), .B(n2964), .Y(n918) );
  INVX1 U2687 ( .A(n918), .Y(n919) );
  AND2X2 U2688 ( .A(\mem<56><4> ), .B(n1487), .Y(n920) );
  INVX1 U2689 ( .A(n920), .Y(n921) );
  AND2X2 U2690 ( .A(\mem<59><4> ), .B(n2602), .Y(n922) );
  INVX1 U2691 ( .A(n922), .Y(n923) );
  AND2X2 U2692 ( .A(\mem<53><4> ), .B(n482), .Y(n924) );
  INVX1 U2693 ( .A(n924), .Y(n925) );
  AND2X2 U2694 ( .A(\mem<55><4> ), .B(n1477), .Y(n926) );
  INVX1 U2695 ( .A(n926), .Y(n927) );
  AND2X2 U2696 ( .A(\mem<49><4> ), .B(n440), .Y(n928) );
  INVX1 U2697 ( .A(n928), .Y(n929) );
  AND2X2 U2698 ( .A(\mem<51><4> ), .B(n1491), .Y(n930) );
  INVX1 U2699 ( .A(n930), .Y(n931) );
  AND2X2 U2700 ( .A(\mem<29><2> ), .B(n3849), .Y(n932) );
  INVX1 U2701 ( .A(n932), .Y(n933) );
  AND2X2 U2702 ( .A(\mem<31><2> ), .B(n433), .Y(n934) );
  INVX1 U2703 ( .A(n934), .Y(n935) );
  AND2X2 U2704 ( .A(\mem<24><2> ), .B(n465), .Y(n936) );
  INVX1 U2705 ( .A(n936), .Y(n937) );
  AND2X2 U2706 ( .A(\mem<27><2> ), .B(n3901), .Y(n938) );
  INVX1 U2707 ( .A(n938), .Y(n939) );
  AND2X2 U2708 ( .A(\mem<21><2> ), .B(n79), .Y(n940) );
  INVX1 U2709 ( .A(n940), .Y(n941) );
  AND2X2 U2710 ( .A(\mem<23><2> ), .B(n437), .Y(n942) );
  INVX1 U2711 ( .A(n942), .Y(n943) );
  AND2X2 U2712 ( .A(\mem<17><2> ), .B(n77), .Y(n944) );
  INVX1 U2713 ( .A(n944), .Y(n945) );
  AND2X2 U2714 ( .A(\mem<19><2> ), .B(n566), .Y(n946) );
  INVX1 U2715 ( .A(n946), .Y(n947) );
  AND2X2 U2716 ( .A(\mem<45><2> ), .B(n1501), .Y(n948) );
  INVX1 U2717 ( .A(n948), .Y(n949) );
  AND2X2 U2718 ( .A(\mem<47><2> ), .B(n1433), .Y(n950) );
  INVX1 U2719 ( .A(n950), .Y(n951) );
  AND2X2 U2720 ( .A(\mem<40><2> ), .B(n483), .Y(n952) );
  INVX1 U2721 ( .A(n952), .Y(n953) );
  AND2X2 U2722 ( .A(\mem<43><2> ), .B(n17), .Y(n954) );
  INVX1 U2723 ( .A(n954), .Y(n955) );
  AND2X2 U2724 ( .A(\mem<37><2> ), .B(n543), .Y(n956) );
  INVX1 U2725 ( .A(n956), .Y(n957) );
  AND2X2 U2726 ( .A(\mem<39><2> ), .B(n1494), .Y(n958) );
  INVX1 U2727 ( .A(n958), .Y(n959) );
  AND2X2 U2728 ( .A(\mem<33><2> ), .B(n439), .Y(n960) );
  INVX1 U2729 ( .A(n960), .Y(n961) );
  AND2X2 U2730 ( .A(\mem<35><2> ), .B(n1508), .Y(n962) );
  INVX1 U2731 ( .A(n962), .Y(n963) );
  AND2X2 U2732 ( .A(\mem<29><3> ), .B(n3849), .Y(n964) );
  INVX1 U2733 ( .A(n964), .Y(n965) );
  AND2X2 U2734 ( .A(\mem<31><3> ), .B(n433), .Y(n966) );
  INVX1 U2735 ( .A(n966), .Y(n967) );
  AND2X2 U2736 ( .A(\mem<24><3> ), .B(n465), .Y(n968) );
  INVX1 U2737 ( .A(n968), .Y(n969) );
  AND2X2 U2738 ( .A(\mem<27><3> ), .B(n3901), .Y(n970) );
  INVX1 U2739 ( .A(n970), .Y(n971) );
  AND2X2 U2740 ( .A(\mem<21><3> ), .B(n461), .Y(n972) );
  INVX1 U2741 ( .A(n972), .Y(n973) );
  AND2X2 U2742 ( .A(\mem<23><3> ), .B(n437), .Y(n974) );
  INVX1 U2743 ( .A(n974), .Y(n975) );
  AND2X2 U2744 ( .A(\mem<17><3> ), .B(n77), .Y(n976) );
  INVX1 U2745 ( .A(n976), .Y(n977) );
  AND2X2 U2746 ( .A(\mem<19><3> ), .B(n566), .Y(n978) );
  INVX1 U2747 ( .A(n978), .Y(n979) );
  AND2X2 U2748 ( .A(\mem<45><3> ), .B(n1501), .Y(n980) );
  INVX1 U2749 ( .A(n980), .Y(n981) );
  AND2X2 U2750 ( .A(\mem<47><3> ), .B(n1433), .Y(n982) );
  INVX1 U2751 ( .A(n982), .Y(n983) );
  AND2X2 U2752 ( .A(\mem<40><3> ), .B(n483), .Y(n984) );
  INVX1 U2753 ( .A(n984), .Y(n985) );
  AND2X2 U2754 ( .A(\mem<43><3> ), .B(n17), .Y(n986) );
  INVX1 U2755 ( .A(n986), .Y(n987) );
  AND2X2 U2756 ( .A(\mem<37><3> ), .B(n518), .Y(n988) );
  INVX1 U2757 ( .A(n988), .Y(n989) );
  AND2X2 U2758 ( .A(\mem<39><3> ), .B(n1494), .Y(n990) );
  INVX1 U2759 ( .A(n990), .Y(n991) );
  AND2X2 U2760 ( .A(\mem<33><3> ), .B(n439), .Y(n992) );
  INVX1 U2761 ( .A(n992), .Y(n993) );
  AND2X2 U2762 ( .A(\mem<35><3> ), .B(n1508), .Y(n994) );
  INVX1 U2763 ( .A(n994), .Y(n995) );
  AND2X2 U2764 ( .A(\mem<29><4> ), .B(n3849), .Y(n996) );
  INVX1 U2765 ( .A(n996), .Y(n997) );
  AND2X2 U2766 ( .A(\mem<31><4> ), .B(n433), .Y(n998) );
  INVX1 U2767 ( .A(n998), .Y(n999) );
  AND2X2 U2768 ( .A(\mem<24><4> ), .B(n465), .Y(n1000) );
  INVX1 U2769 ( .A(n1000), .Y(n1001) );
  AND2X2 U2770 ( .A(\mem<27><4> ), .B(n3901), .Y(n1002) );
  INVX1 U2771 ( .A(n1002), .Y(n1003) );
  AND2X2 U2772 ( .A(\mem<21><4> ), .B(n461), .Y(n1004) );
  INVX1 U2773 ( .A(n1004), .Y(n1005) );
  AND2X2 U2774 ( .A(\mem<23><4> ), .B(n437), .Y(n1006) );
  INVX1 U2775 ( .A(n1006), .Y(n1007) );
  AND2X2 U2776 ( .A(\mem<17><4> ), .B(n77), .Y(n1008) );
  INVX1 U2777 ( .A(n1008), .Y(n1009) );
  AND2X2 U2778 ( .A(\mem<19><4> ), .B(n566), .Y(n1010) );
  INVX1 U2779 ( .A(n1010), .Y(n1011) );
  AND2X2 U2780 ( .A(\mem<45><4> ), .B(n1501), .Y(n1012) );
  INVX1 U2781 ( .A(n1012), .Y(n1013) );
  AND2X2 U2782 ( .A(\mem<47><4> ), .B(n1433), .Y(n1014) );
  INVX1 U2783 ( .A(n1014), .Y(n1015) );
  AND2X2 U2784 ( .A(\mem<40><4> ), .B(n483), .Y(n1016) );
  INVX1 U2785 ( .A(n1016), .Y(n1017) );
  AND2X2 U2786 ( .A(\mem<43><4> ), .B(n17), .Y(n1018) );
  INVX1 U2787 ( .A(n1018), .Y(n1019) );
  AND2X2 U2788 ( .A(\mem<37><4> ), .B(n544), .Y(n1020) );
  INVX1 U2789 ( .A(n1020), .Y(n1021) );
  AND2X2 U2790 ( .A(\mem<39><4> ), .B(n1494), .Y(n1022) );
  INVX1 U2791 ( .A(n1022), .Y(n1023) );
  AND2X2 U2792 ( .A(\mem<33><4> ), .B(n439), .Y(n1024) );
  INVX1 U2793 ( .A(n1024), .Y(n1025) );
  AND2X2 U2794 ( .A(\mem<35><4> ), .B(n1508), .Y(n1026) );
  INVX1 U2795 ( .A(n1026), .Y(n1027) );
  AND2X2 U2796 ( .A(n2647), .B(n2646), .Y(n1028) );
  INVX1 U2797 ( .A(n1028), .Y(n1029) );
  INVX1 U2798 ( .A(n106), .Y(n1030) );
  AND2X2 U2799 ( .A(n2862), .B(n2861), .Y(n1031) );
  INVX1 U2800 ( .A(n1031), .Y(n1032) );
  AND2X2 U2801 ( .A(n2608), .B(n1505), .Y(n1033) );
  INVX1 U2802 ( .A(n1033), .Y(n1034) );
  INVX1 U2803 ( .A(n1035), .Y(n1036) );
  INVX1 U2804 ( .A(n1037), .Y(n1038) );
  INVX1 U2805 ( .A(n1039), .Y(n1040) );
  INVX1 U2806 ( .A(n1041), .Y(n1042) );
  INVX1 U2807 ( .A(n1043), .Y(n1044) );
  INVX1 U2808 ( .A(n1045), .Y(n1046) );
  AND2X2 U2809 ( .A(n2962), .B(n473), .Y(n1047) );
  INVX1 U2810 ( .A(n1047), .Y(n1048) );
  INVX1 U2811 ( .A(n1049), .Y(n1050) );
  INVX1 U2812 ( .A(n1051), .Y(n1052) );
  INVX1 U2813 ( .A(n1053), .Y(n1054) );
  INVX1 U2814 ( .A(n1055), .Y(n1056) );
  INVX1 U2815 ( .A(n1057), .Y(n1058) );
  INVX1 U2816 ( .A(n1059), .Y(n1060) );
  AND2X2 U2817 ( .A(n2650), .B(n2649), .Y(n1061) );
  INVX1 U2818 ( .A(n1061), .Y(n1062) );
  INVX1 U2819 ( .A(n108), .Y(n1063) );
  AND2X2 U2820 ( .A(n2729), .B(n2728), .Y(n1064) );
  INVX1 U2821 ( .A(n1064), .Y(n1065) );
  AND2X2 U2822 ( .A(n2864), .B(n2863), .Y(n1066) );
  INVX1 U2823 ( .A(n1066), .Y(n1067) );
  AND2X2 U2824 ( .A(n1500), .B(n4586), .Y(n1068) );
  AND2X2 U2825 ( .A(n2964), .B(n4586), .Y(n1069) );
  AND2X1 U2826 ( .A(n2625), .B(n1165), .Y(n1070) );
  AND2X2 U2827 ( .A(n2598), .B(n1167), .Y(n1071) );
  AND2X2 U2828 ( .A(n2585), .B(n1171), .Y(n1073) );
  AND2X1 U2829 ( .A(n2624), .B(n1173), .Y(n1074) );
  AND2X1 U2830 ( .A(n3167), .B(n1177), .Y(n1076) );
  AND2X1 U2831 ( .A(n1478), .B(n3192), .Y(n1077) );
  AND2X1 U2832 ( .A(n3242), .B(n1179), .Y(n1078) );
  AND2X1 U2833 ( .A(n1290), .B(n1181), .Y(n1079) );
  AND2X1 U2834 ( .A(n1468), .B(n3294), .Y(n1081) );
  AND2X1 U2835 ( .A(n3322), .B(n3321), .Y(n1082) );
  AND2X1 U2836 ( .A(n1289), .B(n3348), .Y(n1083) );
  AND2X1 U2837 ( .A(n3398), .B(n1183), .Y(n1084) );
  AND2X1 U2838 ( .A(n3423), .B(n1185), .Y(n1085) );
  AND2X1 U2839 ( .A(n3448), .B(n1187), .Y(n1086) );
  AND2X1 U2840 ( .A(n3473), .B(n1189), .Y(n1087) );
  AND2X1 U2841 ( .A(n411), .B(n1191), .Y(n1088) );
  AND2X1 U2842 ( .A(n3522), .B(n1193), .Y(n1089) );
  AND2X1 U2843 ( .A(n3547), .B(n1195), .Y(n1090) );
  AND2X1 U2844 ( .A(n3572), .B(n1197), .Y(n1091) );
  AND2X1 U2845 ( .A(n3597), .B(n1199), .Y(n1092) );
  AND2X1 U2846 ( .A(n1277), .B(n1201), .Y(n1093) );
  AND2X1 U2847 ( .A(n3646), .B(n1203), .Y(n1094) );
  AND2X1 U2848 ( .A(n3671), .B(n1205), .Y(n1095) );
  AND2X1 U2849 ( .A(n3696), .B(n1207), .Y(n1096) );
  AND2X1 U2850 ( .A(n3721), .B(n1209), .Y(n1097) );
  AND2X1 U2851 ( .A(n3746), .B(n1211), .Y(n1098) );
  AND2X1 U2852 ( .A(n1213), .B(n1288), .Y(n1099) );
  AND2X1 U2853 ( .A(n1518), .B(n1215), .Y(n1100) );
  AND2X1 U2854 ( .A(n1217), .B(n1287), .Y(n1101) );
  AND2X1 U2855 ( .A(n2601), .B(n1219), .Y(n1102) );
  AND2X1 U2856 ( .A(n1453), .B(n1221), .Y(n1103) );
  AND2X1 U2857 ( .A(n1480), .B(n1223), .Y(n1104) );
  AND2X2 U2858 ( .A(n549), .B(n1225), .Y(n1105) );
  AND2X1 U2859 ( .A(n2591), .B(n1227), .Y(n1106) );
  AND2X1 U2860 ( .A(n1485), .B(n1229), .Y(n1107) );
  AND2X1 U2861 ( .A(n4003), .B(n1231), .Y(n1108) );
  AND2X1 U2862 ( .A(n4028), .B(n1233), .Y(n1109) );
  AND2X1 U2863 ( .A(n4053), .B(n1235), .Y(n1110) );
  AND2X1 U2864 ( .A(n4078), .B(n1237), .Y(n1111) );
  AND2X1 U2865 ( .A(n4103), .B(n1239), .Y(n1112) );
  AND2X1 U2866 ( .A(n4128), .B(n1241), .Y(n1113) );
  AND2X1 U2867 ( .A(n4153), .B(n1243), .Y(n1114) );
  AND2X1 U2868 ( .A(n1245), .B(n1292), .Y(n1115) );
  AND2X1 U2869 ( .A(n4202), .B(n1247), .Y(n1116) );
  AND2X1 U2870 ( .A(n1456), .B(n1249), .Y(n1117) );
  AND2X1 U2871 ( .A(n4252), .B(n1251), .Y(n1118) );
  AND2X1 U2872 ( .A(n4277), .B(n1253), .Y(n1119) );
  AND2X1 U2873 ( .A(n4302), .B(n1255), .Y(n1120) );
  AND2X1 U2874 ( .A(n4327), .B(n1257), .Y(n1121) );
  AND2X1 U2875 ( .A(n4352), .B(n1259), .Y(n1122) );
  AND2X1 U2876 ( .A(n4377), .B(n1261), .Y(n1123) );
  AND2X1 U2877 ( .A(n4402), .B(n1263), .Y(n1124) );
  AND2X1 U2878 ( .A(n1265), .B(n1291), .Y(n1125) );
  AND2X2 U2879 ( .A(n4451), .B(n1267), .Y(n1126) );
  AND2X1 U2880 ( .A(n4476), .B(n1269), .Y(n1127) );
  AND2X2 U2881 ( .A(n46), .B(n1271), .Y(n1128) );
  AND2X1 U2882 ( .A(n4526), .B(n1273), .Y(n1129) );
  AND2X2 U2883 ( .A(n4551), .B(n1275), .Y(n1130) );
  AND2X2 U2884 ( .A(n4552), .B(n4574), .Y(n1131) );
  INVX1 U2885 ( .A(n1132), .Y(n1133) );
  OR2X2 U2886 ( .A(n1443), .B(N182), .Y(n1134) );
  INVX1 U2887 ( .A(n1134), .Y(n1135) );
  AND2X2 U2888 ( .A(n16), .B(\mem<31><6> ), .Y(n1136) );
  AND2X2 U2889 ( .A(n50), .B(n33), .Y(n1137) );
  INVX1 U2890 ( .A(n1137), .Y(n1138) );
  INVX1 U2891 ( .A(n1139), .Y(n1140) );
  INVX1 U2892 ( .A(n1141), .Y(n1142) );
  INVX1 U2893 ( .A(n1143), .Y(n1144) );
  INVX1 U2894 ( .A(n1145), .Y(n1146) );
  INVX1 U2895 ( .A(n1147), .Y(n1148) );
  INVX1 U2896 ( .A(n1149), .Y(n1150) );
  AND2X2 U2897 ( .A(n1451), .B(\addr<14> ), .Y(n1151) );
  INVX1 U2898 ( .A(n1151), .Y(n1152) );
  INVX1 U2899 ( .A(n1153), .Y(n1154) );
  INVX1 U2900 ( .A(n1155), .Y(n1156) );
  INVX1 U2901 ( .A(n1157), .Y(n1158) );
  INVX1 U2902 ( .A(n1159), .Y(n1160) );
  INVX1 U2903 ( .A(n1161), .Y(n1162) );
  INVX1 U2904 ( .A(n1163), .Y(n1164) );
  INVX1 U2905 ( .A(n1165), .Y(n1166) );
  INVX1 U2906 ( .A(n1167), .Y(n1168) );
  INVX1 U2907 ( .A(n1169), .Y(n1170) );
  INVX1 U2908 ( .A(n1171), .Y(n1172) );
  INVX1 U2909 ( .A(n1173), .Y(n1174) );
  INVX1 U2910 ( .A(n1175), .Y(n1176) );
  INVX1 U2911 ( .A(n1177), .Y(n1178) );
  INVX1 U2912 ( .A(n1179), .Y(n1180) );
  INVX1 U2913 ( .A(n1181), .Y(n1182) );
  INVX1 U2914 ( .A(n1183), .Y(n1184) );
  INVX1 U2915 ( .A(n1185), .Y(n1186) );
  INVX1 U2916 ( .A(n1187), .Y(n1188) );
  INVX1 U2917 ( .A(n1189), .Y(n1190) );
  INVX1 U2918 ( .A(n1191), .Y(n1192) );
  INVX1 U2919 ( .A(n1193), .Y(n1194) );
  INVX1 U2920 ( .A(n1195), .Y(n1196) );
  INVX1 U2921 ( .A(n1197), .Y(n1198) );
  INVX1 U2922 ( .A(n1199), .Y(n1200) );
  INVX1 U2923 ( .A(n1201), .Y(n1202) );
  INVX1 U2924 ( .A(n1203), .Y(n1204) );
  INVX1 U2925 ( .A(n1205), .Y(n1206) );
  INVX1 U2926 ( .A(n1207), .Y(n1208) );
  INVX1 U2927 ( .A(n1209), .Y(n1210) );
  INVX1 U2928 ( .A(n1211), .Y(n1212) );
  INVX1 U2929 ( .A(n1213), .Y(n1214) );
  INVX1 U2930 ( .A(n1215), .Y(n1216) );
  INVX1 U2931 ( .A(n1217), .Y(n1218) );
  INVX1 U2932 ( .A(n1219), .Y(n1220) );
  INVX1 U2933 ( .A(n1221), .Y(n1222) );
  INVX1 U2934 ( .A(n1223), .Y(n1224) );
  INVX1 U2935 ( .A(n1225), .Y(n1226) );
  INVX1 U2936 ( .A(n1227), .Y(n1228) );
  INVX1 U2937 ( .A(n1229), .Y(n1230) );
  INVX1 U2938 ( .A(n1231), .Y(n1232) );
  INVX1 U2939 ( .A(n1233), .Y(n1234) );
  INVX1 U2940 ( .A(n1235), .Y(n1236) );
  INVX1 U2941 ( .A(n1237), .Y(n1238) );
  INVX1 U2942 ( .A(n1239), .Y(n1240) );
  INVX1 U2943 ( .A(n1241), .Y(n1242) );
  INVX1 U2944 ( .A(n1243), .Y(n1244) );
  INVX1 U2945 ( .A(n1245), .Y(n1246) );
  INVX1 U2946 ( .A(n1247), .Y(n1248) );
  INVX1 U2947 ( .A(n1249), .Y(n1250) );
  INVX1 U2948 ( .A(n1251), .Y(n1252) );
  INVX1 U2949 ( .A(n1253), .Y(n1254) );
  INVX1 U2950 ( .A(n1255), .Y(n1256) );
  INVX1 U2951 ( .A(n1257), .Y(n1258) );
  INVX1 U2952 ( .A(n1259), .Y(n1260) );
  INVX1 U2953 ( .A(n1261), .Y(n1262) );
  INVX1 U2954 ( .A(n1263), .Y(n1264) );
  INVX1 U2955 ( .A(n1265), .Y(n1266) );
  INVX1 U2956 ( .A(n1267), .Y(n1268) );
  INVX1 U2957 ( .A(n1269), .Y(n1270) );
  INVX1 U2958 ( .A(n1271), .Y(n1272) );
  INVX1 U2959 ( .A(n1273), .Y(n1274) );
  INVX1 U2960 ( .A(n1275), .Y(n1276) );
  INVX1 U2961 ( .A(n1494), .Y(n1277) );
  AND2X2 U2962 ( .A(n545), .B(n489), .Y(n1278) );
  INVX1 U2963 ( .A(n1278), .Y(n1279) );
  INVX1 U2964 ( .A(n1278), .Y(n1280) );
  BUFX2 U2965 ( .A(n5055), .Y(\data_out<2> ) );
  BUFX2 U2966 ( .A(n5054), .Y(\data_out<3> ) );
  INVX1 U2967 ( .A(n1283), .Y(n1284) );
  OR2X2 U2968 ( .A(n268), .B(n2695), .Y(n1285) );
  INVX1 U2969 ( .A(n1285), .Y(n1286) );
  INVX1 U2970 ( .A(n63), .Y(n1287) );
  INVX1 U2971 ( .A(n439), .Y(n1288) );
  INVX1 U2972 ( .A(n5), .Y(n1289) );
  INVX1 U2973 ( .A(n458), .Y(n1290) );
  INVX1 U2974 ( .A(n383), .Y(n1291) );
  INVX1 U2975 ( .A(n414), .Y(n1292) );
  BUFX2 U2976 ( .A(n5053), .Y(\data_out<4> ) );
  INVX1 U2977 ( .A(n1295), .Y(n1294) );
  BUFX2 U2978 ( .A(n625), .Y(n1295) );
  INVX1 U2979 ( .A(n1296), .Y(n1297) );
  INVX1 U2980 ( .A(n3039), .Y(n1298) );
  INVX1 U2981 ( .A(n1298), .Y(n1299) );
  INVX1 U2982 ( .A(n1298), .Y(n1300) );
  INVX1 U2983 ( .A(n3797), .Y(n1301) );
  INVX1 U2984 ( .A(n1301), .Y(n1302) );
  INVX1 U2985 ( .A(n1301), .Y(n1303) );
  AND2X2 U2986 ( .A(n3014), .B(n1165), .Y(n1304) );
  INVX1 U2987 ( .A(n1304), .Y(n1305) );
  AND2X1 U2988 ( .A(n428), .B(n1167), .Y(n1306) );
  INVX1 U2989 ( .A(n1306), .Y(n1307) );
  AND2X2 U2990 ( .A(n3065), .B(n1169), .Y(n1308) );
  INVX1 U2991 ( .A(n1308), .Y(n1309) );
  AND2X1 U2992 ( .A(n2602), .B(n1171), .Y(n1310) );
  INVX1 U2993 ( .A(n1310), .Y(n1311) );
  AND2X2 U2994 ( .A(n3116), .B(n1173), .Y(n1312) );
  INVX1 U2995 ( .A(n1312), .Y(n1313) );
  AND2X2 U2996 ( .A(n3141), .B(n1175), .Y(n1314) );
  INVX1 U2997 ( .A(n1314), .Y(n1315) );
  AND2X1 U2998 ( .A(n1487), .B(n1177), .Y(n1316) );
  INVX1 U2999 ( .A(n1316), .Y(n1317) );
  AND2X1 U3000 ( .A(n1477), .B(n3192), .Y(n1318) );
  INVX1 U3001 ( .A(n1318), .Y(n1319) );
  INVX1 U3002 ( .A(n1320), .Y(n1321) );
  INVX1 U3003 ( .A(n1322), .Y(n1323) );
  INVX1 U3004 ( .A(n1324), .Y(n1325) );
  AND2X1 U3005 ( .A(n1491), .B(n3294), .Y(n1326) );
  INVX1 U3006 ( .A(n1326), .Y(n1327) );
  AND2X2 U3007 ( .A(n436), .B(n3321), .Y(n1328) );
  INVX1 U3008 ( .A(n1328), .Y(n1329) );
  INVX1 U3009 ( .A(n1330), .Y(n1331) );
  AND2X1 U3010 ( .A(n1446), .B(n1183), .Y(n1332) );
  INVX1 U3011 ( .A(n1332), .Y(n1333) );
  AND2X2 U3012 ( .A(n1185), .B(n24), .Y(n1334) );
  INVX1 U3013 ( .A(n1334), .Y(n1335) );
  AND2X1 U3014 ( .A(n1460), .B(n1187), .Y(n1336) );
  INVX1 U3015 ( .A(n1336), .Y(n1337) );
  AND2X1 U3016 ( .A(n1501), .B(n1189), .Y(n1338) );
  INVX1 U3017 ( .A(n1338), .Y(n1339) );
  INVX1 U3018 ( .A(n1340), .Y(n1341) );
  INVX1 U3019 ( .A(n1342), .Y(n1343) );
  AND2X1 U3020 ( .A(n1461), .B(n1195), .Y(n1344) );
  INVX1 U3021 ( .A(n1344), .Y(n1345) );
  INVX1 U3022 ( .A(n1346), .Y(n1347) );
  INVX1 U3023 ( .A(n1348), .Y(n1349) );
  AND2X1 U3024 ( .A(n1494), .B(n1201), .Y(n1350) );
  INVX1 U3025 ( .A(n1350), .Y(n1351) );
  AND2X2 U3026 ( .A(n2592), .B(n1203), .Y(n1352) );
  INVX1 U3027 ( .A(n1352), .Y(n1353) );
  AND2X2 U3028 ( .A(n518), .B(n1205), .Y(n1354) );
  INVX1 U3029 ( .A(n1354), .Y(n1355) );
  AND2X2 U3030 ( .A(n435), .B(n1207), .Y(n1356) );
  INVX1 U3031 ( .A(n1356), .Y(n1357) );
  AND2X1 U3032 ( .A(n1508), .B(n1209), .Y(n1358) );
  INVX1 U3033 ( .A(n1358), .Y(n1359) );
  AND2X1 U3034 ( .A(n2607), .B(n1211), .Y(n1360) );
  INVX1 U3035 ( .A(n1360), .Y(n1361) );
  AND2X2 U3036 ( .A(n439), .B(n1213), .Y(n1362) );
  INVX1 U3037 ( .A(n1362), .Y(n1363) );
  INVX1 U3038 ( .A(n1364), .Y(n1365) );
  INVX1 U3039 ( .A(n1366), .Y(n1367) );
  AND2X2 U3040 ( .A(n2600), .B(n1219), .Y(n1368) );
  INVX1 U3041 ( .A(n1368), .Y(n1369) );
  AND2X2 U3042 ( .A(n3849), .B(n1221), .Y(n1370) );
  INVX1 U3043 ( .A(n1370), .Y(n1371) );
  AND2X2 U3044 ( .A(n3875), .B(n1223), .Y(n1372) );
  INVX1 U3045 ( .A(n1372), .Y(n1373) );
  AND2X2 U3046 ( .A(n3901), .B(n1225), .Y(n1374) );
  INVX1 U3047 ( .A(n1374), .Y(n1375) );
  AND2X2 U3048 ( .A(n3927), .B(n1227), .Y(n1376) );
  INVX1 U3049 ( .A(n1376), .Y(n1377) );
  AND2X2 U3050 ( .A(n3953), .B(n1229), .Y(n1378) );
  INVX1 U3051 ( .A(n1378), .Y(n1379) );
  INVX1 U3052 ( .A(n1380), .Y(n1381) );
  AND2X2 U3053 ( .A(n437), .B(n1233), .Y(n1382) );
  INVX1 U3054 ( .A(n1382), .Y(n1383) );
  AND2X2 U3055 ( .A(n496), .B(n1235), .Y(n1384) );
  INVX1 U3056 ( .A(n1384), .Y(n1385) );
  INVX1 U3057 ( .A(n1386), .Y(n1387) );
  AND2X2 U3058 ( .A(n474), .B(n1239), .Y(n1388) );
  INVX1 U3059 ( .A(n1388), .Y(n1389) );
  INVX1 U3060 ( .A(n1390), .Y(n1391) );
  AND2X2 U3061 ( .A(n533), .B(n1243), .Y(n1392) );
  INVX1 U3062 ( .A(n1392), .Y(n1393) );
  INVX1 U3063 ( .A(n1394), .Y(n1395) );
  AND2X2 U3064 ( .A(n6), .B(n1247), .Y(n1396) );
  INVX1 U3065 ( .A(n1396), .Y(n1397) );
  AND2X1 U3066 ( .A(n1442), .B(n1249), .Y(n1398) );
  INVX1 U3067 ( .A(n1398), .Y(n1399) );
  AND2X1 U3068 ( .A(n1441), .B(n1251), .Y(n1400) );
  INVX1 U3069 ( .A(n1400), .Y(n1401) );
  AND2X1 U3070 ( .A(n1436), .B(n1253), .Y(n1402) );
  INVX1 U3071 ( .A(n1402), .Y(n1403) );
  AND2X2 U3072 ( .A(n509), .B(n1255), .Y(n1404) );
  INVX1 U3073 ( .A(n1404), .Y(n1405) );
  AND2X2 U3074 ( .A(n1489), .B(n1257), .Y(n1406) );
  INVX1 U3075 ( .A(n1406), .Y(n1407) );
  AND2X1 U3076 ( .A(n1458), .B(n1259), .Y(n1408) );
  INVX1 U3077 ( .A(n1408), .Y(n1409) );
  AND2X1 U3078 ( .A(n1457), .B(n1261), .Y(n1410) );
  INVX1 U3079 ( .A(n1410), .Y(n1411) );
  AND2X2 U3080 ( .A(n490), .B(n1263), .Y(n1412) );
  INVX1 U3081 ( .A(n1412), .Y(n1413) );
  INVX1 U3082 ( .A(n1414), .Y(n1415) );
  AND2X2 U3083 ( .A(n2618), .B(n1267), .Y(n1416) );
  INVX1 U3084 ( .A(n1416), .Y(n1417) );
  INVX1 U3085 ( .A(n1418), .Y(n1419) );
  INVX1 U3086 ( .A(n1420), .Y(n1421) );
  AND2X2 U3087 ( .A(n535), .B(n1273), .Y(n1422) );
  INVX1 U3088 ( .A(n1422), .Y(n1423) );
  INVX1 U3089 ( .A(n1424), .Y(n1425) );
  INVX1 U3090 ( .A(n1426), .Y(n1427) );
  INVX1 U3091 ( .A(n1517), .Y(n1428) );
  INVX1 U3092 ( .A(n1428), .Y(n1429) );
  INVX1 U3093 ( .A(n40), .Y(n1430) );
  INVX1 U3094 ( .A(n2619), .Y(n1431) );
  INVX1 U3095 ( .A(n1431), .Y(n1432) );
  INVX1 U3096 ( .A(n3423), .Y(n1433) );
  INVX1 U3097 ( .A(N177), .Y(n1434) );
  MUX2X1 U3098 ( .B(\mem<13><0> ), .A(\mem<12><0> ), .S(n418), .Y(n1571) );
  INVX1 U3099 ( .A(n4277), .Y(n1436) );
  INVX1 U3100 ( .A(n2620), .Y(n1437) );
  INVX1 U3101 ( .A(n1437), .Y(n1438) );
  INVX1 U3102 ( .A(n2622), .Y(n1439) );
  INVX1 U3103 ( .A(n1439), .Y(n1440) );
  INVX1 U3104 ( .A(n4252), .Y(n1441) );
  MUX2X1 U3105 ( .B(\mem<33><3> ), .A(\mem<32><3> ), .S(n493), .Y(n1744) );
  INVX1 U3106 ( .A(n1456), .Y(n1442) );
  INVX8 U3107 ( .A(n2564), .Y(n2575) );
  MUX2X1 U3108 ( .B(\mem<3><1> ), .A(\mem<2><1> ), .S(n1444), .Y(n1650) );
  AND2X2 U3109 ( .A(n1472), .B(n565), .Y(n2639) );
  INVX1 U3110 ( .A(n62), .Y(n1443) );
  INVX1 U3111 ( .A(n455), .Y(n1444) );
  MUX2X1 U3112 ( .B(\mem<17><0> ), .A(\mem<16><0> ), .S(n2564), .Y(n1565) );
  MUX2X1 U3113 ( .B(\mem<1><0> ), .A(\mem<0><0> ), .S(n2565), .Y(n1583) );
  MUX2X1 U3114 ( .B(\mem<23><0> ), .A(\mem<22><0> ), .S(n2565), .Y(n1563) );
  AND2X2 U3115 ( .A(n385), .B(n44), .Y(n1445) );
  INVX1 U3116 ( .A(n1508), .Y(n3721) );
  INVX1 U3117 ( .A(n3398), .Y(n1446) );
  MUX2X1 U3118 ( .B(n2389), .A(n2388), .S(n1447), .Y(n2387) );
  MUX2X1 U3119 ( .B(n4871), .A(n4864), .S(n560), .Y(n1448) );
  INVX1 U3120 ( .A(\mem<39><5> ), .Y(n4871) );
  INVX1 U3121 ( .A(\mem<38><5> ), .Y(n4864) );
  INVX1 U3122 ( .A(n551), .Y(n3167) );
  MUX2X1 U3123 ( .B(n1806), .A(n1807), .S(n2561), .Y(n1805) );
  NAND3X1 U3124 ( .A(n2699), .B(n1286), .C(n11), .Y(n1450) );
  INVX1 U3125 ( .A(n1459), .Y(n2374) );
  BUFX2 U3126 ( .A(\addr<15> ), .Y(n1451) );
  INVX4 U3127 ( .A(n1463), .Y(n1465) );
  MUX2X1 U3128 ( .B(n2409), .A(n2410), .S(n2558), .Y(n2408) );
  INVX1 U3129 ( .A(n3849), .Y(n1453) );
  INVX1 U3130 ( .A(n2603), .Y(n1454) );
  MUX2X1 U3131 ( .B(\mem<41><0> ), .A(\mem<40><0> ), .S(n462), .Y(n1543) );
  MUX2X1 U3132 ( .B(\mem<35><0> ), .A(\mem<34><0> ), .S(n1465), .Y(n1550) );
  MUX2X1 U3133 ( .B(n1638), .A(n1637), .S(n1455), .Y(n1636) );
  MUX2X1 U3134 ( .B(\mem<47><1> ), .A(\mem<46><1> ), .S(n2562), .Y(n1608) );
  MUX2X1 U3135 ( .B(\mem<37><1> ), .A(\mem<36><1> ), .S(n560), .Y(n1613) );
  INVX1 U3136 ( .A(n377), .Y(n1456) );
  MUX2X1 U3137 ( .B(\mem<61><0> ), .A(\mem<60><0> ), .S(n1471), .Y(n1522) );
  INVX1 U3138 ( .A(n4377), .Y(n1457) );
  MUX2X1 U3139 ( .B(n1538), .A(n1537), .S(n1455), .Y(n1536) );
  INVX1 U3140 ( .A(n4352), .Y(n1458) );
  MUX2X1 U3141 ( .B(n4902), .A(n4894), .S(n560), .Y(n1459) );
  INVX1 U3142 ( .A(\mem<43><5> ), .Y(n4902) );
  INVX1 U3143 ( .A(\mem<42><5> ), .Y(n4894) );
  INVX1 U3144 ( .A(n3448), .Y(n1460) );
  INVX1 U3145 ( .A(n3547), .Y(n1461) );
  MUX2X1 U3146 ( .B(n2360), .A(n2359), .S(n1462), .Y(n2358) );
  INVX1 U3147 ( .A(n2604), .Y(n1463) );
  INVX1 U3148 ( .A(n1463), .Y(n1464) );
  AND2X2 U3149 ( .A(n1475), .B(n51), .Y(n1467) );
  INVX1 U3150 ( .A(n1491), .Y(n1468) );
  MUX2X1 U3151 ( .B(\mem<21><0> ), .A(\mem<20><0> ), .S(n2564), .Y(n1562) );
  MUX2X1 U3152 ( .B(n1770), .A(n1773), .S(n513), .Y(n1777) );
  AND2X2 U3153 ( .A(\mem<34><5> ), .B(n2586), .Y(n1469) );
  INVX1 U3154 ( .A(\addr<7> ), .Y(n1472) );
  INVX1 U3155 ( .A(n1472), .Y(n1473) );
  MUX2X1 U3156 ( .B(\mem<19><0> ), .A(\mem<18><0> ), .S(n1471), .Y(n1566) );
  MUX2X1 U3157 ( .B(\mem<43><1> ), .A(\mem<42><1> ), .S(n2562), .Y(n1611) );
  INVX1 U3158 ( .A(n68), .Y(n2683) );
  INVX4 U3159 ( .A(n1496), .Y(n2568) );
  MUX2X1 U3160 ( .B(\mem<21><7> ), .A(\mem<20><7> ), .S(n498), .Y(n2515) );
  INVX1 U3161 ( .A(n541), .Y(n1474) );
  INVX1 U3162 ( .A(n1280), .Y(n1475) );
  MUX2X1 U3163 ( .B(n1626), .A(n1625), .S(n2550), .Y(n1624) );
  AND2X2 U3164 ( .A(n2677), .B(n2676), .Y(n1476) );
  INVX1 U3165 ( .A(n437), .Y(n4028) );
  INVX1 U3166 ( .A(n1478), .Y(n1477) );
  INVX1 U3167 ( .A(n521), .Y(n1478) );
  MUX2X1 U3168 ( .B(\mem<7><0> ), .A(\mem<6><0> ), .S(n1444), .Y(n1581) );
  INVX4 U3169 ( .A(n448), .Y(n2543) );
  AND2X2 U3170 ( .A(n34), .B(n27), .Y(n1479) );
  INVX1 U3171 ( .A(n1479), .Y(n2696) );
  INVX1 U3172 ( .A(n1486), .Y(n1617) );
  BUFX2 U3173 ( .A(n1299), .Y(n2625) );
  INVX1 U3174 ( .A(n3875), .Y(n1480) );
  NAND2X1 U3175 ( .A(n2674), .B(n2675), .Y(n1481) );
  AND2X2 U3176 ( .A(n1482), .B(n565), .Y(n2676) );
  INVX1 U3177 ( .A(n1481), .Y(n1482) );
  MUX2X1 U3178 ( .B(n2331), .A(n2330), .S(n2550), .Y(n2329) );
  INVX1 U3179 ( .A(n429), .Y(n4377) );
  INVX1 U3180 ( .A(n1490), .Y(n4103) );
  INVX1 U3181 ( .A(n2547), .Y(n1519) );
  INVX1 U3182 ( .A(n3953), .Y(n1485) );
  MUX2X1 U3183 ( .B(\mem<27><1> ), .A(\mem<26><1> ), .S(n578), .Y(n1626) );
  MUX2X1 U3184 ( .B(n4844), .A(n4836), .S(n2562), .Y(n1486) );
  INVX1 U3185 ( .A(\mem<35><1> ), .Y(n4844) );
  INVX1 U3186 ( .A(\mem<34><1> ), .Y(n4836) );
  MUX2X1 U3187 ( .B(\mem<49><1> ), .A(\mem<48><1> ), .S(n459), .Y(n1600) );
  BUFX2 U3188 ( .A(n25), .Y(n1487) );
  MUX2X1 U3189 ( .B(\mem<31><1> ), .A(\mem<30><1> ), .S(n1471), .Y(n1623) );
  AND2X2 U3190 ( .A(n2634), .B(n564), .Y(n1488) );
  AND2X2 U3191 ( .A(n45), .B(n2610), .Y(n1489) );
  INVX1 U3192 ( .A(n1489), .Y(n4327) );
  INVX1 U3193 ( .A(n502), .Y(n1490) );
  INVX1 U3194 ( .A(n413), .Y(n4003) );
  BUFX2 U3195 ( .A(n524), .Y(n1491) );
  NAND2X1 U3196 ( .A(n2716), .B(n2715), .Y(n1492) );
  INVX1 U3197 ( .A(n1492), .Y(n1493) );
  BUFX2 U3198 ( .A(n379), .Y(n1494) );
  AND2X2 U3199 ( .A(n386), .B(n1454), .Y(n1495) );
  INVX1 U3200 ( .A(n2581), .Y(n1496) );
  INVX2 U3201 ( .A(n491), .Y(n2581) );
  MUX2X1 U3202 ( .B(\mem<29><1> ), .A(\mem<28><1> ), .S(n493), .Y(n1622) );
  INVX1 U3203 ( .A(n109), .Y(n1497) );
  INVX1 U3204 ( .A(n396), .Y(n1499) );
  INVX1 U3205 ( .A(n1499), .Y(n1500) );
  MUX2X1 U3206 ( .B(n1620), .A(n1619), .S(n448), .Y(n1618) );
  INVX1 U3207 ( .A(n412), .Y(n3597) );
  INVX1 U3208 ( .A(n3473), .Y(n1501) );
  INVX1 U3209 ( .A(n1445), .Y(n1502) );
  INVX1 U3210 ( .A(n1502), .Y(n1503) );
  AND2X2 U3211 ( .A(n355), .B(n570), .Y(n1504) );
  INVX1 U3212 ( .A(n24), .Y(n3423) );
  MUX2X1 U3213 ( .B(\mem<5><0> ), .A(\mem<4><0> ), .S(n1471), .Y(n1580) );
  AND2X2 U3214 ( .A(n2677), .B(n2676), .Y(n1505) );
  MUX2X1 U3215 ( .B(\mem<23><4> ), .A(\mem<22><4> ), .S(n2562), .Y(n2331) );
  INVX1 U3216 ( .A(n553), .Y(n4128) );
  INVX2 U3217 ( .A(n2604), .Y(n2605) );
  AND2X2 U3218 ( .A(n353), .B(n2611), .Y(n1506) );
  INVX1 U3219 ( .A(n1506), .Y(n4352) );
  INVX1 U3220 ( .A(n357), .Y(n4476) );
  AND2X2 U3221 ( .A(n540), .B(n3), .Y(n1507) );
  INVX1 U3222 ( .A(n470), .Y(n3522) );
  BUFX2 U3223 ( .A(n1503), .Y(n1508) );
  INVX1 U3224 ( .A(\addr<7> ), .Y(n1509) );
  INVX1 U3225 ( .A(n1509), .Y(n1510) );
  INVX1 U3226 ( .A(n1300), .Y(n3014) );
  AND2X2 U3227 ( .A(n1498), .B(n45), .Y(n1511) );
  INVX1 U3228 ( .A(n535), .Y(n4526) );
  AND2X2 U3229 ( .A(n2722), .B(n569), .Y(n1512) );
  INVX1 U3230 ( .A(n66), .Y(n4078) );
  AND2X2 U3231 ( .A(n2962), .B(n2610), .Y(n1513) );
  INVX1 U3232 ( .A(n6), .Y(n4202) );
  INVX1 U3233 ( .A(n490), .Y(n4402) );
  BUFX2 U3234 ( .A(n1297), .Y(n2624) );
  AND2X2 U3235 ( .A(n353), .B(n2722), .Y(n1514) );
  INVX1 U3236 ( .A(n533), .Y(n4153) );
  INVX1 U3237 ( .A(n405), .Y(n4277) );
  AND2X2 U3238 ( .A(n2718), .B(n1479), .Y(n1515) );
  AND2X2 U3239 ( .A(n2718), .B(n1479), .Y(n1516) );
  INVX1 U3240 ( .A(n1297), .Y(n3116) );
  INVX2 U3241 ( .A(n448), .Y(n2542) );
  AND2X2 U3242 ( .A(n485), .B(n570), .Y(n1517) );
  INVX1 U3243 ( .A(n1429), .Y(n3473) );
  INVX1 U3244 ( .A(n3772), .Y(n1518) );
  MUX2X1 U3245 ( .B(n1796), .A(n1799), .S(n1519), .Y(n1810) );
  INVX1 U3246 ( .A(n543), .Y(n3671) );
  INVX1 U3247 ( .A(n436), .Y(n3322) );
  INVX8 U3248 ( .A(n547), .Y(n2574) );
  MUX2X1 U3249 ( .B(\mem<53><4> ), .A(\mem<52><4> ), .S(n507), .Y(n1788) );
  INVX1 U3250 ( .A(n529), .Y(n2540) );
  MUX2X1 U3251 ( .B(n1522), .A(n1523), .S(n2561), .Y(n1521) );
  MUX2X1 U3252 ( .B(n1528), .A(n1529), .S(n2561), .Y(n1524) );
  MUX2X1 U3253 ( .B(n1540), .A(n1541), .S(n2552), .Y(n1539) );
  MUX2X1 U3254 ( .B(n1546), .A(n1547), .S(n2561), .Y(n1545) );
  MUX2X1 U3255 ( .B(n1549), .A(n1550), .S(n9), .Y(n1548) );
  MUX2X1 U3256 ( .B(n1568), .A(n1569), .S(n2544), .Y(n1567) );
  MUX2X1 U3257 ( .B(n1571), .A(n1572), .S(n512), .Y(n1570) );
  MUX2X1 U3258 ( .B(n1583), .A(n1584), .S(n9), .Y(n1582) );
  MUX2X1 U3259 ( .B(n1586), .A(n1587), .S(n2544), .Y(n1585) );
  MUX2X1 U3260 ( .B(n1588), .A(n1589), .S(n2608), .Y(N192) );
  MUX2X1 U3261 ( .B(n1591), .A(n1592), .S(n2561), .Y(n1590) );
  MUX2X1 U3262 ( .B(n1597), .A(n1598), .S(n2552), .Y(n1596) );
  MUX2X1 U3263 ( .B(n1600), .A(n1601), .S(n2552), .Y(n1599) );
  MUX2X1 U3264 ( .B(n1610), .A(n1611), .S(n2552), .Y(n1609) );
  MUX2X1 U3265 ( .B(n1613), .A(n1614), .S(n2557), .Y(n1612) );
  MUX2X1 U3266 ( .B(n1616), .A(n1617), .S(n2561), .Y(n1615) );
  MUX2X1 U3267 ( .B(n1628), .A(n1632), .S(n2561), .Y(n1627) );
  MUX2X1 U3268 ( .B(n1634), .A(n1635), .S(n2561), .Y(n1633) );
  MUX2X1 U3269 ( .B(n1640), .A(n1641), .S(n2552), .Y(n1639) );
  MUX2X1 U3270 ( .B(n1643), .A(n1644), .S(n2552), .Y(n1642) );
  MUX2X1 U3271 ( .B(n1646), .A(n1647), .S(n510), .Y(n1645) );
  MUX2X1 U3272 ( .B(n1652), .A(n1653), .S(n2544), .Y(n1651) );
  MUX2X1 U3273 ( .B(n1654), .A(n1655), .S(n2608), .Y(N191) );
  MUX2X1 U3274 ( .B(n1658), .A(n1659), .S(n2553), .Y(n1657) );
  MUX2X1 U3275 ( .B(n1661), .A(n1662), .S(n2553), .Y(n1660) );
  MUX2X1 U3276 ( .B(n1664), .A(n1665), .S(n2553), .Y(n1663) );
  MUX2X1 U3277 ( .B(n1667), .A(n1668), .S(n2553), .Y(n1666) );
  MUX2X1 U3278 ( .B(n1670), .A(n1671), .S(n2544), .Y(n1669) );
  MUX2X1 U3279 ( .B(n1673), .A(n1674), .S(n2553), .Y(n1672) );
  MUX2X1 U3280 ( .B(n1676), .A(n1677), .S(n2553), .Y(n1675) );
  MUX2X1 U3281 ( .B(n1679), .A(n1680), .S(n2553), .Y(n1678) );
  MUX2X1 U3282 ( .B(n1682), .A(n1683), .S(n2553), .Y(n1681) );
  MUX2X1 U3283 ( .B(n1685), .A(n1686), .S(n2544), .Y(n1684) );
  MUX2X1 U3284 ( .B(n1688), .A(n1689), .S(n2553), .Y(n1687) );
  MUX2X1 U3285 ( .B(n1691), .A(n1692), .S(n2553), .Y(n1690) );
  MUX2X1 U3286 ( .B(n1694), .A(n1695), .S(n2553), .Y(n1693) );
  MUX2X1 U3287 ( .B(n1697), .A(n1698), .S(n2553), .Y(n1696) );
  MUX2X1 U3288 ( .B(n1700), .A(n1701), .S(n2544), .Y(n1699) );
  MUX2X1 U3289 ( .B(n1703), .A(n1704), .S(n2554), .Y(n1702) );
  MUX2X1 U3290 ( .B(n1706), .A(n1707), .S(n2554), .Y(n1705) );
  MUX2X1 U3291 ( .B(n1709), .A(n1710), .S(n2554), .Y(n1708) );
  MUX2X1 U3292 ( .B(n1712), .A(n1713), .S(n2554), .Y(n1711) );
  MUX2X1 U3293 ( .B(n1715), .A(n1716), .S(n2544), .Y(n1714) );
  MUX2X1 U3294 ( .B(n1717), .A(n1718), .S(n2608), .Y(N190) );
  MUX2X1 U3295 ( .B(n1720), .A(n1721), .S(n2554), .Y(n1719) );
  MUX2X1 U3296 ( .B(n1723), .A(n1724), .S(n2554), .Y(n1722) );
  MUX2X1 U3297 ( .B(n1726), .A(n1727), .S(n2554), .Y(n1725) );
  MUX2X1 U3298 ( .B(n1729), .A(n1730), .S(n2554), .Y(n1728) );
  MUX2X1 U3299 ( .B(n1738), .A(n1739), .S(n2554), .Y(n1737) );
  MUX2X1 U3300 ( .B(n1741), .A(n1742), .S(n2554), .Y(n1740) );
  MUX2X1 U3301 ( .B(n1744), .A(n1745), .S(n2554), .Y(n1743) );
  MUX2X1 U3302 ( .B(n1750), .A(n1751), .S(n2555), .Y(n1749) );
  MUX2X1 U3303 ( .B(n1753), .A(n1754), .S(n2555), .Y(n1752) );
  MUX2X1 U3304 ( .B(n1756), .A(n1757), .S(n2555), .Y(n1755) );
  MUX2X1 U3305 ( .B(n1759), .A(n1760), .S(n2555), .Y(n1758) );
  MUX2X1 U3306 ( .B(n1762), .A(n1763), .S(n2543), .Y(n1761) );
  MUX2X1 U3307 ( .B(n1768), .A(n1769), .S(n2555), .Y(n1767) );
  MUX2X1 U3308 ( .B(n1774), .A(n1775), .S(n2555), .Y(n1773) );
  MUX2X1 U3309 ( .B(n1777), .A(n1778), .S(n2543), .Y(n1776) );
  MUX2X1 U3310 ( .B(n1779), .A(n1780), .S(n2608), .Y(N189) );
  MUX2X1 U3311 ( .B(n1782), .A(n1783), .S(n2555), .Y(n1781) );
  MUX2X1 U3312 ( .B(n1785), .A(n1786), .S(n2555), .Y(n1784) );
  MUX2X1 U3313 ( .B(n1788), .A(n1789), .S(n2555), .Y(n1787) );
  MUX2X1 U3314 ( .B(n1791), .A(n1792), .S(n2555), .Y(n1790) );
  MUX2X1 U3315 ( .B(n1794), .A(n1795), .S(n2543), .Y(n1793) );
  MUX2X1 U3316 ( .B(n1797), .A(n1798), .S(n2556), .Y(n1796) );
  MUX2X1 U3317 ( .B(n1800), .A(n1801), .S(n2556), .Y(n1799) );
  MUX2X1 U3318 ( .B(n1803), .A(n1804), .S(n2556), .Y(n1802) );
  MUX2X1 U3319 ( .B(n1812), .A(n1813), .S(n2556), .Y(n1811) );
  MUX2X1 U3320 ( .B(n1815), .A(n2328), .S(n2556), .Y(n1814) );
  MUX2X1 U3321 ( .B(n2333), .A(n2334), .S(n2556), .Y(n2332) );
  MUX2X1 U3322 ( .B(n2336), .A(n2337), .S(n2543), .Y(n2335) );
  MUX2X1 U3323 ( .B(n2339), .A(n2340), .S(n2556), .Y(n2338) );
  MUX2X1 U3324 ( .B(n2342), .A(n2343), .S(n2556), .Y(n2341) );
  MUX2X1 U3325 ( .B(n2345), .A(n2346), .S(n2556), .Y(n2344) );
  MUX2X1 U3326 ( .B(n2348), .A(n2349), .S(n2556), .Y(n2347) );
  MUX2X1 U3327 ( .B(n2351), .A(n2352), .S(n2543), .Y(n2350) );
  MUX2X1 U3328 ( .B(n2353), .A(n2354), .S(n2608), .Y(N188) );
  MUX2X1 U3329 ( .B(n2362), .A(n2363), .S(n2557), .Y(n2361) );
  MUX2X1 U3330 ( .B(n2365), .A(n2366), .S(n2557), .Y(n2364) );
  MUX2X1 U3331 ( .B(n2376), .A(n2377), .S(n2557), .Y(n2375) );
  MUX2X1 U3332 ( .B(n2379), .A(n2380), .S(n2557), .Y(n2378) );
  MUX2X1 U3333 ( .B(n2382), .A(n2383), .S(n2543), .Y(n2381) );
  MUX2X1 U3334 ( .B(n2385), .A(n2386), .S(n2557), .Y(n2384) );
  MUX2X1 U3335 ( .B(n2391), .A(n2392), .S(n2557), .Y(n2390) );
  MUX2X1 U3336 ( .B(n2394), .A(n2395), .S(n2557), .Y(n2393) );
  MUX2X1 U3337 ( .B(n2397), .A(n2398), .S(n2543), .Y(n2396) );
  MUX2X1 U3338 ( .B(n2400), .A(n2401), .S(n2559), .Y(n2399) );
  MUX2X1 U3339 ( .B(n2412), .A(n2413), .S(n2543), .Y(n2411) );
  MUX2X1 U3340 ( .B(n2414), .A(n2415), .S(n2608), .Y(N187) );
  MUX2X1 U3341 ( .B(n2417), .A(n2418), .S(n2559), .Y(n2416) );
  MUX2X1 U3342 ( .B(n2420), .A(n2421), .S(n2559), .Y(n2419) );
  MUX2X1 U3343 ( .B(n2423), .A(n2424), .S(n2559), .Y(n2422) );
  MUX2X1 U3344 ( .B(n2426), .A(n2427), .S(n2559), .Y(n2425) );
  MUX2X1 U3345 ( .B(n2429), .A(n2430), .S(n2542), .Y(n2428) );
  MUX2X1 U3346 ( .B(n2432), .A(n2433), .S(n2559), .Y(n2431) );
  MUX2X1 U3347 ( .B(n2435), .A(n2436), .S(n2559), .Y(n2434) );
  MUX2X1 U3348 ( .B(n2438), .A(n2439), .S(n2559), .Y(n2437) );
  MUX2X1 U3349 ( .B(n2441), .A(n2442), .S(n2559), .Y(n2440) );
  MUX2X1 U3350 ( .B(n2444), .A(n2445), .S(n2542), .Y(n2443) );
  MUX2X1 U3351 ( .B(n2447), .A(n2448), .S(n2558), .Y(n2446) );
  MUX2X1 U3352 ( .B(n2450), .A(n2451), .S(n2558), .Y(n2449) );
  MUX2X1 U3353 ( .B(n2453), .A(n2454), .S(n2558), .Y(n2452) );
  MUX2X1 U3354 ( .B(n2456), .A(n2457), .S(n2558), .Y(n2455) );
  MUX2X1 U3355 ( .B(n2459), .A(n2460), .S(n2542), .Y(n2458) );
  MUX2X1 U3356 ( .B(n2462), .A(n2463), .S(n2558), .Y(n2461) );
  MUX2X1 U3357 ( .B(n2468), .A(n2469), .S(n2558), .Y(n2467) );
  MUX2X1 U3358 ( .B(n2471), .A(n2472), .S(n2558), .Y(n2470) );
  MUX2X1 U3359 ( .B(n2476), .A(n2477), .S(n2608), .Y(N186) );
  MUX2X1 U3360 ( .B(n2479), .A(n2480), .S(n2558), .Y(n2478) );
  MUX2X1 U3361 ( .B(n2482), .A(n2483), .S(n2558), .Y(n2481) );
  MUX2X1 U3362 ( .B(n2485), .A(n2486), .S(n2558), .Y(n2484) );
  MUX2X1 U3363 ( .B(n2488), .A(n2489), .S(n2558), .Y(n2487) );
  MUX2X1 U3364 ( .B(n2491), .A(n2492), .S(n2542), .Y(n2490) );
  MUX2X1 U3365 ( .B(n2494), .A(n2495), .S(n2559), .Y(n2493) );
  MUX2X1 U3366 ( .B(n2497), .A(n2498), .S(n2559), .Y(n2496) );
  MUX2X1 U3367 ( .B(n2500), .A(n2501), .S(n2559), .Y(n2499) );
  MUX2X1 U3368 ( .B(n2503), .A(n2504), .S(n2559), .Y(n2502) );
  MUX2X1 U3369 ( .B(n2506), .A(n2507), .S(n2542), .Y(n2505) );
  MUX2X1 U3370 ( .B(n2509), .A(n2510), .S(n2559), .Y(n2508) );
  MUX2X1 U3371 ( .B(n2512), .A(n2513), .S(n2559), .Y(n2511) );
  MUX2X1 U3372 ( .B(n2515), .A(n2516), .S(n2559), .Y(n2514) );
  MUX2X1 U3373 ( .B(n2518), .A(n2519), .S(n2559), .Y(n2517) );
  MUX2X1 U3374 ( .B(n2521), .A(n2522), .S(n2542), .Y(n2520) );
  MUX2X1 U3375 ( .B(n2524), .A(n2525), .S(n2559), .Y(n2523) );
  MUX2X1 U3376 ( .B(n2527), .A(n2528), .S(n2559), .Y(n2526) );
  MUX2X1 U3377 ( .B(n2530), .A(n2531), .S(n2559), .Y(n2529) );
  MUX2X1 U3378 ( .B(n2533), .A(n2534), .S(n2559), .Y(n2532) );
  MUX2X1 U3379 ( .B(n2536), .A(n2537), .S(n2542), .Y(n2535) );
  MUX2X1 U3380 ( .B(n2538), .A(n2539), .S(n2608), .Y(N185) );
  MUX2X1 U3381 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n2567), .Y(n1523) );
  MUX2X1 U3382 ( .B(\mem<58><0> ), .A(\mem<59><0> ), .S(n2567), .Y(n1529) );
  MUX2X1 U3383 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n2574), .Y(n1532) );
  MUX2X1 U3384 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n2567), .Y(n1531) );
  MUX2X1 U3385 ( .B(n1533), .A(n1530), .S(n2548), .Y(n1537) );
  MUX2X1 U3386 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n522), .Y(n1544) );
  MUX2X1 U3387 ( .B(n1542), .A(n1539), .S(n2548), .Y(n1554) );
  MUX2X1 U3388 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n559), .Y(n1547) );
  MUX2X1 U3389 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n2569), .Y(n1549) );
  MUX2X1 U3390 ( .B(n1548), .A(n1545), .S(n2548), .Y(n1553) );
  MUX2X1 U3391 ( .B(n1551), .A(n1536), .S(n2541), .Y(n1589) );
  MUX2X1 U3392 ( .B(n1558), .A(n1555), .S(n2548), .Y(n1569) );
  MUX2X1 U3393 ( .B(n1564), .A(n1561), .S(n2548), .Y(n1568) );
  MUX2X1 U3394 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n2567), .Y(n1572) );
  MUX2X1 U3395 ( .B(n1573), .A(n1570), .S(n2548), .Y(n1587) );
  MUX2X1 U3396 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n2569), .Y(n1584) );
  MUX2X1 U3397 ( .B(n1585), .A(n1567), .S(n2541), .Y(n1588) );
  MUX2X1 U3398 ( .B(\mem<62><1> ), .A(\mem<63><1> ), .S(n2574), .Y(n1592) );
  MUX2X1 U3399 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n2573), .Y(n1595) );
  MUX2X1 U3400 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n2578), .Y(n1594) );
  MUX2X1 U3401 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n2579), .Y(n1598) );
  MUX2X1 U3402 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n2568), .Y(n1597) );
  MUX2X1 U3403 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n466), .Y(n1601) );
  MUX2X1 U3404 ( .B(n1599), .A(n1596), .S(n2548), .Y(n1603) );
  MUX2X1 U3405 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n2579), .Y(n1610) );
  MUX2X1 U3406 ( .B(n1609), .A(n1606), .S(n2548), .Y(n1620) );
  MUX2X1 U3407 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n2574), .Y(n1614) );
  MUX2X1 U3408 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n2573), .Y(n1616) );
  MUX2X1 U3409 ( .B(n1615), .A(n1612), .S(n2548), .Y(n1619) );
  MUX2X1 U3410 ( .B(n1618), .A(n1602), .S(n2541), .Y(n1655) );
  MUX2X1 U3411 ( .B(n1624), .A(n1621), .S(n2547), .Y(n1638) );
  MUX2X1 U3412 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n522), .Y(n1632) );
  MUX2X1 U3413 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2567), .Y(n1628) );
  MUX2X1 U3414 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n480), .Y(n1635) );
  MUX2X1 U3415 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n2573), .Y(n1634) );
  MUX2X1 U3416 ( .B(n1633), .A(n1627), .S(n2546), .Y(n1637) );
  MUX2X1 U3417 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n466), .Y(n1641) );
  MUX2X1 U3418 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n2573), .Y(n1644) );
  MUX2X1 U3419 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2573), .Y(n1643) );
  MUX2X1 U3420 ( .B(n1642), .A(n1639), .S(n2546), .Y(n1653) );
  MUX2X1 U3421 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n2574), .Y(n1647) );
  MUX2X1 U3422 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n2569), .Y(n1646) );
  MUX2X1 U3423 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n2569), .Y(n1649) );
  MUX2X1 U3424 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n2570), .Y(n1659) );
  MUX2X1 U3425 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n2574), .Y(n1658) );
  MUX2X1 U3426 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n2575), .Y(n1662) );
  MUX2X1 U3427 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n2571), .Y(n1661) );
  MUX2X1 U3428 ( .B(n1660), .A(n1657), .S(n2546), .Y(n1671) );
  MUX2X1 U3429 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n2572), .Y(n1665) );
  MUX2X1 U3430 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n2570), .Y(n1664) );
  MUX2X1 U3431 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n2570), .Y(n1668) );
  MUX2X1 U3432 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n2572), .Y(n1667) );
  MUX2X1 U3433 ( .B(n1666), .A(n1663), .S(n2547), .Y(n1670) );
  MUX2X1 U3434 ( .B(\mem<46><2> ), .A(\mem<47><2> ), .S(n2572), .Y(n1674) );
  MUX2X1 U3435 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n2571), .Y(n1673) );
  MUX2X1 U3436 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n2572), .Y(n1677) );
  MUX2X1 U3437 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n2570), .Y(n1676) );
  MUX2X1 U3438 ( .B(n1675), .A(n1672), .S(n2546), .Y(n1686) );
  MUX2X1 U3439 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n2570), .Y(n1680) );
  MUX2X1 U3440 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n2570), .Y(n1679) );
  MUX2X1 U3441 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n1452), .Y(n1683) );
  MUX2X1 U3442 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n2572), .Y(n1682) );
  MUX2X1 U3443 ( .B(n1681), .A(n1678), .S(n2546), .Y(n1685) );
  MUX2X1 U3444 ( .B(n1684), .A(n1669), .S(n2541), .Y(n1718) );
  MUX2X1 U3445 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2570), .Y(n1689) );
  MUX2X1 U3446 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1452), .Y(n1688) );
  MUX2X1 U3447 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n2572), .Y(n1692) );
  MUX2X1 U3448 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n2575), .Y(n1691) );
  MUX2X1 U3449 ( .B(n1690), .A(n1687), .S(n2547), .Y(n1701) );
  MUX2X1 U3450 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2572), .Y(n1695) );
  MUX2X1 U3451 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n2572), .Y(n1694) );
  MUX2X1 U3452 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n2573), .Y(n1698) );
  MUX2X1 U3453 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n2570), .Y(n1697) );
  MUX2X1 U3454 ( .B(n1696), .A(n1693), .S(n2546), .Y(n1700) );
  MUX2X1 U3455 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2572), .Y(n1704) );
  MUX2X1 U3456 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n2572), .Y(n1703) );
  MUX2X1 U3457 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n2572), .Y(n1707) );
  MUX2X1 U3458 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n2570), .Y(n1706) );
  MUX2X1 U3459 ( .B(n1705), .A(n1702), .S(n2546), .Y(n1716) );
  MUX2X1 U3460 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n2570), .Y(n1710) );
  MUX2X1 U3461 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n2572), .Y(n1709) );
  MUX2X1 U3462 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n2574), .Y(n1713) );
  MUX2X1 U3463 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2570), .Y(n1712) );
  MUX2X1 U3464 ( .B(n1711), .A(n1708), .S(n2547), .Y(n1715) );
  MUX2X1 U3465 ( .B(n1714), .A(n1699), .S(n2541), .Y(n1717) );
  MUX2X1 U3466 ( .B(\mem<62><3> ), .A(\mem<63><3> ), .S(n2572), .Y(n1721) );
  MUX2X1 U3467 ( .B(\mem<60><3> ), .A(\mem<61><3> ), .S(n1452), .Y(n1720) );
  MUX2X1 U3468 ( .B(\mem<58><3> ), .A(\mem<59><3> ), .S(n2570), .Y(n1724) );
  MUX2X1 U3469 ( .B(\mem<56><3> ), .A(\mem<57><3> ), .S(n2570), .Y(n1723) );
  MUX2X1 U3470 ( .B(n1722), .A(n1719), .S(n2547), .Y(n1733) );
  MUX2X1 U3471 ( .B(\mem<54><3> ), .A(\mem<55><3> ), .S(n2576), .Y(n1727) );
  MUX2X1 U3472 ( .B(\mem<52><3> ), .A(\mem<53><3> ), .S(n2574), .Y(n1726) );
  MUX2X1 U3473 ( .B(\mem<50><3> ), .A(\mem<51><3> ), .S(n2575), .Y(n1730) );
  MUX2X1 U3474 ( .B(\mem<48><3> ), .A(\mem<49><3> ), .S(n2568), .Y(n1729) );
  MUX2X1 U3475 ( .B(\mem<46><3> ), .A(\mem<47><3> ), .S(n2575), .Y(n1736) );
  MUX2X1 U3476 ( .B(\mem<44><3> ), .A(\mem<45><3> ), .S(n2574), .Y(n1735) );
  MUX2X1 U3477 ( .B(\mem<42><3> ), .A(\mem<43><3> ), .S(n466), .Y(n1739) );
  MUX2X1 U3478 ( .B(\mem<40><3> ), .A(\mem<41><3> ), .S(n2576), .Y(n1738) );
  MUX2X1 U3479 ( .B(n1737), .A(n1734), .S(n2547), .Y(n1748) );
  MUX2X1 U3480 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n2573), .Y(n1741) );
  MUX2X1 U3481 ( .B(\mem<34><3> ), .A(\mem<35><3> ), .S(n2573), .Y(n1745) );
  MUX2X1 U3482 ( .B(n1743), .A(n1740), .S(n2547), .Y(n1747) );
  MUX2X1 U3483 ( .B(n1746), .A(n1731), .S(n2541), .Y(n1780) );
  MUX2X1 U3484 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n2573), .Y(n1750) );
  MUX2X1 U3485 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2573), .Y(n1754) );
  MUX2X1 U3486 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n2570), .Y(n1753) );
  MUX2X1 U3487 ( .B(n1752), .A(n1749), .S(n2547), .Y(n1763) );
  MUX2X1 U3488 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n2575), .Y(n1757) );
  MUX2X1 U3489 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n2574), .Y(n1756) );
  MUX2X1 U3490 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n2577), .Y(n1760) );
  MUX2X1 U3491 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n2574), .Y(n1759) );
  MUX2X1 U3492 ( .B(n1758), .A(n1755), .S(n2547), .Y(n1762) );
  MUX2X1 U3493 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1435), .Y(n1766) );
  MUX2X1 U3494 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n2574), .Y(n1765) );
  MUX2X1 U3495 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n2574), .Y(n1769) );
  MUX2X1 U3496 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n2574), .Y(n1768) );
  MUX2X1 U3497 ( .B(n1767), .A(n1764), .S(n2547), .Y(n1778) );
  MUX2X1 U3498 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n2568), .Y(n1772) );
  MUX2X1 U3499 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n2576), .Y(n1771) );
  MUX2X1 U3500 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1452), .Y(n1775) );
  MUX2X1 U3501 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2574), .Y(n1774) );
  MUX2X1 U3502 ( .B(n1776), .A(n1761), .S(n2541), .Y(n1779) );
  MUX2X1 U3503 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n2573), .Y(n1783) );
  MUX2X1 U3504 ( .B(\mem<60><4> ), .A(\mem<61><4> ), .S(n2574), .Y(n1782) );
  MUX2X1 U3505 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n2568), .Y(n1786) );
  MUX2X1 U3506 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n2570), .Y(n1785) );
  MUX2X1 U3507 ( .B(n1784), .A(n1781), .S(n2547), .Y(n1795) );
  MUX2X1 U3508 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n2568), .Y(n1789) );
  MUX2X1 U3509 ( .B(\mem<50><4> ), .A(\mem<51><4> ), .S(n1435), .Y(n1792) );
  MUX2X1 U3510 ( .B(\mem<48><4> ), .A(\mem<49><4> ), .S(n2574), .Y(n1791) );
  MUX2X1 U3511 ( .B(n1790), .A(n1787), .S(n2547), .Y(n1794) );
  MUX2X1 U3512 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n2576), .Y(n1798) );
  MUX2X1 U3513 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n2576), .Y(n1797) );
  MUX2X1 U3514 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n2580), .Y(n1801) );
  MUX2X1 U3515 ( .B(\mem<40><4> ), .A(\mem<41><4> ), .S(n2576), .Y(n1800) );
  MUX2X1 U3516 ( .B(\mem<38><4> ), .A(\mem<39><4> ), .S(n2577), .Y(n1804) );
  MUX2X1 U3517 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n1452), .Y(n1803) );
  MUX2X1 U3518 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n2576), .Y(n1807) );
  MUX2X1 U3519 ( .B(\mem<32><4> ), .A(\mem<33><4> ), .S(n2576), .Y(n1806) );
  MUX2X1 U3520 ( .B(n1805), .A(n1802), .S(n2547), .Y(n1809) );
  MUX2X1 U3521 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1452), .Y(n1813) );
  MUX2X1 U3522 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n2576), .Y(n1812) );
  MUX2X1 U3523 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n2576), .Y(n2328) );
  MUX2X1 U3524 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n466), .Y(n1815) );
  MUX2X1 U3525 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2575), .Y(n2330) );
  MUX2X1 U3526 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n2580), .Y(n2334) );
  MUX2X1 U3527 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n2575), .Y(n2333) );
  MUX2X1 U3528 ( .B(n2332), .A(n2329), .S(n2547), .Y(n2336) );
  MUX2X1 U3529 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2578), .Y(n2340) );
  MUX2X1 U3530 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n2576), .Y(n2339) );
  MUX2X1 U3531 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n2570), .Y(n2343) );
  MUX2X1 U3532 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n2570), .Y(n2342) );
  MUX2X1 U3533 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n2576), .Y(n2346) );
  MUX2X1 U3534 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2575), .Y(n2345) );
  MUX2X1 U3535 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n2576), .Y(n2349) );
  MUX2X1 U3536 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n2575), .Y(n2348) );
  MUX2X1 U3537 ( .B(n2347), .A(n2344), .S(n2547), .Y(n2351) );
  MUX2X1 U3538 ( .B(n2350), .A(n2335), .S(n2541), .Y(n2353) );
  MUX2X1 U3539 ( .B(\mem<62><5> ), .A(\mem<63><5> ), .S(n2576), .Y(n2357) );
  MUX2X1 U3540 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n1452), .Y(n2356) );
  MUX2X1 U3541 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n1452), .Y(n2360) );
  MUX2X1 U3542 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n2576), .Y(n2359) );
  MUX2X1 U3543 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n1452), .Y(n2363) );
  MUX2X1 U3544 ( .B(\mem<52><5> ), .A(\mem<53><5> ), .S(n2570), .Y(n2362) );
  MUX2X1 U3545 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n2571), .Y(n2366) );
  MUX2X1 U3546 ( .B(\mem<48><5> ), .A(\mem<49><5> ), .S(n2572), .Y(n2365) );
  MUX2X1 U3547 ( .B(n2364), .A(n2361), .S(n2547), .Y(n2368) );
  MUX2X1 U3548 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n2572), .Y(n2371) );
  MUX2X1 U3549 ( .B(n2373), .A(n2370), .S(n2547), .Y(n2383) );
  MUX2X1 U3550 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n2577), .Y(n2376) );
  MUX2X1 U3551 ( .B(\mem<32><5> ), .A(\mem<33><5> ), .S(n2579), .Y(n2379) );
  MUX2X1 U3552 ( .B(n2378), .A(n2375), .S(n2547), .Y(n2382) );
  MUX2X1 U3553 ( .B(n2381), .A(n2367), .S(n2541), .Y(n2415) );
  MUX2X1 U3554 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n2577), .Y(n2386) );
  MUX2X1 U3555 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n2577), .Y(n2385) );
  MUX2X1 U3556 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n2577), .Y(n2389) );
  MUX2X1 U3557 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n2578), .Y(n2388) );
  MUX2X1 U3558 ( .B(n2387), .A(n2384), .S(n2547), .Y(n2398) );
  MUX2X1 U3559 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n2577), .Y(n2392) );
  MUX2X1 U3560 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n2577), .Y(n2395) );
  MUX2X1 U3561 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n2579), .Y(n2394) );
  MUX2X1 U3562 ( .B(n2393), .A(n2390), .S(n2547), .Y(n2397) );
  MUX2X1 U3563 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n2578), .Y(n2401) );
  MUX2X1 U3564 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n2577), .Y(n2400) );
  MUX2X1 U3565 ( .B(n2402), .A(n2399), .S(n2547), .Y(n2413) );
  MUX2X1 U3566 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n2578), .Y(n2407) );
  MUX2X1 U3567 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n2575), .Y(n2406) );
  MUX2X1 U3568 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n2579), .Y(n2410) );
  MUX2X1 U3569 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n2579), .Y(n2409) );
  MUX2X1 U3570 ( .B(n2411), .A(n2396), .S(n2541), .Y(n2414) );
  MUX2X1 U3571 ( .B(\mem<62><6> ), .A(\mem<63><6> ), .S(n2577), .Y(n2418) );
  MUX2X1 U3572 ( .B(\mem<60><6> ), .A(\mem<61><6> ), .S(n2577), .Y(n2417) );
  MUX2X1 U3573 ( .B(\mem<58><6> ), .A(\mem<59><6> ), .S(n2578), .Y(n2421) );
  MUX2X1 U3574 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n2577), .Y(n2420) );
  MUX2X1 U3575 ( .B(n2419), .A(n2416), .S(n2546), .Y(n2430) );
  MUX2X1 U3576 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n466), .Y(n2424) );
  MUX2X1 U3577 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n2578), .Y(n2423) );
  MUX2X1 U3578 ( .B(\mem<50><6> ), .A(\mem<51><6> ), .S(n466), .Y(n2427) );
  MUX2X1 U3579 ( .B(\mem<48><6> ), .A(\mem<49><6> ), .S(n2578), .Y(n2426) );
  MUX2X1 U3580 ( .B(n2425), .A(n2422), .S(n2546), .Y(n2429) );
  MUX2X1 U3581 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n2577), .Y(n2433) );
  MUX2X1 U3582 ( .B(\mem<44><6> ), .A(\mem<45><6> ), .S(n466), .Y(n2432) );
  MUX2X1 U3583 ( .B(\mem<42><6> ), .A(\mem<43><6> ), .S(n2568), .Y(n2436) );
  MUX2X1 U3584 ( .B(\mem<40><6> ), .A(\mem<41><6> ), .S(n2578), .Y(n2435) );
  MUX2X1 U3585 ( .B(n2434), .A(n2431), .S(n2546), .Y(n2445) );
  MUX2X1 U3586 ( .B(\mem<38><6> ), .A(\mem<39><6> ), .S(n2577), .Y(n2439) );
  MUX2X1 U3587 ( .B(\mem<36><6> ), .A(\mem<37><6> ), .S(n2577), .Y(n2438) );
  MUX2X1 U3588 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n2577), .Y(n2442) );
  MUX2X1 U3589 ( .B(\mem<32><6> ), .A(\mem<33><6> ), .S(n2578), .Y(n2441) );
  MUX2X1 U3590 ( .B(n2440), .A(n2437), .S(n2546), .Y(n2444) );
  MUX2X1 U3591 ( .B(n2443), .A(n2428), .S(n2541), .Y(n2477) );
  MUX2X1 U3592 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n2577), .Y(n2448) );
  MUX2X1 U3593 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n2573), .Y(n2447) );
  MUX2X1 U3594 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n2580), .Y(n2451) );
  MUX2X1 U3595 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n2580), .Y(n2450) );
  MUX2X1 U3596 ( .B(n2449), .A(n2446), .S(n2546), .Y(n2460) );
  MUX2X1 U3597 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n2580), .Y(n2454) );
  MUX2X1 U3598 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n2575), .Y(n2453) );
  MUX2X1 U3599 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n2573), .Y(n2457) );
  MUX2X1 U3600 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n2571), .Y(n2456) );
  MUX2X1 U3601 ( .B(n2455), .A(n2452), .S(n2546), .Y(n2459) );
  MUX2X1 U3602 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n2573), .Y(n2463) );
  MUX2X1 U3603 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n2571), .Y(n2462) );
  MUX2X1 U3604 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n2575), .Y(n2466) );
  MUX2X1 U3605 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n2580), .Y(n2465) );
  MUX2X1 U3606 ( .B(n2464), .A(n2461), .S(n2546), .Y(n2475) );
  MUX2X1 U3607 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n2570), .Y(n2469) );
  MUX2X1 U3608 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n2580), .Y(n2468) );
  MUX2X1 U3609 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n2580), .Y(n2472) );
  MUX2X1 U3610 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n2580), .Y(n2471) );
  MUX2X1 U3611 ( .B(n2473), .A(n2458), .S(n2541), .Y(n2476) );
  MUX2X1 U3612 ( .B(\mem<62><7> ), .A(\mem<63><7> ), .S(n2579), .Y(n2480) );
  MUX2X1 U3613 ( .B(\mem<60><7> ), .A(\mem<61><7> ), .S(n2577), .Y(n2479) );
  MUX2X1 U3614 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n2580), .Y(n2483) );
  MUX2X1 U3615 ( .B(\mem<56><7> ), .A(\mem<57><7> ), .S(n2580), .Y(n2482) );
  MUX2X1 U3616 ( .B(n2481), .A(n2478), .S(n2546), .Y(n2492) );
  MUX2X1 U3617 ( .B(\mem<54><7> ), .A(\mem<55><7> ), .S(n2580), .Y(n2486) );
  MUX2X1 U3618 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n2574), .Y(n2485) );
  MUX2X1 U3619 ( .B(\mem<50><7> ), .A(\mem<51><7> ), .S(n2575), .Y(n2489) );
  MUX2X1 U3620 ( .B(\mem<48><7> ), .A(\mem<49><7> ), .S(n2570), .Y(n2488) );
  MUX2X1 U3621 ( .B(n2487), .A(n2484), .S(n2546), .Y(n2491) );
  MUX2X1 U3622 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n2580), .Y(n2495) );
  MUX2X1 U3623 ( .B(\mem<44><7> ), .A(\mem<45><7> ), .S(n2580), .Y(n2494) );
  MUX2X1 U3624 ( .B(\mem<42><7> ), .A(\mem<43><7> ), .S(n2577), .Y(n2498) );
  MUX2X1 U3625 ( .B(\mem<40><7> ), .A(\mem<41><7> ), .S(n2580), .Y(n2497) );
  MUX2X1 U3626 ( .B(n2496), .A(n2493), .S(n2546), .Y(n2507) );
  MUX2X1 U3627 ( .B(\mem<38><7> ), .A(\mem<39><7> ), .S(n2577), .Y(n2501) );
  MUX2X1 U3628 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n2580), .Y(n2500) );
  MUX2X1 U3629 ( .B(\mem<34><7> ), .A(\mem<35><7> ), .S(n2570), .Y(n2504) );
  MUX2X1 U3630 ( .B(\mem<32><7> ), .A(\mem<33><7> ), .S(n2575), .Y(n2503) );
  MUX2X1 U3631 ( .B(n2502), .A(n2499), .S(n2546), .Y(n2506) );
  MUX2X1 U3632 ( .B(n2505), .A(n2490), .S(n2541), .Y(n2539) );
  MUX2X1 U3633 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n2576), .Y(n2510) );
  MUX2X1 U3634 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n2580), .Y(n2509) );
  MUX2X1 U3635 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n2580), .Y(n2513) );
  MUX2X1 U3636 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n2580), .Y(n2512) );
  MUX2X1 U3637 ( .B(n2511), .A(n2508), .S(n2547), .Y(n2522) );
  MUX2X1 U3638 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n2575), .Y(n2516) );
  MUX2X1 U3639 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n2573), .Y(n2519) );
  MUX2X1 U3640 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n2570), .Y(n2518) );
  MUX2X1 U3641 ( .B(n2517), .A(n2514), .S(n2547), .Y(n2521) );
  MUX2X1 U3642 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n2577), .Y(n2525) );
  MUX2X1 U3643 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n2575), .Y(n2524) );
  MUX2X1 U3644 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n2574), .Y(n2528) );
  MUX2X1 U3645 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n2576), .Y(n2527) );
  MUX2X1 U3646 ( .B(n2526), .A(n2523), .S(n2547), .Y(n2537) );
  MUX2X1 U3647 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n2574), .Y(n2531) );
  MUX2X1 U3648 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n2573), .Y(n2530) );
  MUX2X1 U3649 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n480), .Y(n2534) );
  MUX2X1 U3650 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n2571), .Y(n2533) );
  MUX2X1 U3651 ( .B(n2532), .A(n2529), .S(n2547), .Y(n2536) );
  MUX2X1 U3652 ( .B(n2535), .A(n2520), .S(n2541), .Y(n2538) );
  INVX8 U3653 ( .A(n2545), .Y(n2547) );
  INVX8 U3654 ( .A(n534), .Y(n2550) );
  INVX8 U3655 ( .A(n451), .Y(n2551) );
  INVX8 U3656 ( .A(n2549), .Y(n2552) );
  INVX8 U3657 ( .A(n2551), .Y(n2554) );
  INVX8 U3658 ( .A(n2551), .Y(n2555) );
  INVX8 U3659 ( .A(n2550), .Y(n2556) );
  INVX8 U3660 ( .A(n2550), .Y(n2558) );
  INVX8 U3661 ( .A(n2550), .Y(n2559) );
  INVX8 U3662 ( .A(n2581), .Y(n2562) );
  INVX8 U3663 ( .A(n2582), .Y(n2563) );
  INVX8 U3664 ( .A(n455), .Y(n2564) );
  INVX8 U3665 ( .A(n2582), .Y(n2565) );
  INVX8 U3666 ( .A(n2563), .Y(n2570) );
  INVX8 U3667 ( .A(n2565), .Y(n2572) );
  INVX8 U3668 ( .A(n547), .Y(n2573) );
  INVX8 U3669 ( .A(n2564), .Y(n2576) );
  INVX8 U3670 ( .A(n2563), .Y(n2577) );
  INVX8 U3671 ( .A(n2565), .Y(n2578) );
  INVX8 U3672 ( .A(n2563), .Y(n2579) );
  INVX8 U3673 ( .A(n2562), .Y(n2580) );
  INVX1 U3674 ( .A(n2588), .Y(n2583) );
  INVX1 U3675 ( .A(n2602), .Y(n2585) );
  AND2X2 U3676 ( .A(n352), .B(n1495), .Y(n2586) );
  INVX1 U3677 ( .A(n488), .Y(n3746) );
  NOR3X1 U3678 ( .A(n2719), .B(n85), .C(n582), .Y(n2587) );
  BUFX2 U3679 ( .A(N177), .Y(n2588) );
  NAND2X1 U3680 ( .A(n2717), .B(n2715), .Y(n2589) );
  AND2X2 U3681 ( .A(n548), .B(n2590), .Y(n2677) );
  INVX1 U3682 ( .A(n2589), .Y(n2590) );
  INVX1 U3683 ( .A(n3927), .Y(n2591) );
  AND2X2 U3684 ( .A(n538), .B(n2594), .Y(n2592) );
  INVX1 U3685 ( .A(n2592), .Y(n3646) );
  INVX1 U3686 ( .A(n435), .Y(n3696) );
  AND2X2 U3687 ( .A(n1454), .B(n385), .Y(n2594) );
  AND2X2 U3688 ( .A(n2677), .B(n2676), .Y(n2595) );
  AND2X2 U3689 ( .A(n438), .B(n1497), .Y(n2596) );
  INVX1 U3690 ( .A(n2597), .Y(n2598) );
  INVX1 U3691 ( .A(n2597), .Y(n2599) );
  INVX1 U3692 ( .A(n2600), .Y(n2601) );
  BUFX2 U3693 ( .A(n2584), .Y(n2602) );
  AND2X2 U3694 ( .A(n169), .B(n139), .Y(n2845) );
  NAND3X1 U3695 ( .A(n2652), .B(n548), .C(n2651), .Y(n2603) );
  INVX1 U3696 ( .A(N177), .Y(n2604) );
  AND2X2 U3697 ( .A(n538), .B(n558), .Y(n2606) );
  INVX1 U3698 ( .A(n501), .Y(n3242) );
  BUFX2 U3699 ( .A(n488), .Y(n2607) );
  BUFX2 U3700 ( .A(n36), .Y(n2608) );
  AND2X2 U3701 ( .A(n2587), .B(n537), .Y(n2609) );
  INVX1 U3702 ( .A(n496), .Y(n4053) );
  INVX1 U3703 ( .A(n375), .Y(n2610) );
  INVX1 U3704 ( .A(n375), .Y(n2611) );
  AND2X2 U3705 ( .A(n2723), .B(n376), .Y(n2614) );
  INVX1 U3706 ( .A(n1474), .Y(n4302) );
  AND2X2 U3707 ( .A(n376), .B(n537), .Y(n2615) );
  INVX1 U3708 ( .A(n2615), .Y(n4252) );
  AND2X2 U3709 ( .A(n438), .B(n540), .Y(n2616) );
  INVX1 U3710 ( .A(n2616), .Y(n3572) );
  AND2X2 U3711 ( .A(n2723), .B(n60), .Y(n2617) );
  AND2X2 U3712 ( .A(n1498), .B(n538), .Y(n2618) );
  INVX4 U3713 ( .A(n2618), .Y(n4451) );
  AND2X2 U3714 ( .A(n540), .B(n2962), .Y(n2619) );
  INVX1 U3715 ( .A(n1432), .Y(n3398) );
  INVX1 U3716 ( .A(\addr<11> ), .Y(n2652) );
  AND2X2 U3717 ( .A(n570), .B(n538), .Y(n2620) );
  INVX1 U3718 ( .A(n1438), .Y(n3448) );
  AND2X2 U3719 ( .A(n352), .B(n1497), .Y(n2621) );
  AND2X2 U3720 ( .A(n352), .B(n570), .Y(n2622) );
  INVX1 U3721 ( .A(n1440), .Y(n3547) );
  NOR2X1 U3722 ( .A(n525), .B(n531), .Y(n2640) );
  NAND3X1 U3723 ( .A(n2675), .B(n2640), .C(n2639), .Y(n2644) );
  NOR3X1 U3724 ( .A(\addr<8> ), .B(\addr<10> ), .C(n1443), .Y(n2642) );
  NOR3X1 U3725 ( .A(n80), .B(n89), .C(n1466), .Y(n2641) );
  NAND3X1 U3726 ( .A(n2642), .B(n2716), .C(n2641), .Y(n2643) );
  NAND3X1 U3727 ( .A(n455), .B(n2635), .C(n523), .Y(n2645) );
  AOI22X1 U3728 ( .A(\mem<11><0> ), .B(n1489), .C(\mem<10><0> ), .D(n1506), 
        .Y(n2647) );
  AOI22X1 U3729 ( .A(\mem<16><0> ), .B(n6), .C(\mem<9><0> ), .D(n429), .Y(
        n2646) );
  NAND3X1 U3730 ( .A(n1465), .B(n2634), .C(n534), .Y(n2648) );
  AOI22X1 U3731 ( .A(\mem<15><0> ), .B(n377), .C(\mem<14><0> ), .D(n2615), .Y(
        n2650) );
  AOI22X1 U3732 ( .A(\mem<13><0> ), .B(n405), .C(\mem<12><0> ), .D(n509), .Y(
        n2649) );
  NOR3X1 U3733 ( .A(\addr<15> ), .B(\addr<8> ), .C(n1510), .Y(n2651) );
  NOR2X1 U3734 ( .A(n43), .B(n80), .Y(n2653) );
  NAND3X1 U3735 ( .A(n28), .B(n1430), .C(n2653), .Y(n2656) );
  NOR2X1 U3736 ( .A(\addr<13> ), .B(\addr<12> ), .Y(n2654) );
  NAND2X1 U3737 ( .A(n2655), .B(n55), .Y(n2706) );
  AOI22X1 U3738 ( .A(\mem<35><0> ), .B(n56), .C(\mem<34><0> ), .D(n460), .Y(
        n2658) );
  AOI22X1 U3739 ( .A(\mem<40><0> ), .B(n412), .C(\mem<33><0> ), .D(n439), .Y(
        n2657) );
  AOI22X1 U3740 ( .A(\mem<39><0> ), .B(n379), .C(\mem<38><0> ), .D(n2592), .Y(
        n2660) );
  AOI22X1 U3741 ( .A(\mem<37><0> ), .B(n544), .C(\mem<36><0> ), .D(n435), .Y(
        n2659) );
  NOR3X1 U3742 ( .A(\addr<10> ), .B(n38), .C(n531), .Y(n2662) );
  NOR3X1 U3743 ( .A(\addr<15> ), .B(\addr<14> ), .C(n464), .Y(n2661) );
  NAND3X1 U3744 ( .A(n80), .B(n89), .C(n2636), .Y(n2664) );
  AOI22X1 U3745 ( .A(\mem<51><0> ), .B(n524), .C(\mem<50><0> ), .D(n436), .Y(
        n2666) );
  AOI22X1 U3746 ( .A(\mem<56><0> ), .B(n25), .C(\mem<49><0> ), .D(n430), .Y(
        n2665) );
  AOI22X1 U3747 ( .A(\mem<55><0> ), .B(n521), .C(\mem<54><0> ), .D(n501), .Y(
        n2668) );
  AOI22X1 U3748 ( .A(\mem<53><0> ), .B(n458), .C(\mem<52><0> ), .D(n1467), .Y(
        n2667) );
  AOI22X1 U3749 ( .A(\mem<42><0> ), .B(n2622), .C(\mem<45><0> ), .D(n1517), 
        .Y(n2671) );
  AOI22X1 U3750 ( .A(\mem<41><0> ), .B(n2616), .C(\mem<43><0> ), .D(n470), .Y(
        n2670) );
  AOI22X1 U3751 ( .A(\mem<46><0> ), .B(n2620), .C(\mem<48><0> ), .D(n30), .Y(
        n2673) );
  AOI22X1 U3752 ( .A(\mem<44><0> ), .B(n410), .C(\mem<47><0> ), .D(n1504), .Y(
        n2672) );
  NOR2X1 U3753 ( .A(\addr<12> ), .B(\addr<11> ), .Y(n2674) );
  NAND3X1 U3754 ( .A(n105), .B(n1505), .C(n584), .Y(n3140) );
  AOI21X1 U3755 ( .A(\mem<58><0> ), .B(n3116), .C(n75), .Y(n2682) );
  NAND3X1 U3756 ( .A(n105), .B(n2595), .C(n438), .Y(n3166) );
  INVX2 U3757 ( .A(n415), .Y(n3141) );
  NOR2X1 U3758 ( .A(n2683), .B(n1471), .Y(n2678) );
  NAND3X1 U3759 ( .A(n1515), .B(n1476), .C(n2678), .Y(n3797) );
  NOR2X1 U3760 ( .A(n1303), .B(n2679), .Y(n2680) );
  AOI21X1 U3761 ( .A(\mem<57><0> ), .B(n3141), .C(n2680), .Y(n2681) );
  NAND3X1 U3762 ( .A(n472), .B(n1505), .C(n538), .Y(n3039) );
  NAND3X1 U3763 ( .A(n105), .B(n1505), .C(n431), .Y(n3013) );
  NOR2X1 U3764 ( .A(n1500), .B(n2684), .Y(n2685) );
  AOI21X1 U3765 ( .A(\mem<62><0> ), .B(n3014), .C(n2685), .Y(n2689) );
  NAND3X1 U3766 ( .A(n105), .B(n2595), .C(n419), .Y(n3090) );
  NAND3X1 U3767 ( .A(n105), .B(n1505), .C(n568), .Y(n3064) );
  NOR2X1 U3768 ( .A(n2599), .B(n2686), .Y(n2687) );
  AOI21X1 U3769 ( .A(\mem<60><0> ), .B(n3065), .C(n2687), .Y(n2688) );
  NAND3X1 U3770 ( .A(n1516), .B(n568), .C(n2595), .Y(n3874) );
  NAND3X1 U3771 ( .A(n1516), .B(n584), .C(n1505), .Y(n3952) );
  AOI21X1 U3772 ( .A(\mem<29><0> ), .B(n3849), .C(n342), .Y(n2694) );
  NAND3X1 U3773 ( .A(n1515), .B(n2595), .C(n45), .Y(n3926) );
  NAND3X1 U3774 ( .A(n19), .B(n1505), .C(n438), .Y(n3978) );
  NOR2X1 U3775 ( .A(n447), .B(n2691), .Y(n2692) );
  AOI21X1 U3776 ( .A(\mem<27><0> ), .B(n3901), .C(n2692), .Y(n2693) );
  NAND3X1 U3777 ( .A(n1516), .B(n2595), .C(n537), .Y(n3848) );
  NAND2X1 U3778 ( .A(\addr<8> ), .B(n1473), .Y(n2695) );
  NAND3X1 U3779 ( .A(\addr<9> ), .B(n31), .C(\addr<10> ), .Y(n2697) );
  NOR3X1 U3780 ( .A(n1138), .B(n2697), .C(n1152), .Y(n2698) );
  NOR2X1 U3781 ( .A(n81), .B(n2700), .Y(n2701) );
  AOI21X1 U3782 ( .A(\mem<30><0> ), .B(n2600), .C(n2701), .Y(n2705) );
  NAND3X1 U3783 ( .A(n431), .B(n1515), .C(n1476), .Y(n3823) );
  NAND3X1 U3784 ( .A(n1516), .B(n419), .C(n2595), .Y(n3900) );
  NOR2X1 U3785 ( .A(n2627), .B(n2702), .Y(n2703) );
  AOI21X1 U3786 ( .A(\mem<31><0> ), .B(n63), .C(n2703), .Y(n2704) );
  NAND3X1 U3787 ( .A(n276), .B(n2707), .C(n1135), .Y(n2708) );
  OAI21X1 U3788 ( .A(n4451), .B(n2709), .C(n821), .Y(n2710) );
  OAI21X1 U3789 ( .A(n4552), .B(n2711), .C(n421), .Y(n2714) );
  OAI21X1 U3790 ( .A(n4551), .B(n2712), .C(n823), .Y(n2713) );
  NOR2X1 U3791 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n2717) );
  NAND3X1 U3792 ( .A(n2715), .B(n2716), .C(n87), .Y(n2719) );
  NOR3X1 U3793 ( .A(n85), .B(n2719), .C(n583), .Y(n2722) );
  AOI22X1 U3794 ( .A(\mem<19><0> ), .B(n567), .C(\mem<18><0> ), .D(n486), .Y(
        n2721) );
  AOI22X1 U3795 ( .A(\mem<24><0> ), .B(n413), .C(\mem<17><0> ), .D(n414), .Y(
        n2720) );
  AOI22X1 U3796 ( .A(\mem<23><0> ), .B(n403), .C(\mem<22><0> ), .D(n2609), .Y(
        n2725) );
  AOI22X1 U3797 ( .A(\mem<21><0> ), .B(n66), .C(\mem<20><0> ), .D(n474), .Y(
        n2724) );
  AOI21X1 U3798 ( .A(n84), .B(n359), .C(n2623), .Y(\data_out<0> ) );
  AOI22X1 U3799 ( .A(\mem<11><1> ), .B(n1489), .C(\mem<10><1> ), .D(n1506), 
        .Y(n2727) );
  AOI22X1 U3800 ( .A(\mem<15><1> ), .B(n4203), .C(\mem<14><1> ), .D(n2615), 
        .Y(n2729) );
  AOI22X1 U3801 ( .A(\mem<13><1> ), .B(n405), .C(\mem<12><1> ), .D(n1474), .Y(
        n2728) );
  AOI22X1 U3802 ( .A(\mem<35><1> ), .B(n56), .C(\mem<34><1> ), .D(n460), .Y(
        n2731) );
  AOI22X1 U3803 ( .A(\mem<40><1> ), .B(n412), .C(\mem<33><1> ), .D(n439), .Y(
        n2730) );
  AOI22X1 U3804 ( .A(\mem<39><1> ), .B(n379), .C(\mem<38><1> ), .D(n2592), .Y(
        n2733) );
  AOI22X1 U3805 ( .A(\mem<37><1> ), .B(n12), .C(\mem<36><1> ), .D(n435), .Y(
        n2732) );
  AOI22X1 U3806 ( .A(\mem<51><1> ), .B(n64), .C(\mem<50><1> ), .D(n436), .Y(
        n2735) );
  AOI22X1 U3807 ( .A(\mem<56><1> ), .B(n551), .C(\mem<49><1> ), .D(n430), .Y(
        n2734) );
  AOI22X1 U3808 ( .A(\mem<55><1> ), .B(n520), .C(\mem<54><1> ), .D(n501), .Y(
        n2737) );
  AOI22X1 U3809 ( .A(\mem<53><1> ), .B(n458), .C(\mem<52><1> ), .D(n1467), .Y(
        n2736) );
  AOI22X1 U3810 ( .A(\mem<42><1> ), .B(n32), .C(\mem<45><1> ), .D(n1517), .Y(
        n2739) );
  AOI22X1 U3811 ( .A(\mem<41><1> ), .B(n2616), .C(\mem<43><1> ), .D(n470), .Y(
        n2738) );
  AOI22X1 U3812 ( .A(\mem<46><1> ), .B(n21), .C(\mem<48><1> ), .D(n30), .Y(
        n2741) );
  AOI22X1 U3813 ( .A(\mem<44><1> ), .B(n410), .C(\mem<47><1> ), .D(n1504), .Y(
        n2740) );
  AOI21X1 U3814 ( .A(\mem<58><1> ), .B(n3116), .C(n344), .Y(n2746) );
  NOR2X1 U3815 ( .A(n1303), .B(n2743), .Y(n2744) );
  AOI21X1 U3816 ( .A(\mem<57><1> ), .B(n3141), .C(n2744), .Y(n2745) );
  NOR2X1 U3817 ( .A(n1500), .B(n2747), .Y(n2748) );
  AOI21X1 U3818 ( .A(\mem<62><1> ), .B(n3014), .C(n2748), .Y(n2752) );
  NOR2X1 U3819 ( .A(n2598), .B(n2749), .Y(n2750) );
  AOI21X1 U3820 ( .A(\mem<60><1> ), .B(n3065), .C(n2750), .Y(n2751) );
  AOI21X1 U3821 ( .A(\mem<29><1> ), .B(n3849), .C(n346), .Y(n2757) );
  NOR2X1 U3822 ( .A(n447), .B(n2754), .Y(n2755) );
  AOI21X1 U3823 ( .A(\mem<27><1> ), .B(n3901), .C(n2755), .Y(n2756) );
  NOR2X1 U3824 ( .A(n409), .B(n2758), .Y(n2759) );
  AOI21X1 U3825 ( .A(\mem<30><1> ), .B(n2600), .C(n2759), .Y(n2762) );
  AOI21X1 U3826 ( .A(\mem<31><1> ), .B(n63), .C(n2760), .Y(n2761) );
  OAI21X1 U3827 ( .A(n46), .B(n2763), .C(n825), .Y(n2766) );
  OAI21X1 U3828 ( .A(n4451), .B(n2764), .C(n827), .Y(n2765) );
  NAND2X1 U3829 ( .A(\mem<8><1> ), .B(n490), .Y(n2767) );
  OAI21X1 U3830 ( .A(n4552), .B(n2768), .C(n2767), .Y(n2771) );
  OAI21X1 U3831 ( .A(n4551), .B(n2769), .C(n829), .Y(n2770) );
  AOI22X1 U3832 ( .A(\mem<19><1> ), .B(n567), .C(\mem<18><1> ), .D(n486), .Y(
        n2773) );
  AOI22X1 U3833 ( .A(\mem<24><1> ), .B(n413), .C(\mem<17><1> ), .D(n414), .Y(
        n2772) );
  AOI22X1 U3834 ( .A(\mem<23><1> ), .B(n403), .C(\mem<22><1> ), .D(n2609), .Y(
        n2775) );
  AOI22X1 U3835 ( .A(\mem<21><1> ), .B(n67), .C(\mem<20><1> ), .D(n1490), .Y(
        n2774) );
  AOI21X1 U3836 ( .A(n69), .B(n58), .C(n2623), .Y(\data_out<1> ) );
  AOI22X1 U3837 ( .A(\mem<24><5> ), .B(n413), .C(\mem<21><5> ), .D(n67), .Y(
        n2776) );
  AOI22X1 U3838 ( .A(\mem<19><5> ), .B(n567), .C(\mem<25><5> ), .D(n3953), .Y(
        n2778) );
  AOI22X1 U3839 ( .A(\mem<22><5> ), .B(n2609), .C(\mem<17><5> ), .D(n414), .Y(
        n2777) );
  AOI22X1 U3840 ( .A(\mem<12><5> ), .B(n2614), .C(\mem<10><5> ), .D(n1506), 
        .Y(n2780) );
  AOI22X1 U3841 ( .A(\mem<16><5> ), .B(n504), .C(\mem<9><5> ), .D(n429), .Y(
        n2779) );
  AOI22X1 U3842 ( .A(\mem<13><5> ), .B(n405), .C(\mem<23><5> ), .D(n403), .Y(
        n2782) );
  AOI22X1 U3843 ( .A(\mem<14><5> ), .B(n2615), .C(\mem<11><5> ), .D(n1489), 
        .Y(n2781) );
  AOI21X1 U3844 ( .A(\mem<61><5> ), .B(n2597), .C(n2784), .Y(n2788) );
  NOR2X1 U3845 ( .A(n415), .B(n2785), .Y(n2786) );
  AOI21X1 U3846 ( .A(\mem<59><5> ), .B(n2584), .C(n2786), .Y(n2787) );
  NOR2X1 U3847 ( .A(n1299), .B(n2789), .Y(n2790) );
  AOI21X1 U3848 ( .A(\mem<1><5> ), .B(n2596), .C(n2790), .Y(n2794) );
  NOR2X1 U3849 ( .A(n442), .B(n2791), .Y(n2792) );
  AOI21X1 U3850 ( .A(\mem<63><5> ), .B(n2964), .C(n2792), .Y(n2793) );
  NOR2X1 U3851 ( .A(n416), .B(n2795), .Y(n2796) );
  AOI21X1 U3852 ( .A(\mem<28><5> ), .B(n3875), .C(n2796), .Y(n2800) );
  NOR2X1 U3853 ( .A(n550), .B(n2797), .Y(n2798) );
  AOI21X1 U3854 ( .A(\mem<26><5> ), .B(n3927), .C(n2798), .Y(n2799) );
  NAND2X1 U3855 ( .A(\mem<30><5> ), .B(n432), .Y(n2802) );
  AOI22X1 U3856 ( .A(\mem<0><5> ), .B(n82), .C(\mem<32><5> ), .D(n3772), .Y(
        n2801) );
  AOI22X1 U3857 ( .A(\mem<39><5> ), .B(n379), .C(\mem<36><5> ), .D(n2593), .Y(
        n2803) );
  AOI22X1 U3858 ( .A(\mem<37><5> ), .B(n543), .C(\mem<44><5> ), .D(n410), .Y(
        n2805) );
  AOI22X1 U3859 ( .A(\mem<40><5> ), .B(n412), .C(\mem<38><5> ), .D(n2592), .Y(
        n2804) );
  AOI22X1 U3860 ( .A(\mem<3><5> ), .B(n572), .C(\mem<5><5> ), .D(n357), .Y(
        n2807) );
  AOI22X1 U3861 ( .A(\mem<2><5> ), .B(n2621), .C(\mem<7><5> ), .D(n383), .Y(
        n2806) );
  AOI22X1 U3862 ( .A(\mem<4><5> ), .B(n2617), .C(\mem<33><5> ), .D(n3747), .Y(
        n2809) );
  AOI22X1 U3863 ( .A(\mem<6><5> ), .B(n2618), .C(\mem<8><5> ), .D(n490), .Y(
        n2808) );
  AOI22X1 U3864 ( .A(\mem<51><5> ), .B(n3320), .C(\mem<53><5> ), .D(n457), .Y(
        n2811) );
  AOI22X1 U3865 ( .A(\mem<56><5> ), .B(n1), .C(\mem<52><5> ), .D(n1467), .Y(
        n2810) );
  AOI22X1 U3866 ( .A(\mem<55><5> ), .B(n520), .C(\mem<15><5> ), .D(n4203), .Y(
        n2813) );
  AOI22X1 U3867 ( .A(\mem<54><5> ), .B(n2606), .C(\mem<50><5> ), .D(n1520), 
        .Y(n2812) );
  AOI22X1 U3868 ( .A(\mem<48><5> ), .B(n2619), .C(\mem<47><5> ), .D(n1504), 
        .Y(n2815) );
  AOI22X1 U3869 ( .A(\mem<42><5> ), .B(n2622), .C(\mem<43><5> ), .D(n469), .Y(
        n2814) );
  AOI22X1 U3870 ( .A(\mem<45><5> ), .B(n1517), .C(\mem<49><5> ), .D(n430), .Y(
        n2817) );
  AOI22X1 U3871 ( .A(\mem<46><5> ), .B(n2620), .C(\mem<41><5> ), .D(n2616), 
        .Y(n2816) );
  AOI21X1 U3872 ( .A(n73), .B(n59), .C(n2623), .Y(\data_out<5> ) );
  AOI22X1 U3873 ( .A(\mem<18><6> ), .B(n2), .C(\mem<20><6> ), .D(n1490), .Y(
        n2819) );
  AOI22X1 U3874 ( .A(\mem<24><6> ), .B(n413), .C(\mem<21><6> ), .D(n79), .Y(
        n2818) );
  AOI22X1 U3875 ( .A(\mem<19><6> ), .B(n567), .C(\mem<25><6> ), .D(n3953), .Y(
        n2821) );
  AOI22X1 U3876 ( .A(\mem<22><6> ), .B(n2609), .C(\mem<17><6> ), .D(n414), .Y(
        n2820) );
  AOI22X1 U3877 ( .A(\mem<12><6> ), .B(n2614), .C(\mem<10><6> ), .D(n1506), 
        .Y(n2823) );
  AOI22X1 U3878 ( .A(\mem<16><6> ), .B(n6), .C(\mem<9><6> ), .D(n429), .Y(
        n2822) );
  AOI22X1 U3879 ( .A(\mem<13><6> ), .B(n405), .C(\mem<23><6> ), .D(n403), .Y(
        n2825) );
  AOI22X1 U3880 ( .A(\mem<14><6> ), .B(n2615), .C(\mem<11><6> ), .D(n1489), 
        .Y(n2824) );
  AOI21X1 U3881 ( .A(\mem<61><6> ), .B(n2597), .C(n2826), .Y(n2830) );
  NOR2X1 U3882 ( .A(n415), .B(n2827), .Y(n2828) );
  AOI21X1 U3883 ( .A(\mem<59><6> ), .B(n3091), .C(n2828), .Y(n2829) );
  NOR2X1 U3884 ( .A(n1299), .B(n2831), .Y(n2832) );
  AOI21X1 U3885 ( .A(\mem<1><6> ), .B(n2596), .C(n2832), .Y(n2836) );
  NOR2X1 U3886 ( .A(n442), .B(n2833), .Y(n2834) );
  AOI21X1 U3887 ( .A(\mem<63><6> ), .B(n2964), .C(n2834), .Y(n2835) );
  NOR2X1 U3888 ( .A(n416), .B(n2837), .Y(n2838) );
  AOI21X1 U3889 ( .A(\mem<28><6> ), .B(n3875), .C(n2838), .Y(n2842) );
  NOR2X1 U3890 ( .A(n549), .B(n2839), .Y(n2840) );
  AOI21X1 U3891 ( .A(\mem<26><6> ), .B(n3927), .C(n2840), .Y(n2841) );
  NAND2X1 U3892 ( .A(\mem<30><6> ), .B(n2600), .Y(n2844) );
  AOI22X1 U3893 ( .A(\mem<0><6> ), .B(n561), .C(\mem<32><6> ), .D(n476), .Y(
        n2843) );
  AOI22X1 U3894 ( .A(\mem<39><6> ), .B(n379), .C(\mem<36><6> ), .D(n2593), .Y(
        n2846) );
  AOI22X1 U3895 ( .A(\mem<37><6> ), .B(n544), .C(\mem<44><6> ), .D(n410), .Y(
        n2848) );
  AOI22X1 U3896 ( .A(\mem<40><6> ), .B(n412), .C(\mem<38><6> ), .D(n2592), .Y(
        n2847) );
  AOI22X1 U3897 ( .A(\mem<3><6> ), .B(n574), .C(\mem<5><6> ), .D(n357), .Y(
        n2850) );
  AOI22X1 U3898 ( .A(\mem<2><6> ), .B(n2621), .C(\mem<7><6> ), .D(n383), .Y(
        n2849) );
  AOI22X1 U3899 ( .A(\mem<4><6> ), .B(n2617), .C(\mem<33><6> ), .D(n3747), .Y(
        n2852) );
  AOI22X1 U3900 ( .A(\mem<6><6> ), .B(n2618), .C(\mem<8><6> ), .D(n490), .Y(
        n2851) );
  AOI22X1 U3901 ( .A(\mem<51><6> ), .B(n380), .C(\mem<53><6> ), .D(n457), .Y(
        n2854) );
  AOI22X1 U3902 ( .A(\mem<56><6> ), .B(n1449), .C(\mem<52><6> ), .D(n1467), 
        .Y(n2853) );
  AOI22X1 U3903 ( .A(\mem<55><6> ), .B(n520), .C(\mem<15><6> ), .D(n377), .Y(
        n2856) );
  AOI22X1 U3904 ( .A(\mem<54><6> ), .B(n2606), .C(\mem<50><6> ), .D(n1520), 
        .Y(n2855) );
  AOI22X1 U3905 ( .A(\mem<48><6> ), .B(n2619), .C(\mem<47><6> ), .D(n1504), 
        .Y(n2858) );
  AOI22X1 U3906 ( .A(\mem<42><6> ), .B(n2622), .C(\mem<43><6> ), .D(n469), .Y(
        n2857) );
  AOI22X1 U3907 ( .A(\mem<45><6> ), .B(n1517), .C(\mem<49><6> ), .D(n430), .Y(
        n2860) );
  AOI22X1 U3908 ( .A(\mem<46><6> ), .B(n2620), .C(\mem<41><6> ), .D(n2616), 
        .Y(n2859) );
  AOI21X1 U3909 ( .A(n76), .B(n86), .C(n2623), .Y(\data_out<6> ) );
  AOI22X1 U3910 ( .A(\mem<11><7> ), .B(n1489), .C(\mem<10><7> ), .D(n1506), 
        .Y(n2862) );
  AOI22X1 U3911 ( .A(\mem<16><7> ), .B(n6), .C(\mem<9><7> ), .D(n429), .Y(
        n2861) );
  AOI22X1 U3912 ( .A(\mem<15><7> ), .B(n377), .C(\mem<14><7> ), .D(n2615), .Y(
        n2864) );
  AOI22X1 U3913 ( .A(\mem<13><7> ), .B(n405), .C(\mem<12><7> ), .D(n1474), .Y(
        n2863) );
  AOI22X1 U3914 ( .A(\mem<35><7> ), .B(n1503), .C(\mem<34><7> ), .D(n488), .Y(
        n2866) );
  AOI22X1 U3915 ( .A(\mem<40><7> ), .B(n412), .C(\mem<33><7> ), .D(n439), .Y(
        n2865) );
  AOI22X1 U3916 ( .A(\mem<39><7> ), .B(n379), .C(\mem<38><7> ), .D(n2592), .Y(
        n2868) );
  AOI22X1 U3917 ( .A(\mem<37><7> ), .B(n518), .C(\mem<36><7> ), .D(n435), .Y(
        n2867) );
  AOI22X1 U3918 ( .A(\mem<51><7> ), .B(n524), .C(\mem<50><7> ), .D(n436), .Y(
        n2870) );
  AOI22X1 U3919 ( .A(\mem<56><7> ), .B(n1), .C(\mem<49><7> ), .D(n5), .Y(n2869) );
  AOI22X1 U3920 ( .A(\mem<55><7> ), .B(n521), .C(\mem<54><7> ), .D(n501), .Y(
        n2872) );
  AOI22X1 U3921 ( .A(\mem<53><7> ), .B(n458), .C(\mem<52><7> ), .D(n1467), .Y(
        n2871) );
  AOI22X1 U3922 ( .A(\mem<42><7> ), .B(n1440), .C(\mem<45><7> ), .D(n1429), 
        .Y(n2874) );
  AOI22X1 U3923 ( .A(\mem<41><7> ), .B(n2616), .C(\mem<43><7> ), .D(n470), .Y(
        n2873) );
  AOI22X1 U3924 ( .A(\mem<46><7> ), .B(n1438), .C(\mem<48><7> ), .D(n1432), 
        .Y(n2876) );
  AOI22X1 U3925 ( .A(\mem<44><7> ), .B(n410), .C(\mem<47><7> ), .D(n24), .Y(
        n2875) );
  AOI21X1 U3926 ( .A(\mem<58><7> ), .B(n3116), .C(n54), .Y(n2881) );
  NOR2X1 U3927 ( .A(n1303), .B(n2878), .Y(n2879) );
  AOI21X1 U3928 ( .A(\mem<57><7> ), .B(n3141), .C(n2879), .Y(n2880) );
  NOR2X1 U3929 ( .A(n1500), .B(n2882), .Y(n2883) );
  AOI21X1 U3930 ( .A(\mem<62><7> ), .B(n3014), .C(n2883), .Y(n2887) );
  NOR2X1 U3931 ( .A(n2598), .B(n2884), .Y(n2885) );
  AOI21X1 U3932 ( .A(\mem<60><7> ), .B(n3065), .C(n2885), .Y(n2886) );
  NOR2X1 U3933 ( .A(n2591), .B(n2888), .Y(n2889) );
  AOI21X1 U3934 ( .A(\mem<29><7> ), .B(n3849), .C(n2889), .Y(n2893) );
  NOR2X1 U3935 ( .A(n447), .B(n2890), .Y(n2891) );
  AOI21X1 U3936 ( .A(\mem<27><7> ), .B(n3901), .C(n2891), .Y(n2892) );
  NOR2X1 U3937 ( .A(n409), .B(n2894), .Y(n2895) );
  AOI21X1 U3938 ( .A(\mem<30><7> ), .B(n2600), .C(n2895), .Y(n2899) );
  NOR2X1 U3939 ( .A(n2627), .B(n2896), .Y(n2897) );
  AOI21X1 U3940 ( .A(\mem<31><7> ), .B(n63), .C(n2897), .Y(n2898) );
  OAI21X1 U3941 ( .A(n46), .B(n2900), .C(n831), .Y(n2903) );
  OAI21X1 U3942 ( .A(n4451), .B(n2901), .C(n833), .Y(n2902) );
  NAND2X1 U3943 ( .A(\mem<8><7> ), .B(n490), .Y(n2904) );
  OAI21X1 U3944 ( .A(n4552), .B(n2905), .C(n2904), .Y(n2908) );
  OAI21X1 U3945 ( .A(n4551), .B(n2906), .C(n835), .Y(n2907) );
  AOI22X1 U3946 ( .A(\mem<19><7> ), .B(n553), .C(\mem<18><7> ), .D(n533), .Y(
        n2910) );
  AOI22X1 U3947 ( .A(\mem<24><7> ), .B(n413), .C(\mem<17><7> ), .D(n414), .Y(
        n2909) );
  AOI22X1 U3948 ( .A(\mem<23><7> ), .B(n437), .C(\mem<22><7> ), .D(n496), .Y(
        n2912) );
  AOI22X1 U3949 ( .A(\mem<21><7> ), .B(n79), .C(\mem<20><7> ), .D(n474), .Y(
        n2911) );
  NAND3X1 U3950 ( .A(n350), .B(n363), .C(n133), .Y(n2913) );
  AOI21X1 U3951 ( .A(n127), .B(n135), .C(n2623), .Y(\data_out<7> ) );
  AND2X2 U3952 ( .A(N192), .B(n393), .Y(\data_out<8> ) );
  AND2X2 U3953 ( .A(N191), .B(n393), .Y(\data_out<9> ) );
  AND2X2 U3954 ( .A(N190), .B(n393), .Y(\data_out<10> ) );
  AND2X2 U3955 ( .A(N189), .B(n393), .Y(\data_out<11> ) );
  AND2X2 U3956 ( .A(N188), .B(n393), .Y(\data_out<12> ) );
  AND2X2 U3957 ( .A(N187), .B(n393), .Y(\data_out<13> ) );
  AND2X2 U3958 ( .A(N186), .B(n393), .Y(\data_out<14> ) );
  AND2X2 U3959 ( .A(N185), .B(n393), .Y(\data_out<15> ) );
  OAI21X1 U3960 ( .A(n4302), .B(n4674), .C(n837), .Y(n2915) );
  OAI21X1 U3961 ( .A(n4252), .B(n4690), .C(n839), .Y(n2914) );
  OAI21X1 U3962 ( .A(n4402), .B(n4642), .C(n841), .Y(n2917) );
  OAI21X1 U3963 ( .A(n4352), .B(n4658), .C(n843), .Y(n2916) );
  OAI21X1 U3964 ( .A(n46), .B(n4614), .C(n845), .Y(n2919) );
  OAI21X1 U3965 ( .A(n4451), .B(n4628), .C(n847), .Y(n2918) );
  OAI21X1 U3966 ( .A(n4552), .B(n4596), .C(n849), .Y(n2921) );
  OAI21X1 U3967 ( .A(n4551), .B(n4601), .C(n851), .Y(n2920) );
  OAI21X1 U3968 ( .A(n2626), .B(n5034), .C(n853), .Y(n2923) );
  OAI21X1 U3969 ( .A(n2625), .B(n5045), .C(n855), .Y(n2922) );
  OAI21X1 U3970 ( .A(n444), .B(n5015), .C(n857), .Y(n2925) );
  OAI21X1 U3971 ( .A(n2624), .B(n5022), .C(n859), .Y(n2924) );
  OAI21X1 U3972 ( .A(n3268), .B(n4977), .C(n861), .Y(n2927) );
  OAI21X1 U3973 ( .A(n3242), .B(n4993), .C(n863), .Y(n2926) );
  OAI21X1 U3974 ( .A(n3398), .B(n4945), .C(n865), .Y(n2929) );
  OAI21X1 U3975 ( .A(n3322), .B(n4961), .C(n867), .Y(n2928) );
  OAI21X1 U3976 ( .A(n4302), .B(n4673), .C(n869), .Y(n2931) );
  OAI21X1 U3977 ( .A(n4252), .B(n4689), .C(n871), .Y(n2930) );
  OAI21X1 U3978 ( .A(n4402), .B(n4641), .C(n873), .Y(n2933) );
  OAI21X1 U3979 ( .A(n4352), .B(n4657), .C(n875), .Y(n2932) );
  OAI21X1 U3980 ( .A(n46), .B(n4613), .C(n877), .Y(n2935) );
  OAI21X1 U3981 ( .A(n4451), .B(n4627), .C(n879), .Y(n2934) );
  OAI21X1 U3982 ( .A(n4552), .B(n4595), .C(n881), .Y(n2937) );
  OAI21X1 U3983 ( .A(n4551), .B(n4600), .C(n883), .Y(n2936) );
  OAI21X1 U3984 ( .A(n2626), .B(n5033), .C(n885), .Y(n2939) );
  OAI21X1 U3985 ( .A(n2625), .B(n5044), .C(n887), .Y(n2938) );
  OAI21X1 U3986 ( .A(n444), .B(n5014), .C(n889), .Y(n2941) );
  OAI21X1 U3987 ( .A(n2624), .B(n5021), .C(n891), .Y(n2940) );
  OAI21X1 U3988 ( .A(n3268), .B(n4976), .C(n893), .Y(n2943) );
  OAI21X1 U3989 ( .A(n3242), .B(n4992), .C(n895), .Y(n2942) );
  OAI21X1 U3990 ( .A(n3398), .B(n4944), .C(n897), .Y(n2945) );
  OAI21X1 U3991 ( .A(n3322), .B(n4960), .C(n899), .Y(n2944) );
  OAI21X1 U3992 ( .A(n4302), .B(n4672), .C(n901), .Y(n2947) );
  OAI21X1 U3993 ( .A(n4252), .B(n4688), .C(n903), .Y(n2946) );
  OAI21X1 U3994 ( .A(n4402), .B(n4640), .C(n905), .Y(n2949) );
  OAI21X1 U3995 ( .A(n4352), .B(n4656), .C(n907), .Y(n2948) );
  OAI21X1 U3996 ( .A(n46), .B(n4612), .C(n909), .Y(n2951) );
  OAI21X1 U3997 ( .A(n4451), .B(n4626), .C(n911), .Y(n2950) );
  OAI21X1 U3998 ( .A(n4552), .B(n4594), .C(n913), .Y(n2953) );
  OAI21X1 U3999 ( .A(n4551), .B(n4599), .C(n915), .Y(n2952) );
  OAI21X1 U4000 ( .A(n2626), .B(n5032), .C(n917), .Y(n2955) );
  OAI21X1 U4001 ( .A(n2625), .B(n5043), .C(n919), .Y(n2954) );
  OAI21X1 U4002 ( .A(n444), .B(n5013), .C(n921), .Y(n2957) );
  OAI21X1 U4003 ( .A(n2624), .B(n5020), .C(n923), .Y(n2956) );
  OAI21X1 U4004 ( .A(n3268), .B(n4975), .C(n925), .Y(n2959) );
  OAI21X1 U4005 ( .A(n3242), .B(n4991), .C(n927), .Y(n2958) );
  OAI21X1 U4006 ( .A(n3398), .B(n4943), .C(n929), .Y(n2961) );
  OAI21X1 U4007 ( .A(n3322), .B(n4959), .C(n931), .Y(n2960) );
  OAI21X1 U4008 ( .A(n1133), .B(n2964), .C(n1294), .Y(n2963) );
  AOI22X1 U4009 ( .A(\data_in<15> ), .B(n1068), .C(\data_in<7> ), .D(n1069), 
        .Y(n608) );
  AOI22X1 U4010 ( .A(\data_in<14> ), .B(n1068), .C(\data_in<6> ), .D(n1069), 
        .Y(n607) );
  AOI22X1 U4011 ( .A(\data_in<13> ), .B(n1068), .C(\data_in<5> ), .D(n1069), 
        .Y(n606) );
  AOI22X1 U4012 ( .A(\data_in<12> ), .B(n1068), .C(\data_in<4> ), .D(n1069), 
        .Y(n605) );
  AOI22X1 U4013 ( .A(\data_in<11> ), .B(n1068), .C(\data_in<3> ), .D(n1069), 
        .Y(n604) );
  AOI22X1 U4014 ( .A(\data_in<10> ), .B(n1068), .C(\data_in<2> ), .D(n1069), 
        .Y(n603) );
  AOI22X1 U4015 ( .A(\data_in<9> ), .B(n1068), .C(\data_in<1> ), .D(n1069), 
        .Y(n602) );
  AOI22X1 U4016 ( .A(\data_in<8> ), .B(n1068), .C(\data_in<0> ), .D(n1069), 
        .Y(n599) );
  OAI21X1 U4017 ( .A(n1480), .B(n4793), .C(n933), .Y(n2966) );
  OAI21X1 U4018 ( .A(n2601), .B(n4806), .C(n935), .Y(n2965) );
  OAI21X1 U4019 ( .A(n1485), .B(n4777), .C(n937), .Y(n2968) );
  OAI21X1 U4020 ( .A(n2591), .B(n4782), .C(n939), .Y(n2967) );
  OAI21X1 U4021 ( .A(n4103), .B(n4738), .C(n941), .Y(n2970) );
  OAI21X1 U4022 ( .A(n4053), .B(n4754), .C(n943), .Y(n2969) );
  OAI21X1 U4023 ( .A(n4202), .B(n4706), .C(n945), .Y(n2972) );
  OAI21X1 U4024 ( .A(n4153), .B(n4722), .C(n947), .Y(n2971) );
  OAI21X1 U4025 ( .A(n411), .B(n4913), .C(n949), .Y(n2974) );
  OAI21X1 U4026 ( .A(n3448), .B(n4929), .C(n951), .Y(n2973) );
  OAI21X1 U4027 ( .A(n3572), .B(n4889), .C(n953), .Y(n2976) );
  OAI21X1 U4028 ( .A(n3547), .B(n4897), .C(n955), .Y(n2975) );
  OAI21X1 U4029 ( .A(n3696), .B(n4851), .C(n957), .Y(n2978) );
  OAI21X1 U4030 ( .A(n3646), .B(n4866), .C(n959), .Y(n2977) );
  OAI21X1 U4031 ( .A(n1518), .B(n4821), .C(n961), .Y(n2980) );
  OAI21X1 U4032 ( .A(n3746), .B(n4835), .C(n963), .Y(n2979) );
  OAI21X1 U4033 ( .A(n1480), .B(n4792), .C(n965), .Y(n2982) );
  OAI21X1 U4034 ( .A(n2601), .B(n4805), .C(n967), .Y(n2981) );
  OAI21X1 U4035 ( .A(n1485), .B(n4776), .C(n969), .Y(n2984) );
  OAI21X1 U4036 ( .A(n2591), .B(n4781), .C(n971), .Y(n2983) );
  OAI21X1 U4037 ( .A(n4103), .B(n4737), .C(n973), .Y(n2986) );
  OAI21X1 U4038 ( .A(n4053), .B(n4753), .C(n975), .Y(n2985) );
  OAI21X1 U4039 ( .A(n4202), .B(n4705), .C(n977), .Y(n2988) );
  OAI21X1 U4040 ( .A(n4153), .B(n4721), .C(n979), .Y(n2987) );
  OAI21X1 U4041 ( .A(n411), .B(n4912), .C(n981), .Y(n2990) );
  OAI21X1 U4042 ( .A(n3448), .B(n4928), .C(n983), .Y(n2989) );
  OAI21X1 U4043 ( .A(n3572), .B(n4888), .C(n985), .Y(n2992) );
  OAI21X1 U4044 ( .A(n3547), .B(n4896), .C(n987), .Y(n2991) );
  OAI21X1 U4045 ( .A(n3696), .B(n4850), .C(n989), .Y(n2994) );
  OAI21X1 U4046 ( .A(n3646), .B(n556), .C(n991), .Y(n2993) );
  OAI21X1 U4047 ( .A(n1518), .B(n4820), .C(n993), .Y(n2996) );
  OAI21X1 U4048 ( .A(n3746), .B(n4834), .C(n995), .Y(n2995) );
  OAI21X1 U4049 ( .A(n1480), .B(n4791), .C(n997), .Y(n2998) );
  OAI21X1 U4050 ( .A(n2601), .B(n4804), .C(n999), .Y(n2997) );
  OAI21X1 U4051 ( .A(n1485), .B(n4775), .C(n1001), .Y(n3000) );
  OAI21X1 U4052 ( .A(n2591), .B(n4780), .C(n1003), .Y(n2999) );
  OAI21X1 U4053 ( .A(n4103), .B(n4736), .C(n1005), .Y(n3002) );
  OAI21X1 U4054 ( .A(n4053), .B(n4752), .C(n1007), .Y(n3001) );
  OAI21X1 U4055 ( .A(n4202), .B(n4704), .C(n1009), .Y(n3004) );
  OAI21X1 U4056 ( .A(n4153), .B(n4720), .C(n1011), .Y(n3003) );
  OAI21X1 U4057 ( .A(n411), .B(n4911), .C(n1013), .Y(n3006) );
  OAI21X1 U4058 ( .A(n3448), .B(n4927), .C(n1015), .Y(n3005) );
  OAI21X1 U4059 ( .A(n3572), .B(n4887), .C(n1017), .Y(n3008) );
  OAI21X1 U4060 ( .A(n3547), .B(n4895), .C(n1019), .Y(n3007) );
  OAI21X1 U4061 ( .A(n3696), .B(n4849), .C(n1021), .Y(n3010) );
  OAI21X1 U4062 ( .A(n3646), .B(n4865), .C(n1023), .Y(n3009) );
  OAI21X1 U4063 ( .A(n1518), .B(n4819), .C(n1025), .Y(n3012) );
  OAI21X1 U4064 ( .A(n3746), .B(n4833), .C(n1027), .Y(n3011) );
  AOI22X1 U4065 ( .A(\data_in<8> ), .B(n1070), .C(n3015), .D(n1166), .Y(n3016)
         );
  OAI21X1 U4066 ( .A(n1305), .B(n3017), .C(n3016), .Y(n1824) );
  AOI22X1 U4067 ( .A(\data_in<9> ), .B(n1070), .C(n3018), .D(n1166), .Y(n3019)
         );
  OAI21X1 U4068 ( .A(n1305), .B(n3020), .C(n3019), .Y(n1825) );
  AOI22X1 U4069 ( .A(\data_in<10> ), .B(n1070), .C(n3021), .D(n1166), .Y(n3022) );
  OAI21X1 U4070 ( .A(n1305), .B(n3023), .C(n3022), .Y(n1826) );
  AOI22X1 U4071 ( .A(\data_in<11> ), .B(n1070), .C(n3024), .D(n1166), .Y(n3025) );
  OAI21X1 U4072 ( .A(n1305), .B(n3026), .C(n3025), .Y(n1827) );
  AOI22X1 U4073 ( .A(\data_in<12> ), .B(n1070), .C(n3027), .D(n1166), .Y(n3028) );
  OAI21X1 U4074 ( .A(n1305), .B(n3029), .C(n3028), .Y(n1828) );
  AOI22X1 U4075 ( .A(\data_in<13> ), .B(n1070), .C(n3030), .D(n1166), .Y(n3031) );
  OAI21X1 U4076 ( .A(n1305), .B(n3032), .C(n3031), .Y(n1829) );
  AOI22X1 U4077 ( .A(\data_in<14> ), .B(n1070), .C(n3033), .D(n1166), .Y(n3034) );
  OAI21X1 U4078 ( .A(n1305), .B(n3035), .C(n3034), .Y(n1830) );
  AOI22X1 U4079 ( .A(\data_in<15> ), .B(n1070), .C(n3036), .D(n1166), .Y(n3037) );
  OAI21X1 U4080 ( .A(n1305), .B(n3038), .C(n3037), .Y(n1831) );
  AOI22X1 U4081 ( .A(\data_in<8> ), .B(n1071), .C(n3040), .D(n1168), .Y(n3041)
         );
  OAI21X1 U4082 ( .A(n1307), .B(n3042), .C(n3041), .Y(n1832) );
  AOI22X1 U4083 ( .A(\data_in<9> ), .B(n1071), .C(n3043), .D(n1168), .Y(n3044)
         );
  OAI21X1 U4084 ( .A(n1307), .B(n3045), .C(n3044), .Y(n1833) );
  AOI22X1 U4085 ( .A(\data_in<10> ), .B(n1071), .C(n3046), .D(n1168), .Y(n3047) );
  OAI21X1 U4086 ( .A(n1307), .B(n3048), .C(n3047), .Y(n1834) );
  AOI22X1 U4087 ( .A(\data_in<11> ), .B(n1071), .C(n3049), .D(n1168), .Y(n3050) );
  OAI21X1 U4088 ( .A(n1307), .B(n3051), .C(n3050), .Y(n1835) );
  AOI22X1 U4089 ( .A(\data_in<12> ), .B(n1071), .C(n3052), .D(n1168), .Y(n3053) );
  OAI21X1 U4090 ( .A(n1307), .B(n3054), .C(n3053), .Y(n1836) );
  AOI22X1 U4091 ( .A(\data_in<13> ), .B(n1071), .C(n3055), .D(n1168), .Y(n3056) );
  OAI21X1 U4092 ( .A(n1307), .B(n3057), .C(n3056), .Y(n1837) );
  AOI22X1 U4093 ( .A(\data_in<14> ), .B(n1071), .C(n3058), .D(n1168), .Y(n3059) );
  OAI21X1 U4094 ( .A(n1307), .B(n3060), .C(n3059), .Y(n1838) );
  AOI22X1 U4095 ( .A(\data_in<15> ), .B(n1071), .C(n3061), .D(n1168), .Y(n3062) );
  OAI21X1 U4096 ( .A(n1307), .B(n3063), .C(n3062), .Y(n1839) );
  AOI22X1 U4097 ( .A(\data_in<8> ), .B(n1072), .C(n3066), .D(n1170), .Y(n3067)
         );
  OAI21X1 U4098 ( .A(n1309), .B(n3068), .C(n3067), .Y(n1840) );
  AOI22X1 U4099 ( .A(\data_in<9> ), .B(n1072), .C(n3069), .D(n1170), .Y(n3070)
         );
  OAI21X1 U4100 ( .A(n1309), .B(n3071), .C(n3070), .Y(n1841) );
  AOI22X1 U4101 ( .A(\data_in<10> ), .B(n1072), .C(n3072), .D(n1170), .Y(n3073) );
  OAI21X1 U4102 ( .A(n1309), .B(n3074), .C(n3073), .Y(n1842) );
  AOI22X1 U4103 ( .A(\data_in<11> ), .B(n1072), .C(n3075), .D(n1170), .Y(n3076) );
  OAI21X1 U4104 ( .A(n1309), .B(n3077), .C(n3076), .Y(n1843) );
  AOI22X1 U4105 ( .A(\data_in<12> ), .B(n1072), .C(n3078), .D(n1170), .Y(n3079) );
  OAI21X1 U4106 ( .A(n1309), .B(n3080), .C(n3079), .Y(n1844) );
  AOI22X1 U4107 ( .A(\data_in<13> ), .B(n1072), .C(n3081), .D(n1170), .Y(n3082) );
  OAI21X1 U4108 ( .A(n1309), .B(n3083), .C(n3082), .Y(n1845) );
  AOI22X1 U4109 ( .A(\data_in<14> ), .B(n1072), .C(n3084), .D(n1170), .Y(n3085) );
  OAI21X1 U4110 ( .A(n1309), .B(n3086), .C(n3085), .Y(n1846) );
  AOI22X1 U4111 ( .A(\data_in<15> ), .B(n1072), .C(n3087), .D(n1170), .Y(n3088) );
  OAI21X1 U4112 ( .A(n1309), .B(n3089), .C(n3088), .Y(n1847) );
  AOI22X1 U4113 ( .A(\data_in<8> ), .B(n1073), .C(n3092), .D(n1172), .Y(n3093)
         );
  OAI21X1 U4114 ( .A(n1311), .B(n3094), .C(n3093), .Y(n1848) );
  AOI22X1 U4115 ( .A(\data_in<9> ), .B(n1073), .C(n3095), .D(n1172), .Y(n3096)
         );
  OAI21X1 U4116 ( .A(n1311), .B(n3097), .C(n3096), .Y(n1849) );
  AOI22X1 U4117 ( .A(\data_in<10> ), .B(n1073), .C(n3098), .D(n1172), .Y(n3099) );
  OAI21X1 U4118 ( .A(n1311), .B(n3100), .C(n3099), .Y(n1850) );
  AOI22X1 U4119 ( .A(\data_in<11> ), .B(n1073), .C(n3101), .D(n1172), .Y(n3102) );
  OAI21X1 U4120 ( .A(n1311), .B(n3103), .C(n3102), .Y(n1851) );
  AOI22X1 U4121 ( .A(\data_in<12> ), .B(n1073), .C(n3104), .D(n1172), .Y(n3105) );
  OAI21X1 U4122 ( .A(n1311), .B(n3106), .C(n3105), .Y(n1852) );
  AOI22X1 U4123 ( .A(\data_in<13> ), .B(n1073), .C(n3107), .D(n1172), .Y(n3108) );
  OAI21X1 U4124 ( .A(n1311), .B(n3109), .C(n3108), .Y(n1853) );
  AOI22X1 U4125 ( .A(\data_in<14> ), .B(n1073), .C(n3110), .D(n1172), .Y(n3111) );
  OAI21X1 U4126 ( .A(n1311), .B(n3112), .C(n3111), .Y(n1854) );
  AOI22X1 U4127 ( .A(\data_in<15> ), .B(n1073), .C(n3113), .D(n1172), .Y(n3114) );
  OAI21X1 U4128 ( .A(n1311), .B(n3115), .C(n3114), .Y(n1855) );
  AOI22X1 U4129 ( .A(\data_in<8> ), .B(n1074), .C(n3117), .D(n1174), .Y(n3118)
         );
  OAI21X1 U4130 ( .A(n1313), .B(n3119), .C(n3118), .Y(n1856) );
  AOI22X1 U4131 ( .A(\data_in<9> ), .B(n1074), .C(n3120), .D(n1174), .Y(n3121)
         );
  OAI21X1 U4132 ( .A(n1313), .B(n3122), .C(n3121), .Y(n1857) );
  AOI22X1 U4133 ( .A(\data_in<10> ), .B(n1074), .C(n3123), .D(n1174), .Y(n3124) );
  OAI21X1 U4134 ( .A(n1313), .B(n3125), .C(n3124), .Y(n1858) );
  AOI22X1 U4135 ( .A(\data_in<11> ), .B(n1074), .C(n3126), .D(n1174), .Y(n3127) );
  OAI21X1 U4136 ( .A(n1313), .B(n3128), .C(n3127), .Y(n1859) );
  AOI22X1 U4137 ( .A(\data_in<12> ), .B(n1074), .C(n3129), .D(n1174), .Y(n3130) );
  OAI21X1 U4138 ( .A(n1313), .B(n3131), .C(n3130), .Y(n1860) );
  AOI22X1 U4139 ( .A(\data_in<13> ), .B(n1074), .C(n536), .D(n1174), .Y(n3132)
         );
  OAI21X1 U4140 ( .A(n1313), .B(n3133), .C(n3132), .Y(n1861) );
  AOI22X1 U4141 ( .A(\data_in<14> ), .B(n1074), .C(n3134), .D(n1174), .Y(n3135) );
  OAI21X1 U4142 ( .A(n1313), .B(n3136), .C(n3135), .Y(n1862) );
  AOI22X1 U4143 ( .A(\data_in<15> ), .B(n1074), .C(n3137), .D(n1174), .Y(n3138) );
  OAI21X1 U4144 ( .A(n1313), .B(n3139), .C(n3138), .Y(n1863) );
  AOI22X1 U4145 ( .A(\data_in<8> ), .B(n1075), .C(n3142), .D(n1176), .Y(n3143)
         );
  OAI21X1 U4146 ( .A(n1315), .B(n3144), .C(n3143), .Y(n1864) );
  AOI22X1 U4147 ( .A(\data_in<9> ), .B(n1075), .C(n3145), .D(n1176), .Y(n3146)
         );
  OAI21X1 U4148 ( .A(n1315), .B(n3147), .C(n3146), .Y(n1865) );
  AOI22X1 U4149 ( .A(\data_in<10> ), .B(n1075), .C(n3148), .D(n1176), .Y(n3149) );
  OAI21X1 U4150 ( .A(n1315), .B(n3150), .C(n3149), .Y(n1866) );
  AOI22X1 U4151 ( .A(\data_in<11> ), .B(n1075), .C(n3151), .D(n1176), .Y(n3152) );
  OAI21X1 U4152 ( .A(n1315), .B(n3153), .C(n3152), .Y(n1867) );
  AOI22X1 U4153 ( .A(\data_in<12> ), .B(n1075), .C(n3154), .D(n1176), .Y(n3155) );
  OAI21X1 U4154 ( .A(n1315), .B(n3156), .C(n3155), .Y(n1868) );
  AOI22X1 U4155 ( .A(\data_in<13> ), .B(n1075), .C(n3157), .D(n1176), .Y(n3158) );
  OAI21X1 U4156 ( .A(n1315), .B(n3159), .C(n3158), .Y(n1869) );
  AOI22X1 U4157 ( .A(\data_in<14> ), .B(n1075), .C(n3160), .D(n1176), .Y(n3161) );
  OAI21X1 U4158 ( .A(n1315), .B(n3162), .C(n3161), .Y(n1870) );
  AOI22X1 U4159 ( .A(\data_in<15> ), .B(n1075), .C(n3163), .D(n1176), .Y(n3164) );
  OAI21X1 U4160 ( .A(n1315), .B(n3165), .C(n3164), .Y(n1871) );
  AOI22X1 U4161 ( .A(\data_in<8> ), .B(n1076), .C(n3168), .D(n1178), .Y(n3169)
         );
  OAI21X1 U4162 ( .A(n1317), .B(n3170), .C(n3169), .Y(n1872) );
  AOI22X1 U4163 ( .A(\data_in<9> ), .B(n1076), .C(n3171), .D(n1178), .Y(n3172)
         );
  OAI21X1 U4164 ( .A(n1317), .B(n3173), .C(n3172), .Y(n1873) );
  AOI22X1 U4165 ( .A(\data_in<10> ), .B(n1076), .C(n3174), .D(n1178), .Y(n3175) );
  OAI21X1 U4166 ( .A(n1317), .B(n3176), .C(n3175), .Y(n1874) );
  AOI22X1 U4167 ( .A(\data_in<11> ), .B(n1076), .C(n3177), .D(n1178), .Y(n3178) );
  OAI21X1 U4168 ( .A(n1317), .B(n3179), .C(n3178), .Y(n1875) );
  AOI22X1 U4169 ( .A(\data_in<12> ), .B(n1076), .C(n3180), .D(n1178), .Y(n3181) );
  OAI21X1 U4170 ( .A(n1317), .B(n3182), .C(n3181), .Y(n1876) );
  AOI22X1 U4171 ( .A(\data_in<13> ), .B(n1076), .C(n3183), .D(n1178), .Y(n3184) );
  OAI21X1 U4172 ( .A(n1317), .B(n3185), .C(n3184), .Y(n1877) );
  AOI22X1 U4173 ( .A(\data_in<14> ), .B(n1076), .C(n3186), .D(n1178), .Y(n3187) );
  OAI21X1 U4174 ( .A(n1317), .B(n3188), .C(n3187), .Y(n1878) );
  AOI22X1 U4175 ( .A(\data_in<15> ), .B(n1076), .C(n3189), .D(n1178), .Y(n3190) );
  OAI21X1 U4176 ( .A(n1317), .B(n3191), .C(n3190), .Y(n1879) );
  OAI21X1 U4177 ( .A(n1487), .B(n1477), .C(n1294), .Y(n3214) );
  AOI22X1 U4178 ( .A(\data_in<8> ), .B(n1077), .C(n3193), .D(n3214), .Y(n3194)
         );
  OAI21X1 U4179 ( .A(n1319), .B(n3195), .C(n3194), .Y(n1880) );
  AOI22X1 U4180 ( .A(\data_in<9> ), .B(n1077), .C(n3196), .D(n3214), .Y(n3197)
         );
  OAI21X1 U4181 ( .A(n1319), .B(n3198), .C(n3197), .Y(n1881) );
  AOI22X1 U4182 ( .A(\data_in<10> ), .B(n1077), .C(n3199), .D(n3214), .Y(n3200) );
  OAI21X1 U4183 ( .A(n1319), .B(n3201), .C(n3200), .Y(n1882) );
  AOI22X1 U4184 ( .A(\data_in<11> ), .B(n1077), .C(n3202), .D(n3214), .Y(n3203) );
  OAI21X1 U4185 ( .A(n1319), .B(n3204), .C(n3203), .Y(n1883) );
  AOI22X1 U4186 ( .A(\data_in<12> ), .B(n1077), .C(n3205), .D(n3214), .Y(n3206) );
  OAI21X1 U4187 ( .A(n1319), .B(n3207), .C(n3206), .Y(n1884) );
  AOI22X1 U4188 ( .A(\data_in<13> ), .B(n1077), .C(n3208), .D(n3214), .Y(n3209) );
  OAI21X1 U4189 ( .A(n1319), .B(n3210), .C(n3209), .Y(n1885) );
  AOI22X1 U4190 ( .A(\data_in<14> ), .B(n1077), .C(n3211), .D(n3214), .Y(n3212) );
  OAI21X1 U4191 ( .A(n1319), .B(n3213), .C(n3212), .Y(n1886) );
  AOI22X1 U4192 ( .A(\data_in<15> ), .B(n1077), .C(n3215), .D(n3214), .Y(n3216) );
  OAI21X1 U4193 ( .A(n1319), .B(n3217), .C(n3216), .Y(n1887) );
  AOI22X1 U4194 ( .A(\data_in<8> ), .B(n1078), .C(n3218), .D(n1180), .Y(n3219)
         );
  OAI21X1 U4195 ( .A(n1321), .B(n3220), .C(n3219), .Y(n1888) );
  AOI22X1 U4196 ( .A(\data_in<9> ), .B(n1078), .C(n3221), .D(n1180), .Y(n3222)
         );
  OAI21X1 U4197 ( .A(n1321), .B(n3223), .C(n3222), .Y(n1889) );
  AOI22X1 U4198 ( .A(\data_in<10> ), .B(n1078), .C(n3224), .D(n1180), .Y(n3225) );
  OAI21X1 U4199 ( .A(n1321), .B(n3226), .C(n3225), .Y(n1890) );
  AOI22X1 U4200 ( .A(\data_in<11> ), .B(n1078), .C(n3227), .D(n1180), .Y(n3228) );
  OAI21X1 U4201 ( .A(n1321), .B(n3229), .C(n3228), .Y(n1891) );
  AOI22X1 U4202 ( .A(\data_in<12> ), .B(n1078), .C(n3230), .D(n1180), .Y(n3231) );
  OAI21X1 U4203 ( .A(n1321), .B(n3232), .C(n3231), .Y(n1892) );
  AOI22X1 U4204 ( .A(\data_in<13> ), .B(n1078), .C(n3233), .D(n1180), .Y(n3234) );
  OAI21X1 U4205 ( .A(n1321), .B(n3235), .C(n3234), .Y(n1893) );
  AOI22X1 U4206 ( .A(\data_in<14> ), .B(n1078), .C(n3236), .D(n1180), .Y(n3237) );
  OAI21X1 U4207 ( .A(n1321), .B(n3238), .C(n3237), .Y(n1894) );
  AOI22X1 U4208 ( .A(\data_in<15> ), .B(n1078), .C(n3239), .D(n1180), .Y(n3240) );
  OAI21X1 U4209 ( .A(n1321), .B(n3241), .C(n3240), .Y(n1895) );
  AOI22X1 U4210 ( .A(\data_in<8> ), .B(n1079), .C(n3243), .D(n1182), .Y(n3244)
         );
  OAI21X1 U4211 ( .A(n1323), .B(n3245), .C(n3244), .Y(n1896) );
  AOI22X1 U4212 ( .A(\data_in<9> ), .B(n1079), .C(n3246), .D(n1182), .Y(n3247)
         );
  OAI21X1 U4213 ( .A(n1323), .B(n3248), .C(n3247), .Y(n1897) );
  AOI22X1 U4214 ( .A(\data_in<10> ), .B(n1079), .C(n3249), .D(n1182), .Y(n3250) );
  OAI21X1 U4215 ( .A(n1323), .B(n3251), .C(n3250), .Y(n1898) );
  AOI22X1 U4216 ( .A(\data_in<11> ), .B(n1079), .C(n3252), .D(n1182), .Y(n3253) );
  OAI21X1 U4217 ( .A(n1323), .B(n3254), .C(n3253), .Y(n1899) );
  AOI22X1 U4218 ( .A(\data_in<12> ), .B(n1079), .C(n3255), .D(n1182), .Y(n3256) );
  OAI21X1 U4219 ( .A(n1323), .B(n3257), .C(n3256), .Y(n1900) );
  AOI22X1 U4220 ( .A(\data_in<13> ), .B(n1079), .C(n3258), .D(n1182), .Y(n3259) );
  OAI21X1 U4221 ( .A(n1323), .B(n3260), .C(n3259), .Y(n1901) );
  AOI22X1 U4222 ( .A(\data_in<14> ), .B(n1079), .C(n3261), .D(n1182), .Y(n3262) );
  OAI21X1 U4223 ( .A(n1323), .B(n3263), .C(n3262), .Y(n1902) );
  AOI22X1 U4224 ( .A(\data_in<15> ), .B(n1079), .C(n3264), .D(n1182), .Y(n3265) );
  OAI21X1 U4225 ( .A(n1323), .B(n3266), .C(n3265), .Y(n1903) );
  OAI21X1 U4226 ( .A(n482), .B(n506), .C(n1294), .Y(n3290) );
  AOI22X1 U4227 ( .A(\data_in<8> ), .B(n1080), .C(n3269), .D(n3290), .Y(n3270)
         );
  OAI21X1 U4228 ( .A(n1325), .B(n3271), .C(n3270), .Y(n1904) );
  AOI22X1 U4229 ( .A(\data_in<9> ), .B(n1080), .C(n3272), .D(n3290), .Y(n3273)
         );
  OAI21X1 U4230 ( .A(n1325), .B(n3274), .C(n3273), .Y(n1905) );
  AOI22X1 U4231 ( .A(\data_in<10> ), .B(n1080), .C(n3275), .D(n3290), .Y(n3276) );
  OAI21X1 U4232 ( .A(n1325), .B(n3277), .C(n3276), .Y(n1906) );
  AOI22X1 U4233 ( .A(\data_in<11> ), .B(n1080), .C(n3278), .D(n3290), .Y(n3279) );
  OAI21X1 U4234 ( .A(n1325), .B(n3280), .C(n3279), .Y(n1907) );
  AOI22X1 U4235 ( .A(\data_in<12> ), .B(n1080), .C(n3281), .D(n3290), .Y(n3282) );
  OAI21X1 U4236 ( .A(n1325), .B(n3283), .C(n3282), .Y(n1908) );
  AOI22X1 U4237 ( .A(\data_in<13> ), .B(n1080), .C(n3284), .D(n3290), .Y(n3285) );
  OAI21X1 U4238 ( .A(n1325), .B(n3286), .C(n3285), .Y(n1909) );
  AOI22X1 U4239 ( .A(\data_in<14> ), .B(n1080), .C(n3287), .D(n3290), .Y(n3288) );
  OAI21X1 U4240 ( .A(n1325), .B(n3289), .C(n3288), .Y(n1910) );
  AOI22X1 U4241 ( .A(\data_in<15> ), .B(n1080), .C(n3291), .D(n3290), .Y(n3292) );
  OAI21X1 U4242 ( .A(n1325), .B(n3293), .C(n3292), .Y(n1911) );
  OAI21X1 U4243 ( .A(n1491), .B(n506), .C(n1294), .Y(n3316) );
  AOI22X1 U4244 ( .A(\data_in<8> ), .B(n1081), .C(n3295), .D(n3316), .Y(n3296)
         );
  OAI21X1 U4245 ( .A(n1327), .B(n3297), .C(n3296), .Y(n1912) );
  AOI22X1 U4246 ( .A(\data_in<9> ), .B(n1081), .C(n3298), .D(n3316), .Y(n3299)
         );
  OAI21X1 U4247 ( .A(n1327), .B(n3300), .C(n3299), .Y(n1913) );
  AOI22X1 U4248 ( .A(\data_in<10> ), .B(n1081), .C(n3301), .D(n3316), .Y(n3302) );
  OAI21X1 U4249 ( .A(n1327), .B(n3303), .C(n3302), .Y(n1914) );
  AOI22X1 U4250 ( .A(\data_in<11> ), .B(n1081), .C(n3304), .D(n3316), .Y(n3305) );
  OAI21X1 U4251 ( .A(n1327), .B(n3306), .C(n3305), .Y(n1915) );
  AOI22X1 U4252 ( .A(\data_in<12> ), .B(n1081), .C(n3307), .D(n3316), .Y(n3308) );
  OAI21X1 U4253 ( .A(n1327), .B(n3309), .C(n3308), .Y(n1916) );
  AOI22X1 U4254 ( .A(\data_in<13> ), .B(n1081), .C(n3310), .D(n3316), .Y(n3311) );
  OAI21X1 U4255 ( .A(n1327), .B(n3312), .C(n3311), .Y(n1917) );
  AOI22X1 U4256 ( .A(\data_in<14> ), .B(n1081), .C(n3313), .D(n3316), .Y(n3314) );
  OAI21X1 U4257 ( .A(n1327), .B(n3315), .C(n3314), .Y(n1918) );
  AOI22X1 U4258 ( .A(\data_in<15> ), .B(n1081), .C(n3317), .D(n3316), .Y(n3318) );
  OAI21X1 U4259 ( .A(n1327), .B(n3319), .C(n3318), .Y(n1919) );
  OAI21X1 U4260 ( .A(n1491), .B(n436), .C(n1294), .Y(n3344) );
  AOI22X1 U4261 ( .A(\data_in<8> ), .B(n1082), .C(n3323), .D(n3344), .Y(n3324)
         );
  OAI21X1 U4262 ( .A(n1329), .B(n3325), .C(n3324), .Y(n1920) );
  AOI22X1 U4263 ( .A(\data_in<9> ), .B(n1082), .C(n3326), .D(n3344), .Y(n3327)
         );
  OAI21X1 U4264 ( .A(n1329), .B(n3328), .C(n3327), .Y(n1921) );
  AOI22X1 U4265 ( .A(\data_in<10> ), .B(n1082), .C(n3329), .D(n3344), .Y(n3330) );
  OAI21X1 U4266 ( .A(n1329), .B(n3331), .C(n3330), .Y(n1922) );
  AOI22X1 U4267 ( .A(\data_in<11> ), .B(n1082), .C(n3332), .D(n3344), .Y(n3333) );
  OAI21X1 U4268 ( .A(n1329), .B(n3334), .C(n3333), .Y(n1923) );
  AOI22X1 U4269 ( .A(\data_in<12> ), .B(n1082), .C(n3335), .D(n3344), .Y(n3336) );
  OAI21X1 U4270 ( .A(n1329), .B(n3337), .C(n3336), .Y(n1924) );
  AOI22X1 U4271 ( .A(\data_in<13> ), .B(n1082), .C(n3338), .D(n3344), .Y(n3339) );
  OAI21X1 U4272 ( .A(n1329), .B(n3340), .C(n3339), .Y(n1925) );
  AOI22X1 U4273 ( .A(\data_in<14> ), .B(n1082), .C(n3341), .D(n3344), .Y(n3342) );
  OAI21X1 U4274 ( .A(n1329), .B(n3343), .C(n3342), .Y(n1926) );
  AOI22X1 U4275 ( .A(\data_in<15> ), .B(n1082), .C(n3345), .D(n3344), .Y(n3346) );
  OAI21X1 U4276 ( .A(n1329), .B(n3347), .C(n3346), .Y(n1927) );
  OAI21X1 U4277 ( .A(n440), .B(n436), .C(n1294), .Y(n3370) );
  AOI22X1 U4278 ( .A(\data_in<8> ), .B(n1083), .C(n3349), .D(n3370), .Y(n3350)
         );
  OAI21X1 U4279 ( .A(n1331), .B(n3351), .C(n3350), .Y(n1928) );
  AOI22X1 U4280 ( .A(\data_in<9> ), .B(n1083), .C(n3352), .D(n3370), .Y(n3353)
         );
  OAI21X1 U4281 ( .A(n1331), .B(n3354), .C(n3353), .Y(n1929) );
  AOI22X1 U4282 ( .A(\data_in<10> ), .B(n1083), .C(n3355), .D(n3370), .Y(n3356) );
  OAI21X1 U4283 ( .A(n1331), .B(n3357), .C(n3356), .Y(n1930) );
  AOI22X1 U4284 ( .A(\data_in<11> ), .B(n1083), .C(n3358), .D(n3370), .Y(n3359) );
  OAI21X1 U4285 ( .A(n1331), .B(n3360), .C(n3359), .Y(n1931) );
  AOI22X1 U4286 ( .A(\data_in<12> ), .B(n1083), .C(n3361), .D(n3370), .Y(n3362) );
  OAI21X1 U4287 ( .A(n1331), .B(n3363), .C(n3362), .Y(n1932) );
  AOI22X1 U4288 ( .A(\data_in<13> ), .B(n1083), .C(n3364), .D(n3370), .Y(n3365) );
  OAI21X1 U4289 ( .A(n1331), .B(n3366), .C(n3365), .Y(n1933) );
  AOI22X1 U4290 ( .A(\data_in<14> ), .B(n1083), .C(n3367), .D(n3370), .Y(n3368) );
  OAI21X1 U4291 ( .A(n1331), .B(n3369), .C(n3368), .Y(n1934) );
  AOI22X1 U4292 ( .A(\data_in<15> ), .B(n1083), .C(n3371), .D(n3370), .Y(n3372) );
  OAI21X1 U4293 ( .A(n1331), .B(n3373), .C(n3372), .Y(n1935) );
  AOI22X1 U4294 ( .A(\data_in<8> ), .B(n1084), .C(n3374), .D(n1184), .Y(n3375)
         );
  OAI21X1 U4295 ( .A(n1333), .B(n3376), .C(n3375), .Y(n1936) );
  AOI22X1 U4296 ( .A(\data_in<9> ), .B(n1084), .C(n3377), .D(n1184), .Y(n3378)
         );
  OAI21X1 U4297 ( .A(n1333), .B(n3379), .C(n3378), .Y(n1937) );
  AOI22X1 U4298 ( .A(\data_in<10> ), .B(n1084), .C(n3380), .D(n1184), .Y(n3381) );
  OAI21X1 U4299 ( .A(n1333), .B(n3382), .C(n3381), .Y(n1938) );
  AOI22X1 U4300 ( .A(\data_in<11> ), .B(n1084), .C(n3383), .D(n1184), .Y(n3384) );
  OAI21X1 U4301 ( .A(n1333), .B(n3385), .C(n3384), .Y(n1939) );
  AOI22X1 U4302 ( .A(\data_in<12> ), .B(n1084), .C(n3386), .D(n1184), .Y(n3387) );
  OAI21X1 U4303 ( .A(n1333), .B(n3388), .C(n3387), .Y(n1940) );
  AOI22X1 U4304 ( .A(\data_in<13> ), .B(n1084), .C(n3389), .D(n1184), .Y(n3390) );
  OAI21X1 U4305 ( .A(n1333), .B(n3391), .C(n3390), .Y(n1941) );
  AOI22X1 U4306 ( .A(\data_in<14> ), .B(n1084), .C(n3392), .D(n1184), .Y(n3393) );
  OAI21X1 U4307 ( .A(n1333), .B(n3394), .C(n3393), .Y(n1942) );
  AOI22X1 U4308 ( .A(\data_in<15> ), .B(n1084), .C(n3395), .D(n1184), .Y(n3396) );
  OAI21X1 U4309 ( .A(n1333), .B(n3397), .C(n3396), .Y(n1943) );
  AOI22X1 U4310 ( .A(\data_in<8> ), .B(n1085), .C(n3399), .D(n1186), .Y(n3400)
         );
  OAI21X1 U4311 ( .A(n1335), .B(n3401), .C(n3400), .Y(n1944) );
  AOI22X1 U4312 ( .A(\data_in<9> ), .B(n1085), .C(n3402), .D(n1186), .Y(n3403)
         );
  OAI21X1 U4313 ( .A(n1335), .B(n3404), .C(n3403), .Y(n1945) );
  AOI22X1 U4314 ( .A(\data_in<10> ), .B(n1085), .C(n3405), .D(n1186), .Y(n3406) );
  OAI21X1 U4315 ( .A(n1335), .B(n3407), .C(n3406), .Y(n1946) );
  AOI22X1 U4316 ( .A(\data_in<11> ), .B(n1085), .C(n3408), .D(n1186), .Y(n3409) );
  OAI21X1 U4317 ( .A(n1335), .B(n3410), .C(n3409), .Y(n1947) );
  AOI22X1 U4318 ( .A(\data_in<12> ), .B(n1085), .C(n3411), .D(n1186), .Y(n3412) );
  OAI21X1 U4319 ( .A(n1335), .B(n3413), .C(n3412), .Y(n1948) );
  AOI22X1 U4320 ( .A(\data_in<13> ), .B(n1085), .C(n3414), .D(n1186), .Y(n3415) );
  OAI21X1 U4321 ( .A(n1335), .B(n3416), .C(n3415), .Y(n1949) );
  AOI22X1 U4322 ( .A(\data_in<14> ), .B(n1085), .C(n3417), .D(n1186), .Y(n3418) );
  OAI21X1 U4323 ( .A(n1335), .B(n3419), .C(n3418), .Y(n1950) );
  AOI22X1 U4324 ( .A(\data_in<15> ), .B(n1085), .C(n3420), .D(n1186), .Y(n3421) );
  OAI21X1 U4325 ( .A(n1335), .B(n3422), .C(n3421), .Y(n1951) );
  AOI22X1 U4326 ( .A(\data_in<8> ), .B(n1086), .C(n3424), .D(n1188), .Y(n3425)
         );
  OAI21X1 U4327 ( .A(n1337), .B(n3426), .C(n3425), .Y(n1952) );
  AOI22X1 U4328 ( .A(\data_in<9> ), .B(n1086), .C(n3427), .D(n1188), .Y(n3428)
         );
  OAI21X1 U4329 ( .A(n1337), .B(n3429), .C(n3428), .Y(n1953) );
  AOI22X1 U4330 ( .A(\data_in<10> ), .B(n1086), .C(n3430), .D(n1188), .Y(n3431) );
  OAI21X1 U4331 ( .A(n1337), .B(n3432), .C(n3431), .Y(n1954) );
  AOI22X1 U4332 ( .A(\data_in<11> ), .B(n1086), .C(n3433), .D(n1188), .Y(n3434) );
  OAI21X1 U4333 ( .A(n1337), .B(n3435), .C(n3434), .Y(n1955) );
  AOI22X1 U4334 ( .A(\data_in<12> ), .B(n1086), .C(n3436), .D(n1188), .Y(n3437) );
  OAI21X1 U4335 ( .A(n1337), .B(n3438), .C(n3437), .Y(n1956) );
  AOI22X1 U4336 ( .A(\data_in<13> ), .B(n1086), .C(n3439), .D(n1188), .Y(n3440) );
  OAI21X1 U4337 ( .A(n1337), .B(n3441), .C(n3440), .Y(n1957) );
  AOI22X1 U4338 ( .A(\data_in<14> ), .B(n1086), .C(n3442), .D(n1188), .Y(n3443) );
  OAI21X1 U4339 ( .A(n1337), .B(n3444), .C(n3443), .Y(n1958) );
  AOI22X1 U4340 ( .A(\data_in<15> ), .B(n1086), .C(n3445), .D(n1188), .Y(n3446) );
  OAI21X1 U4341 ( .A(n1337), .B(n3447), .C(n3446), .Y(n1959) );
  AOI22X1 U4342 ( .A(\data_in<8> ), .B(n1087), .C(n3449), .D(n1190), .Y(n3450)
         );
  OAI21X1 U4343 ( .A(n1339), .B(n3451), .C(n3450), .Y(n1960) );
  AOI22X1 U4344 ( .A(\data_in<9> ), .B(n1087), .C(n3452), .D(n1190), .Y(n3453)
         );
  OAI21X1 U4345 ( .A(n1339), .B(n3454), .C(n3453), .Y(n1961) );
  AOI22X1 U4346 ( .A(\data_in<10> ), .B(n1087), .C(n3455), .D(n1190), .Y(n3456) );
  OAI21X1 U4347 ( .A(n1339), .B(n3457), .C(n3456), .Y(n1962) );
  AOI22X1 U4348 ( .A(\data_in<11> ), .B(n1087), .C(n3458), .D(n1190), .Y(n3459) );
  OAI21X1 U4349 ( .A(n1339), .B(n3460), .C(n3459), .Y(n1963) );
  AOI22X1 U4350 ( .A(\data_in<12> ), .B(n1087), .C(n3461), .D(n1190), .Y(n3462) );
  OAI21X1 U4351 ( .A(n1339), .B(n3463), .C(n3462), .Y(n1964) );
  AOI22X1 U4352 ( .A(\data_in<13> ), .B(n1087), .C(n3464), .D(n1190), .Y(n3465) );
  OAI21X1 U4353 ( .A(n1339), .B(n3466), .C(n3465), .Y(n1965) );
  AOI22X1 U4354 ( .A(\data_in<14> ), .B(n1087), .C(n3467), .D(n1190), .Y(n3468) );
  OAI21X1 U4355 ( .A(n1339), .B(n3469), .C(n3468), .Y(n1966) );
  AOI22X1 U4356 ( .A(\data_in<15> ), .B(n1087), .C(n3470), .D(n1190), .Y(n3471) );
  OAI21X1 U4357 ( .A(n1339), .B(n3472), .C(n3471), .Y(n1967) );
  AOI22X1 U4358 ( .A(\data_in<8> ), .B(n1088), .C(n3474), .D(n1192), .Y(n3475)
         );
  OAI21X1 U4359 ( .A(n1341), .B(n3476), .C(n3475), .Y(n1968) );
  AOI22X1 U4360 ( .A(\data_in<9> ), .B(n1088), .C(n3477), .D(n1192), .Y(n3478)
         );
  OAI21X1 U4361 ( .A(n1341), .B(n3479), .C(n3478), .Y(n1969) );
  AOI22X1 U4362 ( .A(\data_in<10> ), .B(n1088), .C(n3480), .D(n1192), .Y(n3481) );
  OAI21X1 U4363 ( .A(n1341), .B(n3482), .C(n3481), .Y(n1970) );
  AOI22X1 U4364 ( .A(\data_in<11> ), .B(n1088), .C(n3483), .D(n1192), .Y(n3484) );
  OAI21X1 U4365 ( .A(n1341), .B(n3485), .C(n3484), .Y(n1971) );
  AOI22X1 U4366 ( .A(\data_in<12> ), .B(n1088), .C(n3486), .D(n1192), .Y(n3487) );
  OAI21X1 U4367 ( .A(n1341), .B(n3488), .C(n3487), .Y(n1972) );
  AOI22X1 U4368 ( .A(\data_in<13> ), .B(n1088), .C(n3489), .D(n1192), .Y(n3490) );
  OAI21X1 U4369 ( .A(n1341), .B(n3491), .C(n3490), .Y(n1973) );
  AOI22X1 U4370 ( .A(\data_in<14> ), .B(n1088), .C(n3492), .D(n1192), .Y(n3493) );
  OAI21X1 U4371 ( .A(n1341), .B(n3494), .C(n3493), .Y(n1974) );
  AOI22X1 U4372 ( .A(\data_in<15> ), .B(n1088), .C(n3495), .D(n1192), .Y(n3496) );
  OAI21X1 U4373 ( .A(n1341), .B(n3497), .C(n3496), .Y(n1975) );
  AOI22X1 U4374 ( .A(\data_in<8> ), .B(n1089), .C(n3498), .D(n1194), .Y(n3499)
         );
  OAI21X1 U4375 ( .A(n1343), .B(n3500), .C(n3499), .Y(n1976) );
  AOI22X1 U4376 ( .A(\data_in<9> ), .B(n1089), .C(n3501), .D(n1194), .Y(n3502)
         );
  OAI21X1 U4377 ( .A(n1343), .B(n3503), .C(n3502), .Y(n1977) );
  AOI22X1 U4378 ( .A(\data_in<10> ), .B(n1089), .C(n3504), .D(n1194), .Y(n3505) );
  OAI21X1 U4379 ( .A(n1343), .B(n3506), .C(n3505), .Y(n1978) );
  AOI22X1 U4380 ( .A(\data_in<11> ), .B(n1089), .C(n3507), .D(n1194), .Y(n3508) );
  OAI21X1 U4381 ( .A(n1343), .B(n3509), .C(n3508), .Y(n1979) );
  AOI22X1 U4382 ( .A(\data_in<12> ), .B(n1089), .C(n3510), .D(n1194), .Y(n3511) );
  OAI21X1 U4383 ( .A(n1343), .B(n3512), .C(n3511), .Y(n1980) );
  AOI22X1 U4384 ( .A(\data_in<13> ), .B(n1089), .C(n3513), .D(n1194), .Y(n3514) );
  OAI21X1 U4385 ( .A(n1343), .B(n3515), .C(n3514), .Y(n1981) );
  AOI22X1 U4386 ( .A(\data_in<14> ), .B(n1089), .C(n3516), .D(n1194), .Y(n3517) );
  OAI21X1 U4387 ( .A(n1343), .B(n3518), .C(n3517), .Y(n1982) );
  AOI22X1 U4388 ( .A(\data_in<15> ), .B(n1089), .C(n3519), .D(n1194), .Y(n3520) );
  OAI21X1 U4389 ( .A(n1343), .B(n3521), .C(n3520), .Y(n1983) );
  AOI22X1 U4390 ( .A(\data_in<8> ), .B(n1090), .C(n3523), .D(n1196), .Y(n3524)
         );
  OAI21X1 U4391 ( .A(n1345), .B(n3525), .C(n3524), .Y(n1984) );
  AOI22X1 U4392 ( .A(\data_in<9> ), .B(n1090), .C(n3526), .D(n1196), .Y(n3527)
         );
  OAI21X1 U4393 ( .A(n1345), .B(n3528), .C(n3527), .Y(n1985) );
  AOI22X1 U4394 ( .A(\data_in<10> ), .B(n1090), .C(n3529), .D(n1196), .Y(n3530) );
  OAI21X1 U4395 ( .A(n1345), .B(n3531), .C(n3530), .Y(n1986) );
  AOI22X1 U4396 ( .A(\data_in<11> ), .B(n1090), .C(n3532), .D(n1196), .Y(n3533) );
  OAI21X1 U4397 ( .A(n1345), .B(n3534), .C(n3533), .Y(n1987) );
  AOI22X1 U4398 ( .A(\data_in<12> ), .B(n1090), .C(n3535), .D(n1196), .Y(n3536) );
  OAI21X1 U4399 ( .A(n1345), .B(n3537), .C(n3536), .Y(n1988) );
  AOI22X1 U4400 ( .A(\data_in<13> ), .B(n1090), .C(n3538), .D(n1196), .Y(n3539) );
  OAI21X1 U4401 ( .A(n1345), .B(n3540), .C(n3539), .Y(n1989) );
  AOI22X1 U4402 ( .A(\data_in<14> ), .B(n1090), .C(n3541), .D(n1196), .Y(n3542) );
  OAI21X1 U4403 ( .A(n1345), .B(n3543), .C(n3542), .Y(n1990) );
  AOI22X1 U4404 ( .A(\data_in<15> ), .B(n1090), .C(n3544), .D(n1196), .Y(n3545) );
  OAI21X1 U4405 ( .A(n1345), .B(n3546), .C(n3545), .Y(n1991) );
  AOI22X1 U4406 ( .A(\data_in<8> ), .B(n1091), .C(n3548), .D(n1198), .Y(n3549)
         );
  OAI21X1 U4407 ( .A(n1347), .B(n3550), .C(n3549), .Y(n1992) );
  AOI22X1 U4408 ( .A(\data_in<9> ), .B(n1091), .C(n3551), .D(n1198), .Y(n3552)
         );
  OAI21X1 U4409 ( .A(n1347), .B(n3553), .C(n3552), .Y(n1993) );
  AOI22X1 U4410 ( .A(\data_in<10> ), .B(n1091), .C(n3554), .D(n1198), .Y(n3555) );
  OAI21X1 U4411 ( .A(n1347), .B(n3556), .C(n3555), .Y(n1994) );
  AOI22X1 U4412 ( .A(\data_in<11> ), .B(n1091), .C(n3557), .D(n1198), .Y(n3558) );
  OAI21X1 U4413 ( .A(n1347), .B(n3559), .C(n3558), .Y(n1995) );
  AOI22X1 U4414 ( .A(\data_in<12> ), .B(n1091), .C(n3560), .D(n1198), .Y(n3561) );
  OAI21X1 U4415 ( .A(n1347), .B(n3562), .C(n3561), .Y(n1996) );
  AOI22X1 U4416 ( .A(\data_in<13> ), .B(n1091), .C(n3563), .D(n1198), .Y(n3564) );
  OAI21X1 U4417 ( .A(n1347), .B(n3565), .C(n3564), .Y(n1997) );
  AOI22X1 U4418 ( .A(\data_in<14> ), .B(n1091), .C(n3566), .D(n1198), .Y(n3567) );
  OAI21X1 U4419 ( .A(n1347), .B(n3568), .C(n3567), .Y(n1998) );
  AOI22X1 U4420 ( .A(\data_in<15> ), .B(n1091), .C(n3569), .D(n1198), .Y(n3570) );
  OAI21X1 U4421 ( .A(n1347), .B(n3571), .C(n3570), .Y(n1999) );
  AOI22X1 U4422 ( .A(\data_in<8> ), .B(n1092), .C(n3573), .D(n1200), .Y(n3574)
         );
  OAI21X1 U4423 ( .A(n1349), .B(n3575), .C(n3574), .Y(n2000) );
  AOI22X1 U4424 ( .A(\data_in<9> ), .B(n1092), .C(n3576), .D(n1200), .Y(n3577)
         );
  OAI21X1 U4425 ( .A(n1349), .B(n3578), .C(n3577), .Y(n2001) );
  AOI22X1 U4426 ( .A(\data_in<10> ), .B(n1092), .C(n3579), .D(n1200), .Y(n3580) );
  OAI21X1 U4427 ( .A(n1349), .B(n3581), .C(n3580), .Y(n2002) );
  AOI22X1 U4428 ( .A(\data_in<11> ), .B(n1092), .C(n3582), .D(n1200), .Y(n3583) );
  OAI21X1 U4429 ( .A(n1349), .B(n3584), .C(n3583), .Y(n2003) );
  AOI22X1 U4430 ( .A(\data_in<12> ), .B(n1092), .C(n3585), .D(n1200), .Y(n3586) );
  OAI21X1 U4431 ( .A(n1349), .B(n3587), .C(n3586), .Y(n2004) );
  AOI22X1 U4432 ( .A(\data_in<13> ), .B(n1092), .C(n3588), .D(n1200), .Y(n3589) );
  OAI21X1 U4433 ( .A(n1349), .B(n3590), .C(n3589), .Y(n2005) );
  AOI22X1 U4434 ( .A(\data_in<14> ), .B(n1092), .C(n3591), .D(n1200), .Y(n3592) );
  OAI21X1 U4435 ( .A(n1349), .B(n3593), .C(n3592), .Y(n2006) );
  AOI22X1 U4436 ( .A(\data_in<15> ), .B(n1092), .C(n3594), .D(n1200), .Y(n3595) );
  OAI21X1 U4437 ( .A(n1349), .B(n3596), .C(n3595), .Y(n2007) );
  AOI22X1 U4438 ( .A(\data_in<8> ), .B(n1093), .C(n3598), .D(n1202), .Y(n3599)
         );
  OAI21X1 U4439 ( .A(n1351), .B(n3600), .C(n3599), .Y(n2008) );
  AOI22X1 U4440 ( .A(\data_in<9> ), .B(n1093), .C(n3601), .D(n1202), .Y(n3602)
         );
  OAI21X1 U4441 ( .A(n1351), .B(n3603), .C(n3602), .Y(n2009) );
  AOI22X1 U4442 ( .A(\data_in<10> ), .B(n1093), .C(n3604), .D(n1202), .Y(n3605) );
  OAI21X1 U4443 ( .A(n1351), .B(n3606), .C(n3605), .Y(n2010) );
  AOI22X1 U4444 ( .A(\data_in<11> ), .B(n1093), .C(n3607), .D(n1202), .Y(n3608) );
  OAI21X1 U4445 ( .A(n1351), .B(n3609), .C(n3608), .Y(n2011) );
  AOI22X1 U4446 ( .A(\data_in<12> ), .B(n1093), .C(n3610), .D(n1202), .Y(n3611) );
  OAI21X1 U4447 ( .A(n1351), .B(n3612), .C(n3611), .Y(n2012) );
  AOI22X1 U4448 ( .A(\data_in<13> ), .B(n1093), .C(n3613), .D(n1202), .Y(n3614) );
  OAI21X1 U4449 ( .A(n1351), .B(n3615), .C(n3614), .Y(n2013) );
  AOI22X1 U4450 ( .A(\data_in<14> ), .B(n1093), .C(n3616), .D(n1202), .Y(n3617) );
  OAI21X1 U4451 ( .A(n1351), .B(n3618), .C(n3617), .Y(n2014) );
  AOI22X1 U4452 ( .A(\data_in<15> ), .B(n1093), .C(n3619), .D(n1202), .Y(n3620) );
  OAI21X1 U4453 ( .A(n1351), .B(n3621), .C(n3620), .Y(n2015) );
  AOI22X1 U4454 ( .A(\data_in<8> ), .B(n1094), .C(n3622), .D(n1204), .Y(n3623)
         );
  OAI21X1 U4455 ( .A(n1353), .B(n3624), .C(n3623), .Y(n2016) );
  AOI22X1 U4456 ( .A(\data_in<9> ), .B(n1094), .C(n3625), .D(n1204), .Y(n3626)
         );
  OAI21X1 U4457 ( .A(n1353), .B(n3627), .C(n3626), .Y(n2017) );
  AOI22X1 U4458 ( .A(\data_in<10> ), .B(n1094), .C(n3628), .D(n1204), .Y(n3629) );
  OAI21X1 U4459 ( .A(n1353), .B(n3630), .C(n3629), .Y(n2018) );
  AOI22X1 U4460 ( .A(\data_in<11> ), .B(n1094), .C(n3631), .D(n1204), .Y(n3632) );
  OAI21X1 U4461 ( .A(n1353), .B(n3633), .C(n3632), .Y(n2019) );
  AOI22X1 U4462 ( .A(\data_in<12> ), .B(n1094), .C(n3634), .D(n1204), .Y(n3635) );
  OAI21X1 U4463 ( .A(n1353), .B(n3636), .C(n3635), .Y(n2020) );
  AOI22X1 U4464 ( .A(\data_in<13> ), .B(n1094), .C(n3637), .D(n1204), .Y(n3638) );
  OAI21X1 U4465 ( .A(n1353), .B(n3639), .C(n3638), .Y(n2021) );
  AOI22X1 U4466 ( .A(\data_in<14> ), .B(n1094), .C(n3640), .D(n1204), .Y(n3641) );
  OAI21X1 U4467 ( .A(n1353), .B(n3642), .C(n3641), .Y(n2022) );
  AOI22X1 U4468 ( .A(\data_in<15> ), .B(n1094), .C(n3643), .D(n1204), .Y(n3644) );
  OAI21X1 U4469 ( .A(n1353), .B(n3645), .C(n3644), .Y(n2023) );
  AOI22X1 U4470 ( .A(\data_in<8> ), .B(n1095), .C(n3647), .D(n1206), .Y(n3648)
         );
  OAI21X1 U4471 ( .A(n1355), .B(n3649), .C(n3648), .Y(n2024) );
  AOI22X1 U4472 ( .A(\data_in<9> ), .B(n1095), .C(n3650), .D(n1206), .Y(n3651)
         );
  OAI21X1 U4473 ( .A(n1355), .B(n3652), .C(n3651), .Y(n2025) );
  AOI22X1 U4474 ( .A(\data_in<10> ), .B(n1095), .C(n3653), .D(n1206), .Y(n3654) );
  OAI21X1 U4475 ( .A(n1355), .B(n3655), .C(n3654), .Y(n2026) );
  AOI22X1 U4476 ( .A(\data_in<11> ), .B(n1095), .C(n3656), .D(n1206), .Y(n3657) );
  OAI21X1 U4477 ( .A(n1355), .B(n3658), .C(n3657), .Y(n2027) );
  AOI22X1 U4478 ( .A(\data_in<12> ), .B(n1095), .C(n3659), .D(n1206), .Y(n3660) );
  OAI21X1 U4479 ( .A(n1355), .B(n3661), .C(n3660), .Y(n2028) );
  AOI22X1 U4480 ( .A(\data_in<13> ), .B(n1095), .C(n3662), .D(n1206), .Y(n3663) );
  OAI21X1 U4481 ( .A(n1355), .B(n3664), .C(n3663), .Y(n2029) );
  AOI22X1 U4482 ( .A(\data_in<14> ), .B(n1095), .C(n3665), .D(n1206), .Y(n3666) );
  OAI21X1 U4483 ( .A(n1355), .B(n3667), .C(n3666), .Y(n2030) );
  AOI22X1 U4484 ( .A(\data_in<15> ), .B(n1095), .C(n3668), .D(n1206), .Y(n3669) );
  OAI21X1 U4485 ( .A(n1355), .B(n3670), .C(n3669), .Y(n2031) );
  AOI22X1 U4486 ( .A(\data_in<8> ), .B(n1096), .C(n3672), .D(n1208), .Y(n3673)
         );
  OAI21X1 U4487 ( .A(n1357), .B(n3674), .C(n3673), .Y(n2032) );
  AOI22X1 U4488 ( .A(\data_in<9> ), .B(n1096), .C(n3675), .D(n1208), .Y(n3676)
         );
  OAI21X1 U4489 ( .A(n1357), .B(n3677), .C(n3676), .Y(n2033) );
  AOI22X1 U4490 ( .A(\data_in<10> ), .B(n1096), .C(n3678), .D(n1208), .Y(n3679) );
  OAI21X1 U4491 ( .A(n1357), .B(n3680), .C(n3679), .Y(n2034) );
  AOI22X1 U4492 ( .A(\data_in<11> ), .B(n1096), .C(n3681), .D(n1208), .Y(n3682) );
  OAI21X1 U4493 ( .A(n1357), .B(n3683), .C(n3682), .Y(n2035) );
  AOI22X1 U4494 ( .A(\data_in<12> ), .B(n1096), .C(n3684), .D(n1208), .Y(n3685) );
  OAI21X1 U4495 ( .A(n1357), .B(n3686), .C(n3685), .Y(n2036) );
  AOI22X1 U4496 ( .A(\data_in<13> ), .B(n1096), .C(n3687), .D(n1208), .Y(n3688) );
  OAI21X1 U4497 ( .A(n1357), .B(n3689), .C(n3688), .Y(n2037) );
  AOI22X1 U4498 ( .A(\data_in<14> ), .B(n1096), .C(n3690), .D(n1208), .Y(n3691) );
  OAI21X1 U4499 ( .A(n1357), .B(n3692), .C(n3691), .Y(n2038) );
  AOI22X1 U4500 ( .A(\data_in<15> ), .B(n1096), .C(n3693), .D(n1208), .Y(n3694) );
  OAI21X1 U4501 ( .A(n1357), .B(n3695), .C(n3694), .Y(n2039) );
  AOI22X1 U4502 ( .A(\data_in<8> ), .B(n1097), .C(n3697), .D(n1210), .Y(n3698)
         );
  OAI21X1 U4503 ( .A(n1359), .B(n3699), .C(n3698), .Y(n2040) );
  AOI22X1 U4504 ( .A(\data_in<9> ), .B(n1097), .C(n3700), .D(n1210), .Y(n3701)
         );
  OAI21X1 U4505 ( .A(n1359), .B(n3702), .C(n3701), .Y(n2041) );
  AOI22X1 U4506 ( .A(\data_in<10> ), .B(n1097), .C(n3703), .D(n1210), .Y(n3704) );
  OAI21X1 U4507 ( .A(n1359), .B(n3705), .C(n3704), .Y(n2042) );
  AOI22X1 U4508 ( .A(\data_in<11> ), .B(n1097), .C(n3706), .D(n1210), .Y(n3707) );
  OAI21X1 U4509 ( .A(n1359), .B(n3708), .C(n3707), .Y(n2043) );
  AOI22X1 U4510 ( .A(\data_in<12> ), .B(n1097), .C(n3709), .D(n1210), .Y(n3710) );
  OAI21X1 U4511 ( .A(n1359), .B(n3711), .C(n3710), .Y(n2044) );
  AOI22X1 U4512 ( .A(\data_in<13> ), .B(n1097), .C(n3712), .D(n1210), .Y(n3713) );
  OAI21X1 U4513 ( .A(n1359), .B(n3714), .C(n3713), .Y(n2045) );
  AOI22X1 U4514 ( .A(\data_in<14> ), .B(n1097), .C(n3715), .D(n1210), .Y(n3716) );
  OAI21X1 U4515 ( .A(n1359), .B(n3717), .C(n3716), .Y(n2046) );
  AOI22X1 U4516 ( .A(\data_in<15> ), .B(n1097), .C(n3718), .D(n1210), .Y(n3719) );
  OAI21X1 U4517 ( .A(n1359), .B(n3720), .C(n3719), .Y(n2047) );
  AOI22X1 U4518 ( .A(\data_in<8> ), .B(n1098), .C(n3722), .D(n1212), .Y(n3723)
         );
  OAI21X1 U4519 ( .A(n1361), .B(n3724), .C(n3723), .Y(n2048) );
  AOI22X1 U4520 ( .A(\data_in<9> ), .B(n1098), .C(n3725), .D(n1212), .Y(n3726)
         );
  OAI21X1 U4521 ( .A(n1361), .B(n3727), .C(n3726), .Y(n2049) );
  AOI22X1 U4522 ( .A(\data_in<10> ), .B(n1098), .C(n3728), .D(n1212), .Y(n3729) );
  OAI21X1 U4523 ( .A(n1361), .B(n3730), .C(n3729), .Y(n2050) );
  AOI22X1 U4524 ( .A(\data_in<11> ), .B(n1098), .C(n3731), .D(n1212), .Y(n3732) );
  OAI21X1 U4525 ( .A(n1361), .B(n3733), .C(n3732), .Y(n2051) );
  AOI22X1 U4526 ( .A(\data_in<12> ), .B(n1098), .C(n3734), .D(n1212), .Y(n3735) );
  OAI21X1 U4527 ( .A(n1361), .B(n3736), .C(n3735), .Y(n2052) );
  AOI22X1 U4528 ( .A(\data_in<13> ), .B(n1098), .C(n3737), .D(n1212), .Y(n3738) );
  OAI21X1 U4529 ( .A(n1361), .B(n3739), .C(n3738), .Y(n2053) );
  AOI22X1 U4530 ( .A(\data_in<14> ), .B(n1098), .C(n3740), .D(n1212), .Y(n3741) );
  OAI21X1 U4531 ( .A(n1361), .B(n3742), .C(n3741), .Y(n2054) );
  AOI22X1 U4532 ( .A(\data_in<15> ), .B(n1098), .C(n3743), .D(n1212), .Y(n3744) );
  OAI21X1 U4533 ( .A(n1361), .B(n3745), .C(n3744), .Y(n2055) );
  AOI22X1 U4534 ( .A(\data_in<8> ), .B(n1099), .C(n3748), .D(n1214), .Y(n3749)
         );
  OAI21X1 U4535 ( .A(n1363), .B(n3750), .C(n3749), .Y(n2056) );
  AOI22X1 U4536 ( .A(\data_in<9> ), .B(n1099), .C(n3751), .D(n1214), .Y(n3752)
         );
  OAI21X1 U4537 ( .A(n1363), .B(n3753), .C(n3752), .Y(n2057) );
  AOI22X1 U4538 ( .A(\data_in<10> ), .B(n1099), .C(n3754), .D(n1214), .Y(n3755) );
  OAI21X1 U4539 ( .A(n1363), .B(n3756), .C(n3755), .Y(n2058) );
  AOI22X1 U4540 ( .A(\data_in<11> ), .B(n1099), .C(n3757), .D(n1214), .Y(n3758) );
  OAI21X1 U4541 ( .A(n1363), .B(n3759), .C(n3758), .Y(n2059) );
  AOI22X1 U4542 ( .A(\data_in<12> ), .B(n1099), .C(n3760), .D(n1214), .Y(n3761) );
  OAI21X1 U4543 ( .A(n1363), .B(n3762), .C(n3761), .Y(n2060) );
  AOI22X1 U4544 ( .A(\data_in<13> ), .B(n1099), .C(n3763), .D(n1214), .Y(n3764) );
  OAI21X1 U4545 ( .A(n1363), .B(n3765), .C(n3764), .Y(n2061) );
  AOI22X1 U4546 ( .A(\data_in<14> ), .B(n1099), .C(n3766), .D(n1214), .Y(n3767) );
  OAI21X1 U4547 ( .A(n1363), .B(n3768), .C(n3767), .Y(n2062) );
  AOI22X1 U4548 ( .A(\data_in<15> ), .B(n1099), .C(n3769), .D(n1214), .Y(n3770) );
  OAI21X1 U4549 ( .A(n1363), .B(n3771), .C(n3770), .Y(n2063) );
  AOI22X1 U4550 ( .A(\data_in<8> ), .B(n1100), .C(n3773), .D(n1216), .Y(n3774)
         );
  OAI21X1 U4551 ( .A(n1365), .B(n3775), .C(n3774), .Y(n2064) );
  AOI22X1 U4552 ( .A(\data_in<9> ), .B(n1100), .C(n3776), .D(n1216), .Y(n3777)
         );
  OAI21X1 U4553 ( .A(n1365), .B(n3778), .C(n3777), .Y(n2065) );
  AOI22X1 U4554 ( .A(\data_in<10> ), .B(n1100), .C(n3779), .D(n1216), .Y(n3780) );
  OAI21X1 U4555 ( .A(n1365), .B(n3781), .C(n3780), .Y(n2066) );
  AOI22X1 U4556 ( .A(\data_in<11> ), .B(n1100), .C(n3782), .D(n1216), .Y(n3783) );
  OAI21X1 U4557 ( .A(n1365), .B(n3784), .C(n3783), .Y(n2067) );
  AOI22X1 U4558 ( .A(\data_in<12> ), .B(n1100), .C(n3785), .D(n1216), .Y(n3786) );
  OAI21X1 U4559 ( .A(n1365), .B(n3787), .C(n3786), .Y(n2068) );
  AOI22X1 U4560 ( .A(\data_in<13> ), .B(n1100), .C(n3788), .D(n1216), .Y(n3789) );
  OAI21X1 U4561 ( .A(n1365), .B(n3790), .C(n3789), .Y(n2069) );
  AOI22X1 U4562 ( .A(\data_in<14> ), .B(n1100), .C(n3791), .D(n1216), .Y(n3792) );
  OAI21X1 U4563 ( .A(n1365), .B(n3793), .C(n3792), .Y(n2070) );
  AOI22X1 U4564 ( .A(\data_in<15> ), .B(n1100), .C(n3794), .D(n1216), .Y(n3795) );
  OAI21X1 U4565 ( .A(n1365), .B(n3796), .C(n3795), .Y(n2071) );
  AOI22X1 U4566 ( .A(\data_in<8> ), .B(n1101), .C(n3799), .D(n1218), .Y(n3800)
         );
  OAI21X1 U4567 ( .A(n1367), .B(n3801), .C(n3800), .Y(n2072) );
  AOI22X1 U4568 ( .A(\data_in<9> ), .B(n1101), .C(n3802), .D(n1218), .Y(n3803)
         );
  OAI21X1 U4569 ( .A(n1367), .B(n3804), .C(n3803), .Y(n2073) );
  AOI22X1 U4570 ( .A(\data_in<10> ), .B(n1101), .C(n3805), .D(n1218), .Y(n3806) );
  OAI21X1 U4571 ( .A(n1367), .B(n3807), .C(n3806), .Y(n2074) );
  AOI22X1 U4572 ( .A(\data_in<11> ), .B(n1101), .C(n3808), .D(n1218), .Y(n3809) );
  OAI21X1 U4573 ( .A(n1367), .B(n3810), .C(n3809), .Y(n2075) );
  AOI22X1 U4574 ( .A(\data_in<12> ), .B(n1101), .C(n3811), .D(n1218), .Y(n3812) );
  OAI21X1 U4575 ( .A(n1367), .B(n3813), .C(n3812), .Y(n2076) );
  AOI22X1 U4576 ( .A(\data_in<13> ), .B(n1101), .C(n3814), .D(n1218), .Y(n3815) );
  OAI21X1 U4577 ( .A(n1367), .B(n3816), .C(n3815), .Y(n2077) );
  AOI22X1 U4578 ( .A(\data_in<14> ), .B(n1101), .C(n3817), .D(n1218), .Y(n3818) );
  OAI21X1 U4579 ( .A(n1367), .B(n3819), .C(n3818), .Y(n2078) );
  AOI22X1 U4580 ( .A(\data_in<15> ), .B(n1101), .C(n3820), .D(n1218), .Y(n3821) );
  OAI21X1 U4581 ( .A(n1367), .B(n3822), .C(n3821), .Y(n2079) );
  AOI22X1 U4582 ( .A(\data_in<8> ), .B(n1102), .C(n3824), .D(n1220), .Y(n3825)
         );
  OAI21X1 U4583 ( .A(n1369), .B(n3826), .C(n3825), .Y(n2080) );
  AOI22X1 U4584 ( .A(\data_in<9> ), .B(n1102), .C(n3827), .D(n1220), .Y(n3828)
         );
  OAI21X1 U4585 ( .A(n1369), .B(n3829), .C(n3828), .Y(n2081) );
  AOI22X1 U4586 ( .A(\data_in<10> ), .B(n1102), .C(n3830), .D(n1220), .Y(n3831) );
  OAI21X1 U4587 ( .A(n1369), .B(n3832), .C(n3831), .Y(n2082) );
  AOI22X1 U4588 ( .A(\data_in<11> ), .B(n1102), .C(n3833), .D(n1220), .Y(n3834) );
  OAI21X1 U4589 ( .A(n1369), .B(n3835), .C(n3834), .Y(n2083) );
  AOI22X1 U4590 ( .A(\data_in<12> ), .B(n1102), .C(n3836), .D(n1220), .Y(n3837) );
  OAI21X1 U4591 ( .A(n1369), .B(n3838), .C(n3837), .Y(n2084) );
  AOI22X1 U4592 ( .A(\data_in<13> ), .B(n1102), .C(n3839), .D(n1220), .Y(n3840) );
  OAI21X1 U4593 ( .A(n1369), .B(n3841), .C(n3840), .Y(n2085) );
  AOI22X1 U4594 ( .A(\data_in<14> ), .B(n1102), .C(n3842), .D(n1220), .Y(n3843) );
  OAI21X1 U4595 ( .A(n1369), .B(n3844), .C(n3843), .Y(n2086) );
  AOI22X1 U4596 ( .A(\data_in<15> ), .B(n1102), .C(n3845), .D(n1220), .Y(n3846) );
  OAI21X1 U4597 ( .A(n1369), .B(n3847), .C(n3846), .Y(n2087) );
  AOI22X1 U4598 ( .A(\data_in<8> ), .B(n1103), .C(n3850), .D(n1222), .Y(n3851)
         );
  OAI21X1 U4599 ( .A(n1371), .B(n3852), .C(n3851), .Y(n2088) );
  AOI22X1 U4600 ( .A(\data_in<9> ), .B(n1103), .C(n3853), .D(n1222), .Y(n3854)
         );
  OAI21X1 U4601 ( .A(n1371), .B(n3855), .C(n3854), .Y(n2089) );
  AOI22X1 U4602 ( .A(\data_in<10> ), .B(n1103), .C(n3856), .D(n1222), .Y(n3857) );
  OAI21X1 U4603 ( .A(n1371), .B(n3858), .C(n3857), .Y(n2090) );
  AOI22X1 U4604 ( .A(\data_in<11> ), .B(n1103), .C(n3859), .D(n1222), .Y(n3860) );
  OAI21X1 U4605 ( .A(n1371), .B(n3861), .C(n3860), .Y(n2091) );
  AOI22X1 U4606 ( .A(\data_in<12> ), .B(n1103), .C(n3862), .D(n1222), .Y(n3863) );
  OAI21X1 U4607 ( .A(n1371), .B(n3864), .C(n3863), .Y(n2092) );
  AOI22X1 U4608 ( .A(\data_in<13> ), .B(n1103), .C(n3865), .D(n1222), .Y(n3866) );
  OAI21X1 U4609 ( .A(n1371), .B(n3867), .C(n3866), .Y(n2093) );
  AOI22X1 U4610 ( .A(\data_in<14> ), .B(n1103), .C(n3868), .D(n1222), .Y(n3869) );
  OAI21X1 U4611 ( .A(n1371), .B(n3870), .C(n3869), .Y(n2094) );
  AOI22X1 U4612 ( .A(\data_in<15> ), .B(n1103), .C(n3871), .D(n1222), .Y(n3872) );
  OAI21X1 U4613 ( .A(n1371), .B(n3873), .C(n3872), .Y(n2095) );
  AOI22X1 U4614 ( .A(\data_in<8> ), .B(n1104), .C(n3876), .D(n1224), .Y(n3877)
         );
  OAI21X1 U4615 ( .A(n1373), .B(n3878), .C(n3877), .Y(n2096) );
  AOI22X1 U4616 ( .A(\data_in<9> ), .B(n1104), .C(n3879), .D(n1224), .Y(n3880)
         );
  OAI21X1 U4617 ( .A(n1373), .B(n3881), .C(n3880), .Y(n2097) );
  AOI22X1 U4618 ( .A(\data_in<10> ), .B(n1104), .C(n3882), .D(n1224), .Y(n3883) );
  OAI21X1 U4619 ( .A(n1373), .B(n3884), .C(n3883), .Y(n2098) );
  AOI22X1 U4620 ( .A(\data_in<11> ), .B(n1104), .C(n3885), .D(n1224), .Y(n3886) );
  OAI21X1 U4621 ( .A(n1373), .B(n3887), .C(n3886), .Y(n2099) );
  AOI22X1 U4622 ( .A(\data_in<12> ), .B(n1104), .C(n3888), .D(n1224), .Y(n3889) );
  OAI21X1 U4623 ( .A(n1373), .B(n3890), .C(n3889), .Y(n2100) );
  AOI22X1 U4624 ( .A(\data_in<13> ), .B(n1104), .C(n3891), .D(n1224), .Y(n3892) );
  OAI21X1 U4625 ( .A(n1373), .B(n3893), .C(n3892), .Y(n2101) );
  AOI22X1 U4626 ( .A(\data_in<14> ), .B(n1104), .C(n3894), .D(n1224), .Y(n3895) );
  OAI21X1 U4627 ( .A(n1373), .B(n3896), .C(n3895), .Y(n2102) );
  AOI22X1 U4628 ( .A(\data_in<15> ), .B(n1104), .C(n3897), .D(n1224), .Y(n3898) );
  OAI21X1 U4629 ( .A(n1373), .B(n3899), .C(n3898), .Y(n2103) );
  AOI22X1 U4630 ( .A(\data_in<8> ), .B(n1105), .C(n3902), .D(n1226), .Y(n3903)
         );
  OAI21X1 U4631 ( .A(n1375), .B(n3904), .C(n3903), .Y(n2104) );
  AOI22X1 U4632 ( .A(\data_in<9> ), .B(n1105), .C(n3905), .D(n1226), .Y(n3906)
         );
  OAI21X1 U4633 ( .A(n1375), .B(n3907), .C(n3906), .Y(n2105) );
  AOI22X1 U4634 ( .A(\data_in<10> ), .B(n1105), .C(n3908), .D(n1226), .Y(n3909) );
  OAI21X1 U4635 ( .A(n1375), .B(n3910), .C(n3909), .Y(n2106) );
  AOI22X1 U4636 ( .A(\data_in<11> ), .B(n1105), .C(n3911), .D(n1226), .Y(n3912) );
  OAI21X1 U4637 ( .A(n1375), .B(n3913), .C(n3912), .Y(n2107) );
  AOI22X1 U4638 ( .A(\data_in<12> ), .B(n1105), .C(n3914), .D(n1226), .Y(n3915) );
  OAI21X1 U4639 ( .A(n1375), .B(n3916), .C(n3915), .Y(n2108) );
  AOI22X1 U4640 ( .A(\data_in<13> ), .B(n1105), .C(n3917), .D(n1226), .Y(n3918) );
  OAI21X1 U4641 ( .A(n1375), .B(n3919), .C(n3918), .Y(n2109) );
  AOI22X1 U4642 ( .A(\data_in<14> ), .B(n1105), .C(n3920), .D(n1226), .Y(n3921) );
  OAI21X1 U4643 ( .A(n1375), .B(n3922), .C(n3921), .Y(n2110) );
  AOI22X1 U4644 ( .A(\data_in<15> ), .B(n1105), .C(n3923), .D(n1226), .Y(n3924) );
  OAI21X1 U4645 ( .A(n1375), .B(n3925), .C(n3924), .Y(n2111) );
  AOI22X1 U4646 ( .A(\data_in<8> ), .B(n1106), .C(n3928), .D(n1228), .Y(n3929)
         );
  OAI21X1 U4647 ( .A(n1377), .B(n3930), .C(n3929), .Y(n2112) );
  AOI22X1 U4648 ( .A(\data_in<9> ), .B(n1106), .C(n3931), .D(n1228), .Y(n3932)
         );
  OAI21X1 U4649 ( .A(n1377), .B(n3933), .C(n3932), .Y(n2113) );
  AOI22X1 U4650 ( .A(\data_in<10> ), .B(n1106), .C(n3934), .D(n1228), .Y(n3935) );
  OAI21X1 U4651 ( .A(n1377), .B(n3936), .C(n3935), .Y(n2114) );
  AOI22X1 U4652 ( .A(\data_in<11> ), .B(n1106), .C(n3937), .D(n1228), .Y(n3938) );
  OAI21X1 U4653 ( .A(n1377), .B(n3939), .C(n3938), .Y(n2115) );
  AOI22X1 U4654 ( .A(\data_in<12> ), .B(n1106), .C(n3940), .D(n1228), .Y(n3941) );
  OAI21X1 U4655 ( .A(n1377), .B(n3942), .C(n3941), .Y(n2116) );
  AOI22X1 U4656 ( .A(\data_in<13> ), .B(n1106), .C(n3943), .D(n1228), .Y(n3944) );
  OAI21X1 U4657 ( .A(n1377), .B(n3945), .C(n3944), .Y(n2117) );
  AOI22X1 U4658 ( .A(\data_in<14> ), .B(n1106), .C(n3946), .D(n1228), .Y(n3947) );
  OAI21X1 U4659 ( .A(n1377), .B(n3948), .C(n3947), .Y(n2118) );
  AOI22X1 U4660 ( .A(\data_in<15> ), .B(n1106), .C(n3949), .D(n1228), .Y(n3950) );
  OAI21X1 U4661 ( .A(n1377), .B(n3951), .C(n3950), .Y(n2119) );
  AOI22X1 U4662 ( .A(\data_in<8> ), .B(n1107), .C(n3954), .D(n1230), .Y(n3955)
         );
  OAI21X1 U4663 ( .A(n1379), .B(n3956), .C(n3955), .Y(n2120) );
  AOI22X1 U4664 ( .A(\data_in<9> ), .B(n1107), .C(n3957), .D(n1230), .Y(n3958)
         );
  OAI21X1 U4665 ( .A(n1379), .B(n3959), .C(n3958), .Y(n2121) );
  AOI22X1 U4666 ( .A(\data_in<10> ), .B(n1107), .C(n3960), .D(n1230), .Y(n3961) );
  OAI21X1 U4667 ( .A(n1379), .B(n3962), .C(n3961), .Y(n2122) );
  AOI22X1 U4668 ( .A(\data_in<11> ), .B(n1107), .C(n3963), .D(n1230), .Y(n3964) );
  OAI21X1 U4669 ( .A(n1379), .B(n3965), .C(n3964), .Y(n2123) );
  AOI22X1 U4670 ( .A(\data_in<12> ), .B(n1107), .C(n3966), .D(n1230), .Y(n3967) );
  OAI21X1 U4671 ( .A(n1379), .B(n3968), .C(n3967), .Y(n2124) );
  AOI22X1 U4672 ( .A(\data_in<13> ), .B(n1107), .C(n3969), .D(n1230), .Y(n3970) );
  OAI21X1 U4673 ( .A(n1379), .B(n3971), .C(n3970), .Y(n2125) );
  AOI22X1 U4674 ( .A(\data_in<14> ), .B(n1107), .C(n3972), .D(n1230), .Y(n3973) );
  OAI21X1 U4675 ( .A(n1379), .B(n3974), .C(n3973), .Y(n2126) );
  AOI22X1 U4676 ( .A(\data_in<15> ), .B(n1107), .C(n3975), .D(n1230), .Y(n3976) );
  OAI21X1 U4677 ( .A(n1379), .B(n3977), .C(n3976), .Y(n2127) );
  AOI22X1 U4678 ( .A(\data_in<8> ), .B(n1108), .C(n3979), .D(n1232), .Y(n3980)
         );
  OAI21X1 U4679 ( .A(n1381), .B(n3981), .C(n3980), .Y(n2128) );
  AOI22X1 U4680 ( .A(\data_in<9> ), .B(n1108), .C(n3982), .D(n1232), .Y(n3983)
         );
  OAI21X1 U4681 ( .A(n1381), .B(n3984), .C(n3983), .Y(n2129) );
  AOI22X1 U4682 ( .A(\data_in<10> ), .B(n1108), .C(n3985), .D(n1232), .Y(n3986) );
  OAI21X1 U4683 ( .A(n1381), .B(n3987), .C(n3986), .Y(n2130) );
  AOI22X1 U4684 ( .A(\data_in<11> ), .B(n1108), .C(n3988), .D(n1232), .Y(n3989) );
  OAI21X1 U4685 ( .A(n1381), .B(n3990), .C(n3989), .Y(n2131) );
  AOI22X1 U4686 ( .A(\data_in<12> ), .B(n1108), .C(n3991), .D(n1232), .Y(n3992) );
  OAI21X1 U4687 ( .A(n1381), .B(n3993), .C(n3992), .Y(n2132) );
  AOI22X1 U4688 ( .A(\data_in<13> ), .B(n1108), .C(n3994), .D(n1232), .Y(n3995) );
  OAI21X1 U4689 ( .A(n1381), .B(n3996), .C(n3995), .Y(n2133) );
  AOI22X1 U4690 ( .A(\data_in<14> ), .B(n1108), .C(n3997), .D(n1232), .Y(n3998) );
  OAI21X1 U4691 ( .A(n1381), .B(n3999), .C(n3998), .Y(n2134) );
  AOI22X1 U4692 ( .A(\data_in<15> ), .B(n1108), .C(n4000), .D(n1232), .Y(n4001) );
  OAI21X1 U4693 ( .A(n1381), .B(n4002), .C(n4001), .Y(n2135) );
  AOI22X1 U4694 ( .A(\data_in<8> ), .B(n1109), .C(n4004), .D(n1234), .Y(n4005)
         );
  OAI21X1 U4695 ( .A(n1383), .B(n4006), .C(n4005), .Y(n2136) );
  AOI22X1 U4696 ( .A(\data_in<9> ), .B(n1109), .C(n4007), .D(n1234), .Y(n4008)
         );
  OAI21X1 U4697 ( .A(n1383), .B(n4009), .C(n4008), .Y(n2137) );
  AOI22X1 U4698 ( .A(\data_in<10> ), .B(n1109), .C(n4010), .D(n1234), .Y(n4011) );
  OAI21X1 U4699 ( .A(n1383), .B(n4012), .C(n4011), .Y(n2138) );
  AOI22X1 U4700 ( .A(\data_in<11> ), .B(n1109), .C(n4013), .D(n1234), .Y(n4014) );
  OAI21X1 U4701 ( .A(n1383), .B(n4015), .C(n4014), .Y(n2139) );
  AOI22X1 U4702 ( .A(\data_in<12> ), .B(n1109), .C(n4016), .D(n1234), .Y(n4017) );
  OAI21X1 U4703 ( .A(n1383), .B(n4018), .C(n4017), .Y(n2140) );
  AOI22X1 U4704 ( .A(\data_in<13> ), .B(n1109), .C(n4019), .D(n1234), .Y(n4020) );
  OAI21X1 U4705 ( .A(n1383), .B(n4021), .C(n4020), .Y(n2141) );
  AOI22X1 U4706 ( .A(\data_in<14> ), .B(n1109), .C(n4022), .D(n1234), .Y(n4023) );
  OAI21X1 U4707 ( .A(n1383), .B(n4024), .C(n4023), .Y(n2142) );
  AOI22X1 U4708 ( .A(\data_in<15> ), .B(n1109), .C(n4025), .D(n1234), .Y(n4026) );
  OAI21X1 U4709 ( .A(n1383), .B(n4027), .C(n4026), .Y(n2143) );
  AOI22X1 U4710 ( .A(\data_in<8> ), .B(n1110), .C(n4029), .D(n1236), .Y(n4030)
         );
  OAI21X1 U4711 ( .A(n1385), .B(n4031), .C(n4030), .Y(n2144) );
  AOI22X1 U4712 ( .A(\data_in<9> ), .B(n1110), .C(n4032), .D(n1236), .Y(n4033)
         );
  OAI21X1 U4713 ( .A(n1385), .B(n4034), .C(n4033), .Y(n2145) );
  AOI22X1 U4714 ( .A(\data_in<10> ), .B(n1110), .C(n4035), .D(n1236), .Y(n4036) );
  OAI21X1 U4715 ( .A(n1385), .B(n4037), .C(n4036), .Y(n2146) );
  AOI22X1 U4716 ( .A(\data_in<11> ), .B(n1110), .C(n4038), .D(n1236), .Y(n4039) );
  OAI21X1 U4717 ( .A(n1385), .B(n4040), .C(n4039), .Y(n2147) );
  AOI22X1 U4718 ( .A(\data_in<12> ), .B(n1110), .C(n4041), .D(n1236), .Y(n4042) );
  OAI21X1 U4719 ( .A(n1385), .B(n4043), .C(n4042), .Y(n2148) );
  AOI22X1 U4720 ( .A(\data_in<13> ), .B(n1110), .C(n4044), .D(n1236), .Y(n4045) );
  OAI21X1 U4721 ( .A(n1385), .B(n4046), .C(n4045), .Y(n2149) );
  AOI22X1 U4722 ( .A(\data_in<14> ), .B(n1110), .C(n4047), .D(n1236), .Y(n4048) );
  OAI21X1 U4723 ( .A(n1385), .B(n4049), .C(n4048), .Y(n2150) );
  AOI22X1 U4724 ( .A(\data_in<15> ), .B(n1110), .C(n4050), .D(n1236), .Y(n4051) );
  OAI21X1 U4725 ( .A(n1385), .B(n4052), .C(n4051), .Y(n2151) );
  AOI22X1 U4726 ( .A(\data_in<8> ), .B(n1111), .C(n4054), .D(n1238), .Y(n4055)
         );
  OAI21X1 U4727 ( .A(n1387), .B(n4056), .C(n4055), .Y(n2152) );
  AOI22X1 U4728 ( .A(\data_in<9> ), .B(n1111), .C(n4057), .D(n1238), .Y(n4058)
         );
  OAI21X1 U4729 ( .A(n1387), .B(n4059), .C(n4058), .Y(n2153) );
  AOI22X1 U4730 ( .A(\data_in<10> ), .B(n1111), .C(n4060), .D(n1238), .Y(n4061) );
  OAI21X1 U4731 ( .A(n1387), .B(n4062), .C(n4061), .Y(n2154) );
  AOI22X1 U4732 ( .A(\data_in<11> ), .B(n1111), .C(n4063), .D(n1238), .Y(n4064) );
  OAI21X1 U4733 ( .A(n1387), .B(n4065), .C(n4064), .Y(n2155) );
  AOI22X1 U4734 ( .A(\data_in<12> ), .B(n1111), .C(n4066), .D(n1238), .Y(n4067) );
  OAI21X1 U4735 ( .A(n1387), .B(n4068), .C(n4067), .Y(n2156) );
  AOI22X1 U4736 ( .A(\data_in<13> ), .B(n1111), .C(n4069), .D(n1238), .Y(n4070) );
  OAI21X1 U4737 ( .A(n1387), .B(n4071), .C(n4070), .Y(n2157) );
  AOI22X1 U4738 ( .A(\data_in<14> ), .B(n1111), .C(n4072), .D(n1238), .Y(n4073) );
  OAI21X1 U4739 ( .A(n1387), .B(n4074), .C(n4073), .Y(n2158) );
  AOI22X1 U4740 ( .A(\data_in<15> ), .B(n1111), .C(n4075), .D(n1238), .Y(n4076) );
  OAI21X1 U4741 ( .A(n1387), .B(n4077), .C(n4076), .Y(n2159) );
  AOI22X1 U4742 ( .A(\data_in<8> ), .B(n1112), .C(n4079), .D(n1240), .Y(n4080)
         );
  OAI21X1 U4743 ( .A(n1389), .B(n4081), .C(n4080), .Y(n2160) );
  AOI22X1 U4744 ( .A(\data_in<9> ), .B(n1112), .C(n4082), .D(n1240), .Y(n4083)
         );
  OAI21X1 U4745 ( .A(n1389), .B(n4084), .C(n4083), .Y(n2161) );
  AOI22X1 U4746 ( .A(\data_in<10> ), .B(n1112), .C(n4085), .D(n1240), .Y(n4086) );
  OAI21X1 U4747 ( .A(n1389), .B(n4087), .C(n4086), .Y(n2162) );
  AOI22X1 U4748 ( .A(\data_in<11> ), .B(n1112), .C(n4088), .D(n1240), .Y(n4089) );
  OAI21X1 U4749 ( .A(n1389), .B(n4090), .C(n4089), .Y(n2163) );
  AOI22X1 U4750 ( .A(\data_in<12> ), .B(n1112), .C(n4091), .D(n1240), .Y(n4092) );
  OAI21X1 U4751 ( .A(n1389), .B(n4093), .C(n4092), .Y(n2164) );
  AOI22X1 U4752 ( .A(\data_in<13> ), .B(n1112), .C(n4094), .D(n1240), .Y(n4095) );
  OAI21X1 U4753 ( .A(n1389), .B(n4096), .C(n4095), .Y(n2165) );
  AOI22X1 U4754 ( .A(\data_in<14> ), .B(n1112), .C(n4097), .D(n1240), .Y(n4098) );
  OAI21X1 U4755 ( .A(n1389), .B(n4099), .C(n4098), .Y(n2166) );
  AOI22X1 U4756 ( .A(\data_in<15> ), .B(n1112), .C(n4100), .D(n1240), .Y(n4101) );
  OAI21X1 U4757 ( .A(n1389), .B(n4102), .C(n4101), .Y(n2167) );
  AOI22X1 U4758 ( .A(\data_in<8> ), .B(n1113), .C(n4104), .D(n1242), .Y(n4105)
         );
  OAI21X1 U4759 ( .A(n1391), .B(n4106), .C(n4105), .Y(n2168) );
  AOI22X1 U4760 ( .A(\data_in<9> ), .B(n1113), .C(n4107), .D(n1242), .Y(n4108)
         );
  OAI21X1 U4761 ( .A(n1391), .B(n4109), .C(n4108), .Y(n2169) );
  AOI22X1 U4762 ( .A(\data_in<10> ), .B(n1113), .C(n4110), .D(n1242), .Y(n4111) );
  OAI21X1 U4763 ( .A(n1391), .B(n4112), .C(n4111), .Y(n2170) );
  AOI22X1 U4764 ( .A(\data_in<11> ), .B(n1113), .C(n4113), .D(n1242), .Y(n4114) );
  OAI21X1 U4765 ( .A(n1391), .B(n4115), .C(n4114), .Y(n2171) );
  AOI22X1 U4766 ( .A(\data_in<12> ), .B(n1113), .C(n4116), .D(n1242), .Y(n4117) );
  OAI21X1 U4767 ( .A(n1391), .B(n4118), .C(n4117), .Y(n2172) );
  AOI22X1 U4768 ( .A(\data_in<13> ), .B(n1113), .C(n4119), .D(n1242), .Y(n4120) );
  OAI21X1 U4769 ( .A(n1391), .B(n4121), .C(n4120), .Y(n2173) );
  AOI22X1 U4770 ( .A(\data_in<14> ), .B(n1113), .C(n4122), .D(n1242), .Y(n4123) );
  OAI21X1 U4771 ( .A(n1391), .B(n4124), .C(n4123), .Y(n2174) );
  AOI22X1 U4772 ( .A(\data_in<15> ), .B(n1113), .C(n4125), .D(n1242), .Y(n4126) );
  OAI21X1 U4773 ( .A(n1391), .B(n4127), .C(n4126), .Y(n2175) );
  AOI22X1 U4774 ( .A(\data_in<8> ), .B(n1114), .C(n4129), .D(n1244), .Y(n4130)
         );
  OAI21X1 U4775 ( .A(n1393), .B(n4131), .C(n4130), .Y(n2176) );
  AOI22X1 U4776 ( .A(\data_in<9> ), .B(n1114), .C(n4132), .D(n1244), .Y(n4133)
         );
  OAI21X1 U4777 ( .A(n1393), .B(n4134), .C(n4133), .Y(n2177) );
  AOI22X1 U4778 ( .A(\data_in<10> ), .B(n1114), .C(n4135), .D(n1244), .Y(n4136) );
  OAI21X1 U4779 ( .A(n1393), .B(n4137), .C(n4136), .Y(n2178) );
  AOI22X1 U4780 ( .A(\data_in<11> ), .B(n1114), .C(n4138), .D(n1244), .Y(n4139) );
  OAI21X1 U4781 ( .A(n1393), .B(n4140), .C(n4139), .Y(n2179) );
  AOI22X1 U4782 ( .A(\data_in<12> ), .B(n1114), .C(n4141), .D(n1244), .Y(n4142) );
  OAI21X1 U4783 ( .A(n1393), .B(n4143), .C(n4142), .Y(n2180) );
  AOI22X1 U4784 ( .A(\data_in<13> ), .B(n1114), .C(n4144), .D(n1244), .Y(n4145) );
  OAI21X1 U4785 ( .A(n1393), .B(n4146), .C(n4145), .Y(n2181) );
  AOI22X1 U4786 ( .A(\data_in<14> ), .B(n1114), .C(n4147), .D(n1244), .Y(n4148) );
  OAI21X1 U4787 ( .A(n1393), .B(n4149), .C(n4148), .Y(n2182) );
  AOI22X1 U4788 ( .A(\data_in<15> ), .B(n1114), .C(n4150), .D(n1244), .Y(n4151) );
  OAI21X1 U4789 ( .A(n1393), .B(n4152), .C(n4151), .Y(n2183) );
  AOI22X1 U4790 ( .A(\data_in<8> ), .B(n1115), .C(n4154), .D(n1246), .Y(n4155)
         );
  OAI21X1 U4791 ( .A(n1395), .B(n4156), .C(n4155), .Y(n2184) );
  AOI22X1 U4792 ( .A(\data_in<9> ), .B(n1115), .C(n4157), .D(n1246), .Y(n4158)
         );
  OAI21X1 U4793 ( .A(n1395), .B(n4159), .C(n4158), .Y(n2185) );
  AOI22X1 U4794 ( .A(\data_in<10> ), .B(n1115), .C(n4160), .D(n1246), .Y(n4161) );
  OAI21X1 U4795 ( .A(n1395), .B(n4162), .C(n4161), .Y(n2186) );
  AOI22X1 U4796 ( .A(\data_in<11> ), .B(n1115), .C(n4163), .D(n1246), .Y(n4164) );
  OAI21X1 U4797 ( .A(n1395), .B(n4165), .C(n4164), .Y(n2187) );
  AOI22X1 U4798 ( .A(\data_in<12> ), .B(n1115), .C(n4166), .D(n1246), .Y(n4167) );
  OAI21X1 U4799 ( .A(n1395), .B(n4168), .C(n4167), .Y(n2188) );
  AOI22X1 U4800 ( .A(\data_in<13> ), .B(n1115), .C(n4169), .D(n1246), .Y(n4170) );
  OAI21X1 U4801 ( .A(n1395), .B(n4171), .C(n4170), .Y(n2189) );
  AOI22X1 U4802 ( .A(\data_in<14> ), .B(n1115), .C(n4172), .D(n1246), .Y(n4173) );
  OAI21X1 U4803 ( .A(n1395), .B(n4174), .C(n4173), .Y(n2190) );
  AOI22X1 U4804 ( .A(\data_in<15> ), .B(n1115), .C(n4175), .D(n1246), .Y(n4176) );
  OAI21X1 U4805 ( .A(n1395), .B(n4177), .C(n4176), .Y(n2191) );
  AOI22X1 U4806 ( .A(\data_in<8> ), .B(n1116), .C(n4178), .D(n1248), .Y(n4179)
         );
  OAI21X1 U4807 ( .A(n1397), .B(n4180), .C(n4179), .Y(n2192) );
  AOI22X1 U4808 ( .A(\data_in<9> ), .B(n1116), .C(n4181), .D(n1248), .Y(n4182)
         );
  OAI21X1 U4809 ( .A(n1397), .B(n4183), .C(n4182), .Y(n2193) );
  AOI22X1 U4810 ( .A(\data_in<10> ), .B(n1116), .C(n4184), .D(n1248), .Y(n4185) );
  OAI21X1 U4811 ( .A(n1397), .B(n4186), .C(n4185), .Y(n2194) );
  AOI22X1 U4812 ( .A(\data_in<11> ), .B(n1116), .C(n4187), .D(n1248), .Y(n4188) );
  OAI21X1 U4813 ( .A(n1397), .B(n4189), .C(n4188), .Y(n2195) );
  AOI22X1 U4814 ( .A(\data_in<12> ), .B(n1116), .C(n4190), .D(n1248), .Y(n4191) );
  OAI21X1 U4815 ( .A(n1397), .B(n4192), .C(n4191), .Y(n2196) );
  AOI22X1 U4816 ( .A(\data_in<13> ), .B(n1116), .C(n4193), .D(n1248), .Y(n4194) );
  OAI21X1 U4817 ( .A(n1397), .B(n4195), .C(n4194), .Y(n2197) );
  AOI22X1 U4818 ( .A(\data_in<14> ), .B(n1116), .C(n4196), .D(n1248), .Y(n4197) );
  OAI21X1 U4819 ( .A(n1397), .B(n4198), .C(n4197), .Y(n2198) );
  AOI22X1 U4820 ( .A(\data_in<15> ), .B(n1116), .C(n4199), .D(n1248), .Y(n4200) );
  OAI21X1 U4821 ( .A(n1397), .B(n4201), .C(n4200), .Y(n2199) );
  AOI22X1 U4822 ( .A(\data_in<8> ), .B(n1117), .C(n4204), .D(n1250), .Y(n4205)
         );
  OAI21X1 U4823 ( .A(n1399), .B(n4206), .C(n4205), .Y(n2200) );
  AOI22X1 U4824 ( .A(\data_in<9> ), .B(n1117), .C(n4207), .D(n1250), .Y(n4208)
         );
  OAI21X1 U4825 ( .A(n1399), .B(n4209), .C(n4208), .Y(n2201) );
  AOI22X1 U4826 ( .A(\data_in<10> ), .B(n1117), .C(n4210), .D(n1250), .Y(n4211) );
  OAI21X1 U4827 ( .A(n1399), .B(n4212), .C(n4211), .Y(n2202) );
  AOI22X1 U4828 ( .A(\data_in<11> ), .B(n1117), .C(n4213), .D(n1250), .Y(n4214) );
  OAI21X1 U4829 ( .A(n1399), .B(n4215), .C(n4214), .Y(n2203) );
  AOI22X1 U4830 ( .A(\data_in<12> ), .B(n1117), .C(n4216), .D(n1250), .Y(n4217) );
  OAI21X1 U4831 ( .A(n1399), .B(n4218), .C(n4217), .Y(n2204) );
  AOI22X1 U4832 ( .A(\data_in<13> ), .B(n1117), .C(n4219), .D(n1250), .Y(n4220) );
  OAI21X1 U4833 ( .A(n1399), .B(n4221), .C(n4220), .Y(n2205) );
  AOI22X1 U4834 ( .A(\data_in<14> ), .B(n1117), .C(n4222), .D(n1250), .Y(n4223) );
  OAI21X1 U4835 ( .A(n1399), .B(n4224), .C(n4223), .Y(n2206) );
  AOI22X1 U4836 ( .A(\data_in<15> ), .B(n1117), .C(n4225), .D(n1250), .Y(n4226) );
  OAI21X1 U4837 ( .A(n1399), .B(n4227), .C(n4226), .Y(n2207) );
  AOI22X1 U4838 ( .A(\data_in<8> ), .B(n1118), .C(n4228), .D(n1252), .Y(n4229)
         );
  OAI21X1 U4839 ( .A(n1401), .B(n4230), .C(n4229), .Y(n2208) );
  AOI22X1 U4840 ( .A(\data_in<9> ), .B(n1118), .C(n4231), .D(n1252), .Y(n4232)
         );
  OAI21X1 U4841 ( .A(n1401), .B(n4233), .C(n4232), .Y(n2209) );
  AOI22X1 U4842 ( .A(\data_in<10> ), .B(n1118), .C(n4234), .D(n1252), .Y(n4235) );
  OAI21X1 U4843 ( .A(n1401), .B(n4236), .C(n4235), .Y(n2210) );
  AOI22X1 U4844 ( .A(\data_in<11> ), .B(n1118), .C(n4237), .D(n1252), .Y(n4238) );
  OAI21X1 U4845 ( .A(n1401), .B(n4239), .C(n4238), .Y(n2211) );
  AOI22X1 U4846 ( .A(\data_in<12> ), .B(n1118), .C(n4240), .D(n1252), .Y(n4241) );
  OAI21X1 U4847 ( .A(n1401), .B(n4242), .C(n4241), .Y(n2212) );
  AOI22X1 U4848 ( .A(\data_in<13> ), .B(n1118), .C(n4243), .D(n1252), .Y(n4244) );
  OAI21X1 U4849 ( .A(n1401), .B(n4245), .C(n4244), .Y(n2213) );
  AOI22X1 U4850 ( .A(\data_in<14> ), .B(n1118), .C(n4246), .D(n1252), .Y(n4247) );
  OAI21X1 U4851 ( .A(n1401), .B(n4248), .C(n4247), .Y(n2214) );
  AOI22X1 U4852 ( .A(\data_in<15> ), .B(n1118), .C(n4249), .D(n1252), .Y(n4250) );
  OAI21X1 U4853 ( .A(n1401), .B(n4251), .C(n4250), .Y(n2215) );
  AOI22X1 U4854 ( .A(\data_in<8> ), .B(n1119), .C(n4253), .D(n1254), .Y(n4254)
         );
  OAI21X1 U4855 ( .A(n1403), .B(n4255), .C(n4254), .Y(n2216) );
  AOI22X1 U4856 ( .A(\data_in<9> ), .B(n1119), .C(n4256), .D(n1254), .Y(n4257)
         );
  OAI21X1 U4857 ( .A(n1403), .B(n4258), .C(n4257), .Y(n2217) );
  AOI22X1 U4858 ( .A(\data_in<10> ), .B(n1119), .C(n4259), .D(n1254), .Y(n4260) );
  OAI21X1 U4859 ( .A(n1403), .B(n4261), .C(n4260), .Y(n2218) );
  AOI22X1 U4860 ( .A(\data_in<11> ), .B(n1119), .C(n4262), .D(n1254), .Y(n4263) );
  OAI21X1 U4861 ( .A(n1403), .B(n4264), .C(n4263), .Y(n2219) );
  AOI22X1 U4862 ( .A(\data_in<12> ), .B(n1119), .C(n4265), .D(n1254), .Y(n4266) );
  OAI21X1 U4863 ( .A(n1403), .B(n4267), .C(n4266), .Y(n2220) );
  AOI22X1 U4864 ( .A(\data_in<13> ), .B(n1119), .C(n4268), .D(n1254), .Y(n4269) );
  OAI21X1 U4865 ( .A(n1403), .B(n4270), .C(n4269), .Y(n2221) );
  AOI22X1 U4866 ( .A(\data_in<14> ), .B(n1119), .C(n4271), .D(n1254), .Y(n4272) );
  OAI21X1 U4867 ( .A(n1403), .B(n4273), .C(n4272), .Y(n2222) );
  AOI22X1 U4868 ( .A(\data_in<15> ), .B(n1119), .C(n4274), .D(n1254), .Y(n4275) );
  OAI21X1 U4869 ( .A(n1403), .B(n4276), .C(n4275), .Y(n2223) );
  AOI22X1 U4870 ( .A(\data_in<8> ), .B(n1120), .C(n4278), .D(n1256), .Y(n4279)
         );
  OAI21X1 U4871 ( .A(n1405), .B(n4280), .C(n4279), .Y(n2224) );
  AOI22X1 U4872 ( .A(\data_in<9> ), .B(n1120), .C(n4281), .D(n1256), .Y(n4282)
         );
  OAI21X1 U4873 ( .A(n1405), .B(n4283), .C(n4282), .Y(n2225) );
  AOI22X1 U4874 ( .A(\data_in<10> ), .B(n1120), .C(n4284), .D(n1256), .Y(n4285) );
  OAI21X1 U4875 ( .A(n1405), .B(n4286), .C(n4285), .Y(n2226) );
  AOI22X1 U4876 ( .A(\data_in<11> ), .B(n1120), .C(n4287), .D(n1256), .Y(n4288) );
  OAI21X1 U4877 ( .A(n1405), .B(n4289), .C(n4288), .Y(n2227) );
  AOI22X1 U4878 ( .A(\data_in<12> ), .B(n1120), .C(n4290), .D(n1256), .Y(n4291) );
  OAI21X1 U4879 ( .A(n1405), .B(n4292), .C(n4291), .Y(n2228) );
  AOI22X1 U4880 ( .A(\data_in<13> ), .B(n1120), .C(n4293), .D(n1256), .Y(n4294) );
  OAI21X1 U4881 ( .A(n1405), .B(n4295), .C(n4294), .Y(n2229) );
  AOI22X1 U4882 ( .A(\data_in<14> ), .B(n1120), .C(n4296), .D(n1256), .Y(n4297) );
  OAI21X1 U4883 ( .A(n1405), .B(n4298), .C(n4297), .Y(n2230) );
  AOI22X1 U4884 ( .A(\data_in<15> ), .B(n1120), .C(n4299), .D(n1256), .Y(n4300) );
  OAI21X1 U4885 ( .A(n1405), .B(n4301), .C(n4300), .Y(n2231) );
  AOI22X1 U4886 ( .A(\data_in<8> ), .B(n1121), .C(n4303), .D(n1258), .Y(n4304)
         );
  OAI21X1 U4887 ( .A(n1407), .B(n4305), .C(n4304), .Y(n2232) );
  AOI22X1 U4888 ( .A(\data_in<9> ), .B(n1121), .C(n4306), .D(n1258), .Y(n4307)
         );
  OAI21X1 U4889 ( .A(n1407), .B(n4308), .C(n4307), .Y(n2233) );
  AOI22X1 U4890 ( .A(\data_in<10> ), .B(n1121), .C(n4309), .D(n1258), .Y(n4310) );
  OAI21X1 U4891 ( .A(n1407), .B(n4311), .C(n4310), .Y(n2234) );
  AOI22X1 U4892 ( .A(\data_in<11> ), .B(n1121), .C(n4312), .D(n1258), .Y(n4313) );
  OAI21X1 U4893 ( .A(n1407), .B(n4314), .C(n4313), .Y(n2235) );
  AOI22X1 U4894 ( .A(\data_in<12> ), .B(n1121), .C(n4315), .D(n1258), .Y(n4316) );
  OAI21X1 U4895 ( .A(n1407), .B(n4317), .C(n4316), .Y(n2236) );
  AOI22X1 U4896 ( .A(\data_in<13> ), .B(n1121), .C(n4318), .D(n1258), .Y(n4319) );
  OAI21X1 U4897 ( .A(n1407), .B(n4320), .C(n4319), .Y(n2237) );
  AOI22X1 U4898 ( .A(\data_in<14> ), .B(n1121), .C(n4321), .D(n1258), .Y(n4322) );
  OAI21X1 U4899 ( .A(n1407), .B(n4323), .C(n4322), .Y(n2238) );
  AOI22X1 U4900 ( .A(\data_in<15> ), .B(n1121), .C(n4324), .D(n1258), .Y(n4325) );
  OAI21X1 U4901 ( .A(n1407), .B(n4326), .C(n4325), .Y(n2239) );
  AOI22X1 U4902 ( .A(\data_in<8> ), .B(n1122), .C(n4328), .D(n1260), .Y(n4329)
         );
  OAI21X1 U4903 ( .A(n1409), .B(n4330), .C(n4329), .Y(n2240) );
  AOI22X1 U4904 ( .A(\data_in<9> ), .B(n1122), .C(n4331), .D(n1260), .Y(n4332)
         );
  OAI21X1 U4905 ( .A(n1409), .B(n4333), .C(n4332), .Y(n2241) );
  AOI22X1 U4906 ( .A(\data_in<10> ), .B(n1122), .C(n4334), .D(n1260), .Y(n4335) );
  OAI21X1 U4907 ( .A(n1409), .B(n4336), .C(n4335), .Y(n2242) );
  AOI22X1 U4908 ( .A(\data_in<11> ), .B(n1122), .C(n4337), .D(n1260), .Y(n4338) );
  OAI21X1 U4909 ( .A(n1409), .B(n4339), .C(n4338), .Y(n2243) );
  AOI22X1 U4910 ( .A(\data_in<12> ), .B(n1122), .C(n4340), .D(n1260), .Y(n4341) );
  OAI21X1 U4911 ( .A(n1409), .B(n4342), .C(n4341), .Y(n2244) );
  AOI22X1 U4912 ( .A(\data_in<13> ), .B(n1122), .C(n4343), .D(n1260), .Y(n4344) );
  OAI21X1 U4913 ( .A(n1409), .B(n4345), .C(n4344), .Y(n2245) );
  AOI22X1 U4914 ( .A(\data_in<14> ), .B(n1122), .C(n4346), .D(n1260), .Y(n4347) );
  OAI21X1 U4915 ( .A(n1409), .B(n4348), .C(n4347), .Y(n2246) );
  AOI22X1 U4916 ( .A(\data_in<15> ), .B(n1122), .C(n4349), .D(n1260), .Y(n4350) );
  OAI21X1 U4917 ( .A(n1409), .B(n4351), .C(n4350), .Y(n2247) );
  AOI22X1 U4918 ( .A(\data_in<8> ), .B(n1123), .C(n4353), .D(n1262), .Y(n4354)
         );
  OAI21X1 U4919 ( .A(n1411), .B(n4355), .C(n4354), .Y(n2248) );
  AOI22X1 U4920 ( .A(\data_in<9> ), .B(n1123), .C(n4356), .D(n1262), .Y(n4357)
         );
  OAI21X1 U4921 ( .A(n1411), .B(n4358), .C(n4357), .Y(n2249) );
  AOI22X1 U4922 ( .A(\data_in<10> ), .B(n1123), .C(n4359), .D(n1262), .Y(n4360) );
  OAI21X1 U4923 ( .A(n1411), .B(n4361), .C(n4360), .Y(n2250) );
  AOI22X1 U4924 ( .A(\data_in<11> ), .B(n1123), .C(n4362), .D(n1262), .Y(n4363) );
  OAI21X1 U4925 ( .A(n1411), .B(n4364), .C(n4363), .Y(n2251) );
  AOI22X1 U4926 ( .A(\data_in<12> ), .B(n1123), .C(n4365), .D(n1262), .Y(n4366) );
  OAI21X1 U4927 ( .A(n1411), .B(n4367), .C(n4366), .Y(n2252) );
  AOI22X1 U4928 ( .A(\data_in<13> ), .B(n1123), .C(n4368), .D(n1262), .Y(n4369) );
  OAI21X1 U4929 ( .A(n1411), .B(n4370), .C(n4369), .Y(n2253) );
  AOI22X1 U4930 ( .A(\data_in<14> ), .B(n1123), .C(n4371), .D(n1262), .Y(n4372) );
  OAI21X1 U4931 ( .A(n1411), .B(n4373), .C(n4372), .Y(n2254) );
  AOI22X1 U4932 ( .A(\data_in<15> ), .B(n1123), .C(n4374), .D(n1262), .Y(n4375) );
  OAI21X1 U4933 ( .A(n1411), .B(n4376), .C(n4375), .Y(n2255) );
  AOI22X1 U4934 ( .A(\data_in<8> ), .B(n1124), .C(n4378), .D(n1264), .Y(n4379)
         );
  OAI21X1 U4935 ( .A(n1413), .B(n4380), .C(n4379), .Y(n2256) );
  AOI22X1 U4936 ( .A(\data_in<9> ), .B(n1124), .C(n4381), .D(n1264), .Y(n4382)
         );
  OAI21X1 U4937 ( .A(n1413), .B(n4383), .C(n4382), .Y(n2257) );
  AOI22X1 U4938 ( .A(\data_in<10> ), .B(n1124), .C(n4384), .D(n1264), .Y(n4385) );
  OAI21X1 U4939 ( .A(n1413), .B(n4386), .C(n4385), .Y(n2258) );
  AOI22X1 U4940 ( .A(\data_in<11> ), .B(n1124), .C(n4387), .D(n1264), .Y(n4388) );
  OAI21X1 U4941 ( .A(n1413), .B(n4389), .C(n4388), .Y(n2259) );
  AOI22X1 U4942 ( .A(\data_in<12> ), .B(n1124), .C(n4390), .D(n1264), .Y(n4391) );
  OAI21X1 U4943 ( .A(n1413), .B(n4392), .C(n4391), .Y(n2260) );
  AOI22X1 U4944 ( .A(\data_in<13> ), .B(n1124), .C(n4393), .D(n1264), .Y(n4394) );
  OAI21X1 U4945 ( .A(n1413), .B(n4395), .C(n4394), .Y(n2261) );
  AOI22X1 U4946 ( .A(\data_in<14> ), .B(n1124), .C(n4396), .D(n1264), .Y(n4397) );
  OAI21X1 U4947 ( .A(n1413), .B(n4398), .C(n4397), .Y(n2262) );
  AOI22X1 U4948 ( .A(\data_in<15> ), .B(n1124), .C(n4399), .D(n1264), .Y(n4400) );
  OAI21X1 U4949 ( .A(n1413), .B(n4401), .C(n4400), .Y(n2263) );
  AOI22X1 U4950 ( .A(\data_in<8> ), .B(n1125), .C(n4403), .D(n1266), .Y(n4404)
         );
  OAI21X1 U4951 ( .A(n1415), .B(n4405), .C(n4404), .Y(n2264) );
  AOI22X1 U4952 ( .A(\data_in<9> ), .B(n1125), .C(n4406), .D(n1266), .Y(n4407)
         );
  OAI21X1 U4953 ( .A(n1415), .B(n4408), .C(n4407), .Y(n2265) );
  AOI22X1 U4954 ( .A(\data_in<10> ), .B(n1125), .C(n4409), .D(n1266), .Y(n4410) );
  OAI21X1 U4955 ( .A(n1415), .B(n4411), .C(n4410), .Y(n2266) );
  AOI22X1 U4956 ( .A(\data_in<11> ), .B(n1125), .C(n4412), .D(n1266), .Y(n4413) );
  OAI21X1 U4957 ( .A(n1415), .B(n4414), .C(n4413), .Y(n2267) );
  AOI22X1 U4958 ( .A(\data_in<12> ), .B(n1125), .C(n4415), .D(n1266), .Y(n4416) );
  OAI21X1 U4959 ( .A(n1415), .B(n4417), .C(n4416), .Y(n2268) );
  AOI22X1 U4960 ( .A(\data_in<13> ), .B(n1125), .C(n4418), .D(n1266), .Y(n4419) );
  OAI21X1 U4961 ( .A(n1415), .B(n4420), .C(n4419), .Y(n2269) );
  AOI22X1 U4962 ( .A(\data_in<14> ), .B(n1125), .C(n4421), .D(n1266), .Y(n4422) );
  OAI21X1 U4963 ( .A(n1415), .B(n4423), .C(n4422), .Y(n2270) );
  AOI22X1 U4964 ( .A(\data_in<15> ), .B(n1125), .C(n4424), .D(n1266), .Y(n4425) );
  OAI21X1 U4965 ( .A(n1415), .B(n4426), .C(n4425), .Y(n2271) );
  AOI22X1 U4966 ( .A(\data_in<8> ), .B(n1126), .C(n4427), .D(n1268), .Y(n4428)
         );
  OAI21X1 U4967 ( .A(n1417), .B(n4429), .C(n4428), .Y(n2272) );
  AOI22X1 U4968 ( .A(\data_in<9> ), .B(n1126), .C(n4430), .D(n1268), .Y(n4431)
         );
  OAI21X1 U4969 ( .A(n1417), .B(n4432), .C(n4431), .Y(n2273) );
  AOI22X1 U4970 ( .A(\data_in<10> ), .B(n1126), .C(n4433), .D(n1268), .Y(n4434) );
  OAI21X1 U4971 ( .A(n1417), .B(n4435), .C(n4434), .Y(n2274) );
  AOI22X1 U4972 ( .A(\data_in<11> ), .B(n1126), .C(n4436), .D(n1268), .Y(n4437) );
  OAI21X1 U4973 ( .A(n1417), .B(n4438), .C(n4437), .Y(n2275) );
  AOI22X1 U4974 ( .A(\data_in<12> ), .B(n1126), .C(n4439), .D(n1268), .Y(n4440) );
  OAI21X1 U4975 ( .A(n1417), .B(n4441), .C(n4440), .Y(n2276) );
  AOI22X1 U4976 ( .A(\data_in<13> ), .B(n1126), .C(n4442), .D(n1268), .Y(n4443) );
  OAI21X1 U4977 ( .A(n1417), .B(n4444), .C(n4443), .Y(n2277) );
  AOI22X1 U4978 ( .A(\data_in<14> ), .B(n1126), .C(n4445), .D(n1268), .Y(n4446) );
  OAI21X1 U4979 ( .A(n1417), .B(n4447), .C(n4446), .Y(n2278) );
  AOI22X1 U4980 ( .A(\data_in<15> ), .B(n1126), .C(n4448), .D(n1268), .Y(n4449) );
  OAI21X1 U4981 ( .A(n1417), .B(n4450), .C(n4449), .Y(n2279) );
  AOI22X1 U4982 ( .A(\data_in<8> ), .B(n1127), .C(n4452), .D(n1270), .Y(n4453)
         );
  OAI21X1 U4983 ( .A(n1419), .B(n4454), .C(n4453), .Y(n2280) );
  AOI22X1 U4984 ( .A(\data_in<9> ), .B(n1127), .C(n4455), .D(n1270), .Y(n4456)
         );
  OAI21X1 U4985 ( .A(n1419), .B(n4457), .C(n4456), .Y(n2281) );
  AOI22X1 U4986 ( .A(\data_in<10> ), .B(n1127), .C(n4458), .D(n1270), .Y(n4459) );
  OAI21X1 U4987 ( .A(n1419), .B(n4460), .C(n4459), .Y(n2282) );
  AOI22X1 U4988 ( .A(\data_in<11> ), .B(n1127), .C(n4461), .D(n1270), .Y(n4462) );
  OAI21X1 U4989 ( .A(n1419), .B(n4463), .C(n4462), .Y(n2283) );
  AOI22X1 U4990 ( .A(\data_in<12> ), .B(n1127), .C(n4464), .D(n1270), .Y(n4465) );
  OAI21X1 U4991 ( .A(n1419), .B(n4466), .C(n4465), .Y(n2284) );
  AOI22X1 U4992 ( .A(\data_in<13> ), .B(n1127), .C(n4467), .D(n1270), .Y(n4468) );
  OAI21X1 U4993 ( .A(n1419), .B(n4469), .C(n4468), .Y(n2285) );
  AOI22X1 U4994 ( .A(\data_in<14> ), .B(n1127), .C(n4470), .D(n1270), .Y(n4471) );
  OAI21X1 U4995 ( .A(n1419), .B(n4472), .C(n4471), .Y(n2286) );
  AOI22X1 U4996 ( .A(\data_in<15> ), .B(n1127), .C(n4473), .D(n1270), .Y(n4474) );
  OAI21X1 U4997 ( .A(n1419), .B(n4475), .C(n4474), .Y(n2287) );
  AOI22X1 U4998 ( .A(\data_in<8> ), .B(n1128), .C(n4477), .D(n1272), .Y(n4478)
         );
  OAI21X1 U4999 ( .A(n1421), .B(n4479), .C(n4478), .Y(n2288) );
  AOI22X1 U5000 ( .A(\data_in<9> ), .B(n1128), .C(n4480), .D(n1272), .Y(n4481)
         );
  OAI21X1 U5001 ( .A(n1421), .B(n4482), .C(n4481), .Y(n2289) );
  AOI22X1 U5002 ( .A(\data_in<10> ), .B(n1128), .C(n4483), .D(n1272), .Y(n4484) );
  OAI21X1 U5003 ( .A(n1421), .B(n4485), .C(n4484), .Y(n2290) );
  AOI22X1 U5004 ( .A(\data_in<11> ), .B(n1128), .C(n4486), .D(n1272), .Y(n4487) );
  OAI21X1 U5005 ( .A(n1421), .B(n4488), .C(n4487), .Y(n2291) );
  AOI22X1 U5006 ( .A(\data_in<12> ), .B(n1128), .C(n4489), .D(n1272), .Y(n4490) );
  OAI21X1 U5007 ( .A(n1421), .B(n4491), .C(n4490), .Y(n2292) );
  AOI22X1 U5008 ( .A(\data_in<13> ), .B(n1128), .C(n4492), .D(n1272), .Y(n4493) );
  OAI21X1 U5009 ( .A(n1421), .B(n4494), .C(n4493), .Y(n2293) );
  AOI22X1 U5010 ( .A(\data_in<14> ), .B(n1128), .C(n4495), .D(n1272), .Y(n4496) );
  OAI21X1 U5011 ( .A(n1421), .B(n4497), .C(n4496), .Y(n2294) );
  AOI22X1 U5012 ( .A(\data_in<15> ), .B(n1128), .C(n4498), .D(n1272), .Y(n4499) );
  OAI21X1 U5013 ( .A(n1421), .B(n4500), .C(n4499), .Y(n2295) );
  AOI22X1 U5014 ( .A(\data_in<8> ), .B(n1129), .C(n4502), .D(n1274), .Y(n4503)
         );
  OAI21X1 U5015 ( .A(n1423), .B(n4504), .C(n4503), .Y(n2296) );
  AOI22X1 U5016 ( .A(\data_in<9> ), .B(n1129), .C(n4505), .D(n1274), .Y(n4506)
         );
  OAI21X1 U5017 ( .A(n1423), .B(n4507), .C(n4506), .Y(n2297) );
  AOI22X1 U5018 ( .A(\data_in<10> ), .B(n1129), .C(n4508), .D(n1274), .Y(n4509) );
  OAI21X1 U5019 ( .A(n1423), .B(n4510), .C(n4509), .Y(n2298) );
  AOI22X1 U5020 ( .A(\data_in<11> ), .B(n1129), .C(n4511), .D(n1274), .Y(n4512) );
  OAI21X1 U5021 ( .A(n1423), .B(n4513), .C(n4512), .Y(n2299) );
  AOI22X1 U5022 ( .A(\data_in<12> ), .B(n1129), .C(n4514), .D(n1274), .Y(n4515) );
  OAI21X1 U5023 ( .A(n1423), .B(n4516), .C(n4515), .Y(n2300) );
  AOI22X1 U5024 ( .A(\data_in<13> ), .B(n1129), .C(n4517), .D(n1274), .Y(n4518) );
  OAI21X1 U5025 ( .A(n1423), .B(n4519), .C(n4518), .Y(n2301) );
  AOI22X1 U5026 ( .A(\data_in<14> ), .B(n1129), .C(n4520), .D(n1274), .Y(n4521) );
  OAI21X1 U5027 ( .A(n1423), .B(n4522), .C(n4521), .Y(n2302) );
  AOI22X1 U5028 ( .A(\data_in<15> ), .B(n1129), .C(n4523), .D(n1274), .Y(n4524) );
  OAI21X1 U5029 ( .A(n1423), .B(n4525), .C(n4524), .Y(n2303) );
  AOI22X1 U5030 ( .A(\data_in<8> ), .B(n1130), .C(n4527), .D(n1276), .Y(n4528)
         );
  OAI21X1 U5031 ( .A(n1425), .B(n4529), .C(n4528), .Y(n2304) );
  AOI22X1 U5032 ( .A(\data_in<9> ), .B(n1130), .C(n4530), .D(n1276), .Y(n4531)
         );
  OAI21X1 U5033 ( .A(n1425), .B(n4532), .C(n4531), .Y(n2305) );
  AOI22X1 U5034 ( .A(\data_in<10> ), .B(n1130), .C(n4533), .D(n1276), .Y(n4534) );
  OAI21X1 U5035 ( .A(n1425), .B(n4535), .C(n4534), .Y(n2306) );
  AOI22X1 U5036 ( .A(\data_in<11> ), .B(n1130), .C(n4536), .D(n1276), .Y(n4537) );
  OAI21X1 U5037 ( .A(n1425), .B(n4538), .C(n4537), .Y(n2307) );
  AOI22X1 U5038 ( .A(\data_in<12> ), .B(n1130), .C(n4539), .D(n1276), .Y(n4540) );
  OAI21X1 U5039 ( .A(n1425), .B(n4541), .C(n4540), .Y(n2308) );
  AOI22X1 U5040 ( .A(\data_in<13> ), .B(n1130), .C(n4542), .D(n1276), .Y(n4543) );
  OAI21X1 U5041 ( .A(n1425), .B(n4544), .C(n4543), .Y(n2309) );
  AOI22X1 U5042 ( .A(\data_in<14> ), .B(n1130), .C(n4545), .D(n1276), .Y(n4546) );
  OAI21X1 U5043 ( .A(n1425), .B(n4547), .C(n4546), .Y(n2310) );
  AOI22X1 U5044 ( .A(\data_in<15> ), .B(n1130), .C(n4548), .D(n1276), .Y(n4549) );
  OAI21X1 U5045 ( .A(n1425), .B(n4550), .C(n4549), .Y(n2311) );
  OAI21X1 U5046 ( .A(n4551), .B(n1295), .C(n1284), .Y(n4574) );
  NOR2X1 U5047 ( .A(n4574), .B(n2711), .Y(n4553) );
  AOI21X1 U5048 ( .A(\data_in<8> ), .B(n1131), .C(n4553), .Y(n4554) );
  OAI21X1 U5049 ( .A(n1427), .B(n4555), .C(n810), .Y(n2312) );
  NOR2X1 U5050 ( .A(n4574), .B(n2768), .Y(n4556) );
  AOI21X1 U5051 ( .A(\data_in<9> ), .B(n1131), .C(n4556), .Y(n4557) );
  OAI21X1 U5052 ( .A(n1427), .B(n4558), .C(n811), .Y(n2313) );
  NOR2X1 U5053 ( .A(n4574), .B(n4596), .Y(n4559) );
  AOI21X1 U5054 ( .A(\data_in<10> ), .B(n1131), .C(n4559), .Y(n4560) );
  OAI21X1 U5055 ( .A(n1427), .B(n4561), .C(n812), .Y(n2314) );
  NOR2X1 U5056 ( .A(n4574), .B(n4595), .Y(n4562) );
  AOI21X1 U5057 ( .A(\data_in<11> ), .B(n1131), .C(n4562), .Y(n4563) );
  OAI21X1 U5058 ( .A(n1427), .B(n4564), .C(n813), .Y(n2315) );
  NOR2X1 U5059 ( .A(n4574), .B(n4594), .Y(n4565) );
  AOI21X1 U5060 ( .A(\data_in<12> ), .B(n1131), .C(n4565), .Y(n4566) );
  OAI21X1 U5061 ( .A(n1427), .B(n4567), .C(n814), .Y(n2316) );
  NOR2X1 U5062 ( .A(n4574), .B(n4593), .Y(n4568) );
  AOI21X1 U5063 ( .A(\data_in<13> ), .B(n1131), .C(n4568), .Y(n4569) );
  OAI21X1 U5064 ( .A(n1427), .B(n4570), .C(n815), .Y(n2317) );
  NOR2X1 U5065 ( .A(n4574), .B(n4592), .Y(n4571) );
  AOI21X1 U5066 ( .A(\data_in<14> ), .B(n1131), .C(n4571), .Y(n4572) );
  OAI21X1 U5067 ( .A(n1427), .B(n4573), .C(n816), .Y(n2318) );
  NOR2X1 U5068 ( .A(n4574), .B(n2905), .Y(n4575) );
  AOI21X1 U5069 ( .A(\data_in<15> ), .B(n1131), .C(n4575), .Y(n4576) );
  OAI21X1 U5070 ( .A(n1427), .B(n4577), .C(n817), .Y(n2319) );
  MUX2X1 U5071 ( .B(n2700), .A(n4578), .S(n1283), .Y(n2320) );
  MUX2X1 U5072 ( .B(n2758), .A(n4579), .S(n1283), .Y(n2321) );
  MUX2X1 U5073 ( .B(n4591), .A(n4580), .S(n1283), .Y(n2322) );
  MUX2X1 U5074 ( .B(n4590), .A(n4581), .S(n1283), .Y(n2323) );
  MUX2X1 U5075 ( .B(n4589), .A(n4582), .S(n1283), .Y(n2324) );
  MUX2X1 U5076 ( .B(n4588), .A(n4583), .S(n1283), .Y(n2325) );
  MUX2X1 U5077 ( .B(n4587), .A(n4584), .S(n1283), .Y(n2326) );
  MUX2X1 U5078 ( .B(n2894), .A(n4585), .S(n1283), .Y(n2327) );
endmodule


module cla16_2 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14;

  cla4_11 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_10 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n14), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_9 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n13), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_8 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n12), .S({\S<15> , \S<14> , \S<13> , \S<12> }), .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  INVX1 U1 ( .A(Cin), .Y(n4) );
  INVX1 U2 ( .A(\G<0> ), .Y(n3) );
  INVX1 U3 ( .A(\G<1> ), .Y(n6) );
  INVX1 U4 ( .A(\G<3> ), .Y(n10) );
  AND2X2 U5 ( .A(\P<3> ), .B(n12), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  INVX1 U7 ( .A(n9), .Y(n12) );
  INVX1 U8 ( .A(\P<1> ), .Y(n7) );
  INVX1 U9 ( .A(\P<0> ), .Y(n5) );
  OAI21X1 U10 ( .A(n5), .B(n4), .C(n3), .Y(n14) );
  INVX2 U11 ( .A(n14), .Y(n8) );
  OAI21X1 U12 ( .A(n8), .B(n7), .C(n6), .Y(n13) );
  AOI21X1 U13 ( .A(\P<2> ), .B(n13), .C(\G<2> ), .Y(n9) );
  NAND2X1 U14 ( .A(n10), .B(n2), .Y(Cout) );
endmodule


module rf ( .read1data({\read1data<15> , \read1data<14> , \read1data<13> , 
        \read1data<12> , \read1data<11> , \read1data<10> , \read1data<9> , 
        \read1data<8> , \read1data<7> , \read1data<6> , \read1data<5> , 
        \read1data<4> , \read1data<3> , \read1data<2> , \read1data<1> , 
        \read1data<0> }), .read2data({\read2data<15> , \read2data<14> , 
        \read2data<13> , \read2data<12> , \read2data<11> , \read2data<10> , 
        \read2data<9> , \read2data<8> , \read2data<7> , \read2data<6> , 
        \read2data<5> , \read2data<4> , \read2data<3> , \read2data<2> , 
        \read2data<1> , \read2data<0> }), err, clk, rst, .read1regsel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .read2regsel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .writeregsel({
        \writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   \rf_wr_en<7> , \rf_wr_en<6> , \rf_wr_en<5> , \rf_wr_en<4> ,
         \rf_wr_en<3> , \rf_wr_en<2> , \rf_wr_en<1> , \rf_wr_en<0> ,
         \write_en<7> , \write_en<6> , \write_en<5> , \write_en<4> ,
         \write_en<3> , \write_en<2> , \write_en<1> , \write_en<0> ,
         \reg_in<127> , \reg_in<126> , \reg_in<125> , \reg_in<124> ,
         \reg_in<123> , \reg_in<122> , \reg_in<121> , \reg_in<120> ,
         \reg_in<119> , \reg_in<118> , \reg_in<117> , \reg_in<116> ,
         \reg_in<115> , \reg_in<114> , \reg_in<113> , \reg_in<112> ,
         \reg_in<111> , \reg_in<110> , \reg_in<109> , \reg_in<108> ,
         \reg_in<107> , \reg_in<106> , \reg_in<105> , \reg_in<104> ,
         \reg_in<103> , \reg_in<102> , \reg_in<101> , \reg_in<100> ,
         \reg_in<99> , \reg_in<98> , \reg_in<97> , \reg_in<96> , \reg_in<95> ,
         \reg_in<94> , \reg_in<93> , \reg_in<92> , \reg_in<91> , \reg_in<90> ,
         \reg_in<89> , \reg_in<88> , \reg_in<87> , \reg_in<86> , \reg_in<85> ,
         \reg_in<84> , \reg_in<83> , \reg_in<82> , \reg_in<81> , \reg_in<80> ,
         \reg_in<79> , \reg_in<78> , \reg_in<77> , \reg_in<76> , \reg_in<75> ,
         \reg_in<74> , \reg_in<73> , \reg_in<72> , \reg_in<71> , \reg_in<70> ,
         \reg_in<69> , \reg_in<68> , \reg_in<67> , \reg_in<66> , \reg_in<65> ,
         \reg_in<64> , \reg_in<63> , \reg_in<62> , \reg_in<61> , \reg_in<60> ,
         \reg_in<59> , \reg_in<58> , \reg_in<57> , \reg_in<56> , \reg_in<55> ,
         \reg_in<54> , \reg_in<53> , \reg_in<52> , \reg_in<51> , \reg_in<50> ,
         \reg_in<49> , \reg_in<48> , \reg_in<47> , \reg_in<46> , \reg_in<45> ,
         \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> ,
         \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> ,
         \reg_in<34> , \reg_in<33> , \reg_in<32> , \reg_in<31> , \reg_in<30> ,
         \reg_in<29> , \reg_in<28> , \reg_in<27> , \reg_in<26> , \reg_in<25> ,
         \reg_in<24> , \reg_in<23> , \reg_in<22> , \reg_in<21> , \reg_in<20> ,
         \reg_in<19> , \reg_in<18> , \reg_in<17> , \reg_in<16> , \reg_in<15> ,
         \reg_in<14> , \reg_in<13> , \reg_in<12> , \reg_in<11> , \reg_in<10> ,
         \reg_in<9> , \reg_in<8> , \reg_in<7> , \reg_in<6> , \reg_in<5> ,
         \reg_in<4> , \reg_in<3> , \reg_in<2> , \reg_in<1> , \reg_in<0> ,
         \reg_out<127> , \reg_out<126> , \reg_out<125> , \reg_out<124> ,
         \reg_out<123> , \reg_out<122> , \reg_out<121> , \reg_out<120> ,
         \reg_out<119> , \reg_out<118> , \reg_out<117> , \reg_out<116> ,
         \reg_out<115> , \reg_out<114> , \reg_out<113> , \reg_out<112> ,
         \reg_out<111> , \reg_out<110> , \reg_out<109> , \reg_out<108> ,
         \reg_out<107> , \reg_out<106> , \reg_out<105> , \reg_out<104> ,
         \reg_out<103> , \reg_out<102> , \reg_out<101> , \reg_out<100> ,
         \reg_out<99> , \reg_out<98> , \reg_out<97> , \reg_out<96> ,
         \reg_out<95> , \reg_out<94> , \reg_out<93> , \reg_out<92> ,
         \reg_out<91> , \reg_out<90> , \reg_out<89> , \reg_out<88> ,
         \reg_out<87> , \reg_out<86> , \reg_out<85> , \reg_out<84> ,
         \reg_out<83> , \reg_out<82> , \reg_out<81> , \reg_out<80> ,
         \reg_out<79> , \reg_out<78> , \reg_out<77> , \reg_out<76> ,
         \reg_out<75> , \reg_out<74> , \reg_out<73> , \reg_out<72> ,
         \reg_out<71> , \reg_out<70> , \reg_out<69> , \reg_out<68> ,
         \reg_out<67> , \reg_out<66> , \reg_out<65> , \reg_out<64> ,
         \reg_out<63> , \reg_out<62> , \reg_out<61> , \reg_out<60> ,
         \reg_out<59> , \reg_out<58> , \reg_out<57> , \reg_out<56> ,
         \reg_out<55> , \reg_out<54> , \reg_out<53> , \reg_out<52> ,
         \reg_out<51> , \reg_out<50> , \reg_out<49> , \reg_out<48> ,
         \reg_out<47> , \reg_out<46> , \reg_out<45> , \reg_out<44> ,
         \reg_out<43> , \reg_out<42> , \reg_out<41> , \reg_out<40> ,
         \reg_out<39> , \reg_out<38> , \reg_out<37> , \reg_out<36> ,
         \reg_out<35> , \reg_out<34> , \reg_out<33> , \reg_out<32> ,
         \reg_out<31> , \reg_out<30> , \reg_out<29> , \reg_out<28> ,
         \reg_out<27> , \reg_out<26> , \reg_out<25> , \reg_out<24> ,
         \reg_out<23> , \reg_out<22> , \reg_out<21> , \reg_out<20> ,
         \reg_out<19> , \reg_out<18> , \reg_out<17> , \reg_out<16> ,
         \reg_out<15> , \reg_out<14> , \reg_out<13> , \reg_out<12> ,
         \reg_out<11> , \reg_out<10> , \reg_out<9> , \reg_out<8> ,
         \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , \reg_out<3> ,
         \reg_out<2> , \reg_out<1> , \reg_out<0> , n1, n2, n3, n4;
  assign err = 1'b0;

  AND2X2 U2 ( .A(\write_en<7> ), .B(write), .Y(\rf_wr_en<7> ) );
  AND2X2 U3 ( .A(\write_en<6> ), .B(write), .Y(\rf_wr_en<6> ) );
  AND2X2 U4 ( .A(\write_en<5> ), .B(write), .Y(\rf_wr_en<5> ) );
  AND2X2 U5 ( .A(\write_en<4> ), .B(write), .Y(\rf_wr_en<4> ) );
  AND2X2 U6 ( .A(\write_en<3> ), .B(write), .Y(\rf_wr_en<3> ) );
  AND2X2 U7 ( .A(\write_en<2> ), .B(write), .Y(\rf_wr_en<2> ) );
  AND2X2 U8 ( .A(\write_en<1> ), .B(write), .Y(\rf_wr_en<1> ) );
  AND2X2 U9 ( .A(\write_en<0> ), .B(write), .Y(\rf_wr_en<0> ) );
  register16_0 \registers[0]  ( .d({\reg_in<15> , \reg_in<14> , \reg_in<13> , 
        \reg_in<12> , \reg_in<11> , \reg_in<10> , \reg_in<9> , \reg_in<8> , 
        \reg_in<7> , \reg_in<6> , \reg_in<5> , \reg_in<4> , \reg_in<3> , 
        \reg_in<2> , \reg_in<1> , \reg_in<0> }), .clk(clk), .wr_en(
        \rf_wr_en<0> ), .rst(n4), .q({\reg_out<15> , \reg_out<14> , 
        \reg_out<13> , \reg_out<12> , \reg_out<11> , \reg_out<10> , 
        \reg_out<9> , \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , 
        \reg_out<4> , \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> })
         );
  register16_1 \registers[1]  ( .d({\reg_in<31> , \reg_in<30> , \reg_in<29> , 
        \reg_in<28> , \reg_in<27> , \reg_in<26> , \reg_in<25> , \reg_in<24> , 
        \reg_in<23> , \reg_in<22> , \reg_in<21> , \reg_in<20> , \reg_in<19> , 
        \reg_in<18> , \reg_in<17> , \reg_in<16> }), .clk(clk), .wr_en(
        \rf_wr_en<1> ), .rst(n3), .q({\reg_out<31> , \reg_out<30> , 
        \reg_out<29> , \reg_out<28> , \reg_out<27> , \reg_out<26> , 
        \reg_out<25> , \reg_out<24> , \reg_out<23> , \reg_out<22> , 
        \reg_out<21> , \reg_out<20> , \reg_out<19> , \reg_out<18> , 
        \reg_out<17> , \reg_out<16> }) );
  register16_2 \registers[2]  ( .d({\reg_in<47> , \reg_in<46> , \reg_in<45> , 
        \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> , 
        \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> , 
        \reg_in<34> , \reg_in<33> , \reg_in<32> }), .clk(clk), .wr_en(
        \rf_wr_en<2> ), .rst(n3), .q({\reg_out<47> , \reg_out<46> , 
        \reg_out<45> , \reg_out<44> , \reg_out<43> , \reg_out<42> , 
        \reg_out<41> , \reg_out<40> , \reg_out<39> , \reg_out<38> , 
        \reg_out<37> , \reg_out<36> , \reg_out<35> , \reg_out<34> , 
        \reg_out<33> , \reg_out<32> }) );
  register16_3 \registers[3]  ( .d({\reg_in<63> , \reg_in<62> , \reg_in<61> , 
        \reg_in<60> , \reg_in<59> , \reg_in<58> , \reg_in<57> , \reg_in<56> , 
        \reg_in<55> , \reg_in<54> , \reg_in<53> , \reg_in<52> , \reg_in<51> , 
        \reg_in<50> , \reg_in<49> , \reg_in<48> }), .clk(clk), .wr_en(
        \rf_wr_en<3> ), .rst(n3), .q({\reg_out<63> , \reg_out<62> , 
        \reg_out<61> , \reg_out<60> , \reg_out<59> , \reg_out<58> , 
        \reg_out<57> , \reg_out<56> , \reg_out<55> , \reg_out<54> , 
        \reg_out<53> , \reg_out<52> , \reg_out<51> , \reg_out<50> , 
        \reg_out<49> , \reg_out<48> }) );
  register16_4 \registers[4]  ( .d({\reg_in<79> , \reg_in<78> , \reg_in<77> , 
        \reg_in<76> , \reg_in<75> , \reg_in<74> , \reg_in<73> , \reg_in<72> , 
        \reg_in<71> , \reg_in<70> , \reg_in<69> , \reg_in<68> , \reg_in<67> , 
        \reg_in<66> , \reg_in<65> , \reg_in<64> }), .clk(clk), .wr_en(
        \rf_wr_en<4> ), .rst(n3), .q({\reg_out<79> , \reg_out<78> , 
        \reg_out<77> , \reg_out<76> , \reg_out<75> , \reg_out<74> , 
        \reg_out<73> , \reg_out<72> , \reg_out<71> , \reg_out<70> , 
        \reg_out<69> , \reg_out<68> , \reg_out<67> , \reg_out<66> , 
        \reg_out<65> , \reg_out<64> }) );
  register16_5 \registers[5]  ( .d({\reg_in<95> , \reg_in<94> , \reg_in<93> , 
        \reg_in<92> , \reg_in<91> , \reg_in<90> , \reg_in<89> , \reg_in<88> , 
        \reg_in<87> , \reg_in<86> , \reg_in<85> , \reg_in<84> , \reg_in<83> , 
        \reg_in<82> , \reg_in<81> , \reg_in<80> }), .clk(clk), .wr_en(
        \rf_wr_en<5> ), .rst(n4), .q({\reg_out<95> , \reg_out<94> , 
        \reg_out<93> , \reg_out<92> , \reg_out<91> , \reg_out<90> , 
        \reg_out<89> , \reg_out<88> , \reg_out<87> , \reg_out<86> , 
        \reg_out<85> , \reg_out<84> , \reg_out<83> , \reg_out<82> , 
        \reg_out<81> , \reg_out<80> }) );
  register16_6 \registers[6]  ( .d({\reg_in<111> , \reg_in<110> , 
        \reg_in<109> , \reg_in<108> , \reg_in<107> , \reg_in<106> , 
        \reg_in<105> , \reg_in<104> , \reg_in<103> , \reg_in<102> , 
        \reg_in<101> , \reg_in<100> , \reg_in<99> , \reg_in<98> , \reg_in<97> , 
        \reg_in<96> }), .clk(clk), .wr_en(\rf_wr_en<6> ), .rst(n4), .q({
        \reg_out<111> , \reg_out<110> , \reg_out<109> , \reg_out<108> , 
        \reg_out<107> , \reg_out<106> , \reg_out<105> , \reg_out<104> , 
        \reg_out<103> , \reg_out<102> , \reg_out<101> , \reg_out<100> , 
        \reg_out<99> , \reg_out<98> , \reg_out<97> , \reg_out<96> }) );
  register16_7 \registers[7]  ( .d({\reg_in<127> , \reg_in<126> , 
        \reg_in<125> , \reg_in<124> , \reg_in<123> , \reg_in<122> , 
        \reg_in<121> , \reg_in<120> , \reg_in<119> , \reg_in<118> , 
        \reg_in<117> , \reg_in<116> , \reg_in<115> , \reg_in<114> , 
        \reg_in<113> , \reg_in<112> }), .clk(clk), .wr_en(\rf_wr_en<7> ), 
        .rst(n4), .q({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> }) );
  decoder3to8 wr_dec ( .In({\writeregsel<2> , \writeregsel<1> , n1}), .Out({
        \write_en<7> , \write_en<6> , \write_en<5> , \write_en<4> , 
        \write_en<3> , \write_en<2> , \write_en<1> , \write_en<0> }) );
  mux8to1_16_1 read1_mux ( .In({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> , \reg_out<111> , \reg_out<110> , \reg_out<109> , 
        \reg_out<108> , \reg_out<107> , \reg_out<106> , \reg_out<105> , 
        \reg_out<104> , \reg_out<103> , \reg_out<102> , \reg_out<101> , 
        \reg_out<100> , \reg_out<99> , \reg_out<98> , \reg_out<97> , 
        \reg_out<96> , \reg_out<95> , \reg_out<94> , \reg_out<93> , 
        \reg_out<92> , \reg_out<91> , \reg_out<90> , \reg_out<89> , 
        \reg_out<88> , \reg_out<87> , \reg_out<86> , \reg_out<85> , 
        \reg_out<84> , \reg_out<83> , \reg_out<82> , \reg_out<81> , 
        \reg_out<80> , \reg_out<79> , \reg_out<78> , \reg_out<77> , 
        \reg_out<76> , \reg_out<75> , \reg_out<74> , \reg_out<73> , 
        \reg_out<72> , \reg_out<71> , \reg_out<70> , \reg_out<69> , 
        \reg_out<68> , \reg_out<67> , \reg_out<66> , \reg_out<65> , 
        \reg_out<64> , \reg_out<63> , \reg_out<62> , \reg_out<61> , 
        \reg_out<60> , \reg_out<59> , \reg_out<58> , \reg_out<57> , 
        \reg_out<56> , \reg_out<55> , \reg_out<54> , \reg_out<53> , 
        \reg_out<52> , \reg_out<51> , \reg_out<50> , \reg_out<49> , 
        \reg_out<48> , \reg_out<47> , \reg_out<46> , \reg_out<45> , 
        \reg_out<44> , \reg_out<43> , \reg_out<42> , \reg_out<41> , 
        \reg_out<40> , \reg_out<39> , \reg_out<38> , \reg_out<37> , 
        \reg_out<36> , \reg_out<35> , \reg_out<34> , \reg_out<33> , 
        \reg_out<32> , \reg_out<31> , \reg_out<30> , \reg_out<29> , 
        \reg_out<28> , \reg_out<27> , \reg_out<26> , \reg_out<25> , 
        \reg_out<24> , \reg_out<23> , \reg_out<22> , \reg_out<21> , 
        \reg_out<20> , \reg_out<19> , \reg_out<18> , \reg_out<17> , 
        \reg_out<16> , \reg_out<15> , \reg_out<14> , \reg_out<13> , 
        \reg_out<12> , \reg_out<11> , \reg_out<10> , \reg_out<9> , 
        \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , 
        \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> }), .Sel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .Out({
        \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> , 
        \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> , 
        \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> , 
        \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> }) );
  mux8to1_16_0 read2_mux ( .In({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> , \reg_out<111> , \reg_out<110> , \reg_out<109> , 
        \reg_out<108> , \reg_out<107> , \reg_out<106> , \reg_out<105> , 
        \reg_out<104> , \reg_out<103> , \reg_out<102> , \reg_out<101> , 
        \reg_out<100> , \reg_out<99> , \reg_out<98> , \reg_out<97> , 
        \reg_out<96> , \reg_out<95> , \reg_out<94> , \reg_out<93> , 
        \reg_out<92> , \reg_out<91> , \reg_out<90> , \reg_out<89> , 
        \reg_out<88> , \reg_out<87> , \reg_out<86> , \reg_out<85> , 
        \reg_out<84> , \reg_out<83> , \reg_out<82> , \reg_out<81> , 
        \reg_out<80> , \reg_out<79> , \reg_out<78> , \reg_out<77> , 
        \reg_out<76> , \reg_out<75> , \reg_out<74> , \reg_out<73> , 
        \reg_out<72> , \reg_out<71> , \reg_out<70> , \reg_out<69> , 
        \reg_out<68> , \reg_out<67> , \reg_out<66> , \reg_out<65> , 
        \reg_out<64> , \reg_out<63> , \reg_out<62> , \reg_out<61> , 
        \reg_out<60> , \reg_out<59> , \reg_out<58> , \reg_out<57> , 
        \reg_out<56> , \reg_out<55> , \reg_out<54> , \reg_out<53> , 
        \reg_out<52> , \reg_out<51> , \reg_out<50> , \reg_out<49> , 
        \reg_out<48> , \reg_out<47> , \reg_out<46> , \reg_out<45> , 
        \reg_out<44> , \reg_out<43> , \reg_out<42> , \reg_out<41> , 
        \reg_out<40> , \reg_out<39> , \reg_out<38> , \reg_out<37> , 
        \reg_out<36> , \reg_out<35> , \reg_out<34> , \reg_out<33> , 
        \reg_out<32> , \reg_out<31> , \reg_out<30> , \reg_out<29> , 
        \reg_out<28> , \reg_out<27> , \reg_out<26> , \reg_out<25> , 
        \reg_out<24> , \reg_out<23> , \reg_out<22> , \reg_out<21> , 
        \reg_out<20> , \reg_out<19> , \reg_out<18> , \reg_out<17> , 
        \reg_out<16> , \reg_out<15> , \reg_out<14> , \reg_out<13> , 
        \reg_out<12> , \reg_out<11> , \reg_out<10> , \reg_out<9> , 
        \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , 
        \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> }), .Sel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .Out({
        \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> , 
        \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> , 
        \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> , 
        \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> }) );
  demux1to8_16 wr_demux ( .In({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .S({\writeregsel<2> , 
        \writeregsel<1> , n1}), .Out0({\reg_in<15> , \reg_in<14> , 
        \reg_in<13> , \reg_in<12> , \reg_in<11> , \reg_in<10> , \reg_in<9> , 
        \reg_in<8> , \reg_in<7> , \reg_in<6> , \reg_in<5> , \reg_in<4> , 
        \reg_in<3> , \reg_in<2> , \reg_in<1> , \reg_in<0> }), .Out1({
        \reg_in<31> , \reg_in<30> , \reg_in<29> , \reg_in<28> , \reg_in<27> , 
        \reg_in<26> , \reg_in<25> , \reg_in<24> , \reg_in<23> , \reg_in<22> , 
        \reg_in<21> , \reg_in<20> , \reg_in<19> , \reg_in<18> , \reg_in<17> , 
        \reg_in<16> }), .Out2({\reg_in<47> , \reg_in<46> , \reg_in<45> , 
        \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> , 
        \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> , 
        \reg_in<34> , \reg_in<33> , \reg_in<32> }), .Out3({\reg_in<63> , 
        \reg_in<62> , \reg_in<61> , \reg_in<60> , \reg_in<59> , \reg_in<58> , 
        \reg_in<57> , \reg_in<56> , \reg_in<55> , \reg_in<54> , \reg_in<53> , 
        \reg_in<52> , \reg_in<51> , \reg_in<50> , \reg_in<49> , \reg_in<48> }), 
        .Out4({\reg_in<79> , \reg_in<78> , \reg_in<77> , \reg_in<76> , 
        \reg_in<75> , \reg_in<74> , \reg_in<73> , \reg_in<72> , \reg_in<71> , 
        \reg_in<70> , \reg_in<69> , \reg_in<68> , \reg_in<67> , \reg_in<66> , 
        \reg_in<65> , \reg_in<64> }), .Out5({\reg_in<95> , \reg_in<94> , 
        \reg_in<93> , \reg_in<92> , \reg_in<91> , \reg_in<90> , \reg_in<89> , 
        \reg_in<88> , \reg_in<87> , \reg_in<86> , \reg_in<85> , \reg_in<84> , 
        \reg_in<83> , \reg_in<82> , \reg_in<81> , \reg_in<80> }), .Out6({
        \reg_in<111> , \reg_in<110> , \reg_in<109> , \reg_in<108> , 
        \reg_in<107> , \reg_in<106> , \reg_in<105> , \reg_in<104> , 
        \reg_in<103> , \reg_in<102> , \reg_in<101> , \reg_in<100> , 
        \reg_in<99> , \reg_in<98> , \reg_in<97> , \reg_in<96> }), .Out7({
        \reg_in<127> , \reg_in<126> , \reg_in<125> , \reg_in<124> , 
        \reg_in<123> , \reg_in<122> , \reg_in<121> , \reg_in<120> , 
        \reg_in<119> , \reg_in<118> , \reg_in<117> , \reg_in<116> , 
        \reg_in<115> , \reg_in<114> , \reg_in<113> , \reg_in<112> }) );
  BUFX2 U10 ( .A(rst), .Y(n3) );
  BUFX2 U11 ( .A(rst), .Y(n4) );
  INVX1 U12 ( .A(n2), .Y(n1) );
  INVX1 U13 ( .A(\writeregsel<0> ), .Y(n2) );
endmodule


module control_unit ( .opcode({\opcode<4> , \opcode<3> , \opcode<2> , 
        \opcode<1> , \opcode<0> }), .func({\func<1> , \func<0> }), .aluop({
        \aluop<2> , \aluop<1> , \aluop<0> }), alusrc, branch, jump, i1, i2, r, 
        jumpreg, set, btr, regwrite, memwrite, memread, memtoreg, invA, invB, 
        cin, excp, zeroext, halt, slbi, link, lbi, stu, rti );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ,
         \func<1> , \func<0> ;
  output \aluop<2> , \aluop<1> , \aluop<0> , alusrc, branch, jump, i1, i2, r,
         jumpreg, set, btr, regwrite, memwrite, memread, memtoreg, invA, invB,
         cin, excp, zeroext, halt, slbi, link, lbi, stu, rti;
  wire   n162, N20, N55, n1, n2, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18,
         n19, n21, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50,
         n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n88, n89, n90, n92, n93, n94, n95, n97, n98,
         n100, n101, n103, n104, n105, n106, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160;
  assign \aluop<2>  = N20;
  assign \aluop<0>  = N55;

  INVX2 U1 ( .A(\func<1> ), .Y(n153) );
  INVX4 U2 ( .A(n10), .Y(invB) );
  INVX1 U3 ( .A(n2), .Y(n141) );
  AND2X1 U4 ( .A(n53), .B(n151), .Y(n41) );
  INVX1 U5 ( .A(n125), .Y(memread) );
  OR2X2 U6 ( .A(n38), .B(n105), .Y(n1) );
  MUX2X1 U7 ( .B(n114), .A(n3), .S(n106), .Y(n2) );
  INVX1 U8 ( .A(n140), .Y(n3) );
  INVX1 U9 ( .A(\func<0> ), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(n5) );
  OR2X2 U11 ( .A(n74), .B(n138), .Y(n6) );
  INVX1 U12 ( .A(n6), .Y(halt) );
  AND2X2 U13 ( .A(n52), .B(n37), .Y(n8) );
  INVX1 U14 ( .A(n8), .Y(cin) );
  AND2X2 U15 ( .A(n53), .B(n51), .Y(n10) );
  OR2X2 U16 ( .A(n40), .B(n154), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(btr) );
  OR2X2 U18 ( .A(n58), .B(n129), .Y(n14) );
  INVX1 U19 ( .A(n14), .Y(jumpreg) );
  AND2X2 U20 ( .A(n83), .B(n35), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(\aluop<1> ) );
  OR2X2 U22 ( .A(n111), .B(n109), .Y(n18) );
  INVX1 U23 ( .A(n18), .Y(n19) );
  AND2X2 U24 ( .A(n55), .B(n121), .Y(lbi) );
  OR2X2 U25 ( .A(n58), .B(n139), .Y(n21) );
  INVX1 U26 ( .A(n21), .Y(link) );
  AND2X2 U27 ( .A(\opcode<1> ), .B(n144), .Y(n23) );
  AND2X2 U28 ( .A(n148), .B(n23), .Y(n24) );
  OR2X2 U29 ( .A(n60), .B(n65), .Y(n25) );
  INVX1 U30 ( .A(n25), .Y(memwrite) );
  AND2X2 U31 ( .A(n146), .B(n119), .Y(n27) );
  INVX1 U32 ( .A(n27), .Y(n28) );
  AND2X2 U33 ( .A(n123), .B(n71), .Y(n29) );
  INVX1 U34 ( .A(n29), .Y(n30) );
  AND2X2 U35 ( .A(n131), .B(n123), .Y(n31) );
  INVX1 U36 ( .A(n31), .Y(n32) );
  AND2X2 U37 ( .A(n131), .B(n158), .Y(n33) );
  INVX1 U38 ( .A(n33), .Y(n34) );
  BUFX2 U39 ( .A(n156), .Y(n35) );
  AND2X2 U40 ( .A(n66), .B(n104), .Y(n36) );
  INVX1 U41 ( .A(n36), .Y(n37) );
  AND2X2 U42 ( .A(\func<1> ), .B(\func<0> ), .Y(n38) );
  AND2X2 U43 ( .A(\opcode<4> ), .B(n127), .Y(n39) );
  INVX1 U44 ( .A(n39), .Y(n40) );
  INVX1 U45 ( .A(n41), .Y(n42) );
  AND2X2 U46 ( .A(n28), .B(n158), .Y(n43) );
  INVX1 U47 ( .A(n43), .Y(n44) );
  AND2X2 U48 ( .A(n64), .B(n108), .Y(n45) );
  INVX1 U49 ( .A(n45), .Y(n46) );
  INVX1 U50 ( .A(n59), .Y(n47) );
  OR2X2 U51 ( .A(n73), .B(n136), .Y(n48) );
  INVX1 U52 ( .A(n48), .Y(slbi) );
  AND2X2 U53 ( .A(n61), .B(set), .Y(n50) );
  INVX1 U54 ( .A(n50), .Y(n51) );
  INVX1 U55 ( .A(n50), .Y(n52) );
  BUFX2 U56 ( .A(n150), .Y(n53) );
  OR2X2 U57 ( .A(n134), .B(n113), .Y(n54) );
  INVX1 U58 ( .A(n54), .Y(n55) );
  INVX1 U59 ( .A(n54), .Y(n56) );
  AND2X2 U60 ( .A(n131), .B(n137), .Y(jump) );
  INVX1 U61 ( .A(jump), .Y(n58) );
  AND2X2 U62 ( .A(n118), .B(n82), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(n60) );
  INVX1 U64 ( .A(n59), .Y(n61) );
  AND2X2 U65 ( .A(n131), .B(n121), .Y(set) );
  AND2X2 U66 ( .A(n148), .B(n132), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(n64) );
  INVX1 U68 ( .A(n63), .Y(n65) );
  AND2X2 U69 ( .A(n135), .B(n111), .Y(n66) );
  AND2X2 U70 ( .A(n63), .B(n127), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(n68) );
  AND2X2 U72 ( .A(n124), .B(n115), .Y(n69) );
  INVX1 U73 ( .A(n69), .Y(n70) );
  AND2X2 U74 ( .A(n131), .B(n111), .Y(n71) );
  BUFX2 U75 ( .A(n143), .Y(n72) );
  INVX1 U76 ( .A(n24), .Y(n73) );
  BUFX2 U77 ( .A(n120), .Y(n74) );
  INVX4 U78 ( .A(n159), .Y(n119) );
  INVX1 U79 ( .A(n123), .Y(n158) );
  AND2X2 U80 ( .A(n146), .B(n119), .Y(n75) );
  OR2X1 U81 ( .A(n94), .B(n77), .Y(i2) );
  OR2X1 U82 ( .A(n92), .B(n93), .Y(n77) );
  AND2X2 U83 ( .A(n123), .B(n112), .Y(n78) );
  INVX1 U84 ( .A(n78), .Y(n79) );
  INVX1 U85 ( .A(memtoreg), .Y(n125) );
  INVX1 U86 ( .A(n68), .Y(memtoreg) );
  AND2X2 U87 ( .A(n5), .B(\opcode<4> ), .Y(n80) );
  INVX1 U88 ( .A(n80), .Y(n81) );
  INVX1 U89 ( .A(n23), .Y(n82) );
  BUFX2 U90 ( .A(n157), .Y(n83) );
  AND2X2 U91 ( .A(n111), .B(n117), .Y(n84) );
  INVX1 U92 ( .A(n84), .Y(n85) );
  INVX1 U93 ( .A(n84), .Y(n86) );
  INVX1 U94 ( .A(n85), .Y(n142) );
  AND2X2 U95 ( .A(n131), .B(n75), .Y(branch) );
  INVX1 U96 ( .A(branch), .Y(n88) );
  INVX1 U97 ( .A(set), .Y(n89) );
  OR2X1 U98 ( .A(n97), .B(n100), .Y(n90) );
  INVX1 U99 ( .A(n90), .Y(stu) );
  INVX1 U100 ( .A(n147), .Y(n92) );
  INVX1 U101 ( .A(n88), .Y(n93) );
  INVX1 U102 ( .A(n133), .Y(n94) );
  AND2X2 U103 ( .A(n133), .B(n83), .Y(n95) );
  INVX1 U104 ( .A(n95), .Y(zeroext) );
  INVX1 U105 ( .A(n138), .Y(n137) );
  BUFX2 U106 ( .A(n86), .Y(n97) );
  OR2X2 U107 ( .A(n112), .B(n138), .Y(n98) );
  INVX1 U108 ( .A(n98), .Y(excp) );
  INVX1 U109 ( .A(n63), .Y(n100) );
  INVX1 U110 ( .A(n162), .Y(n101) );
  INVX1 U111 ( .A(n101), .Y(regwrite) );
  INVX2 U112 ( .A(n135), .Y(n154) );
  INVX1 U113 ( .A(n141), .Y(n103) );
  INVX1 U114 ( .A(n103), .Y(n104) );
  INVX1 U115 ( .A(\opcode<4> ), .Y(n105) );
  INVX1 U116 ( .A(n105), .Y(n106) );
  AND2X2 U117 ( .A(n141), .B(n66), .Y(invA) );
  INVX1 U118 ( .A(n75), .Y(n108) );
  INVX1 U119 ( .A(n114), .Y(n109) );
  BUFX2 U120 ( .A(n19), .Y(n110) );
  INVX1 U121 ( .A(n128), .Y(n111) );
  INVX4 U122 ( .A(n130), .Y(n131) );
  BUFX2 U123 ( .A(n73), .Y(n112) );
  INVX1 U124 ( .A(n116), .Y(n113) );
  INVX1 U125 ( .A(\opcode<1> ), .Y(n114) );
  INVX1 U126 ( .A(n56), .Y(n115) );
  INVX1 U127 ( .A(\opcode<1> ), .Y(n116) );
  INVX1 U128 ( .A(n116), .Y(n117) );
  INVX4 U129 ( .A(\opcode<3> ), .Y(n159) );
  INVX1 U130 ( .A(\opcode<2> ), .Y(n148) );
  OR2X2 U131 ( .A(\opcode<1> ), .B(n128), .Y(n118) );
  INVX1 U132 ( .A(n118), .Y(n127) );
  INVX2 U133 ( .A(\opcode<4> ), .Y(n146) );
  OR2X2 U134 ( .A(n134), .B(n109), .Y(n120) );
  AND2X2 U135 ( .A(\opcode<4> ), .B(\opcode<3> ), .Y(n121) );
  INVX1 U136 ( .A(n121), .Y(n145) );
  INVX1 U137 ( .A(n139), .Y(n122) );
  AND2X2 U138 ( .A(\opcode<4> ), .B(n159), .Y(n123) );
  INVX1 U139 ( .A(n146), .Y(n124) );
  INVX1 U140 ( .A(\opcode<0> ), .Y(n144) );
  INVX1 U141 ( .A(\opcode<0> ), .Y(n128) );
  INVX1 U142 ( .A(\opcode<1> ), .Y(n139) );
  BUFX2 U143 ( .A(n144), .Y(n129) );
  INVX1 U144 ( .A(\opcode<2> ), .Y(n130) );
  AND2X2 U145 ( .A(\opcode<4> ), .B(n159), .Y(n132) );
  BUFX2 U146 ( .A(n151), .Y(n133) );
  INVX1 U147 ( .A(n132), .Y(n136) );
  OR2X2 U148 ( .A(\opcode<0> ), .B(\opcode<2> ), .Y(n134) );
  INVX1 U149 ( .A(slbi), .Y(n151) );
  AND2X2 U150 ( .A(n148), .B(\opcode<3> ), .Y(n135) );
  OR2X2 U151 ( .A(n119), .B(n106), .Y(n138) );
  NOR3X1 U152 ( .A(n97), .B(n138), .C(n131), .Y(rti) );
  NAND3X1 U153 ( .A(n122), .B(n135), .C(n146), .Y(n157) );
  NAND3X1 U154 ( .A(n5), .B(n117), .C(n153), .Y(n140) );
  NAND3X1 U155 ( .A(n135), .B(n142), .C(n1), .Y(n150) );
  NAND3X1 U156 ( .A(n131), .B(n122), .C(n159), .Y(n143) );
  NAND3X1 U157 ( .A(n72), .B(n154), .C(n70), .Y(n162) );
  OAI21X1 U158 ( .A(n110), .B(n145), .C(n89), .Y(r) );
  AOI21X1 U159 ( .A(n146), .B(n71), .C(lbi), .Y(n147) );
  OAI21X1 U160 ( .A(n154), .B(n124), .C(n79), .Y(i1) );
  MUX2X1 U161 ( .B(n130), .A(n120), .S(n119), .Y(n149) );
  OR2X2 U162 ( .A(n149), .B(n44), .Y(alusrc) );
  OAI21X1 U163 ( .A(n81), .B(n112), .C(n30), .Y(n152) );
  OR2X2 U164 ( .A(n42), .B(n152), .Y(N55) );
  OAI21X1 U165 ( .A(n154), .B(n153), .C(n32), .Y(n155) );
  AOI22X1 U166 ( .A(n19), .B(set), .C(n122), .D(n155), .Y(n156) );
  OAI21X1 U167 ( .A(n159), .B(n47), .C(n34), .Y(n160) );
  OR2X2 U168 ( .A(n160), .B(n46), .Y(N20) );
endmodule


module alu ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , 
        \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> 
        }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , 
        \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> 
        }), Cin, .Op({\Op<2> , \Op<1> , \Op<0> }), invA, invB, sign, .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Ofl, Z, Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<2> , \Op<1> , \Op<0> , invA, invB, sign;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Ofl, Z, Cout;
  wire   \A_real<15> , \A_real<14> , \A_real<13> , \A_real<12> , \A_real<11> ,
         \A_real<10> , \A_real<9> , \A_real<8> , \A_real<7> , \A_real<6> ,
         \A_real<5> , \A_real<4> , \A_real<3> , \A_real<2> , \A_real<1> ,
         \A_real<0> , \B_real<15> , \B_real<14> , \B_real<13> , \B_real<12> ,
         \B_real<11> , \B_real<10> , \B_real<9> , \B_real<8> , \B_real<7> ,
         \B_real<6> , \B_real<5> , \B_real<4> , \B_real<3> , \B_real<2> ,
         \B_real<1> , \B_real<0> , \op0_out<15> , \op0_out<14> , \op0_out<13> ,
         \op0_out<12> , \op0_out<11> , \op0_out<10> , \op0_out<9> ,
         \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , \op0_out<4> ,
         \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> , \op1_out<15> ,
         \op1_out<14> , \op1_out<13> , \op1_out<12> , \op1_out<11> ,
         \op1_out<10> , \op1_out<9> , \op1_out<8> , \op1_out<7> , \op1_out<6> ,
         \op1_out<5> , \op1_out<4> , \op1_out<3> , \op1_out<2> , \op1_out<1> ,
         \op1_out<0> , \op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> ,
         \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> ,
         \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> ,
         \op0_A<1> , \op0_A<0> , \op0_B<15> , \op0_B<14> , \op0_B<13> ,
         \op0_B<12> , \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> ,
         \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> ,
         \op0_B<2> , \op0_B<1> , \op0_B<0> , \op1_A<3> , \op1_A<2> ,
         \op1_A<1> , \op1_A<0> , \op1_B<15> , \op1_B<14> , \op1_B<13> ,
         \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> ,
         \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> ,
         \op1_B<2> , \op1_B<1> , \op1_B<0> , n59, n60, n62, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n61, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  OR2X2 U4 ( .A(n72), .B(n74), .Y(n62) );
  NAND3X1 U76 ( .A(Cout), .B(n85), .C(n84), .Y(n59) );
  demux1to2_16_1 demux0 ( .In({\A_real<15> , \A_real<14> , \A_real<13> , 
        \A_real<12> , \A_real<11> , \A_real<10> , \A_real<9> , \A_real<8> , 
        \A_real<7> , \A_real<6> , \A_real<5> , \A_real<4> , \A_real<3> , 
        \A_real<2> , \A_real<1> , \A_real<0> }), .S(n101), .Out0({\op0_A<15> , 
        \op0_A<14> , \op0_A<13> , \op0_A<12> , \op0_A<11> , \op0_A<10> , 
        \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , \op0_A<5> , \op0_A<4> , 
        \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .Out1({\op0_B<15> , 
        \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , \op0_B<10> , 
        \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , 
        \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }) );
  demux1to2_16_0 demux1 ( .In({\B_real<15> , \B_real<14> , \B_real<13> , 
        \B_real<12> , \B_real<11> , \B_real<10> , \B_real<9> , \B_real<8> , 
        \B_real<7> , \B_real<6> , \B_real<5> , \B_real<4> , \B_real<3> , 
        \B_real<2> , \B_real<1> , \B_real<0> }), .S(n99), .Out0({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, \op1_A<3> , 
        \op1_A<2> , \op1_A<1> , \op1_A<0> }), .Out1({\op1_B<15> , \op1_B<14> , 
        \op1_B<13> , \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , 
        \op1_B<8> , \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , 
        \op1_B<2> , \op1_B<1> , \op1_B<0> }) );
  cla_or_xor_and coxa0 ( .A({\op0_B<15> , \op0_B<14> , \op0_B<13> , 
        \op0_B<12> , \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> , 
        \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , 
        \op0_B<1> , \op0_B<0> }), .B({\op1_B<15> , \op1_B<14> , \op1_B<13> , 
        \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , 
        \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> , 
        \op1_B<1> , \op1_B<0> }), .Cin(Cin), .Op({n58, \Op<0> }), .Out({
        \op0_out<15> , \op0_out<14> , \op0_out<13> , \op0_out<12> , 
        \op0_out<11> , \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , 
        \op0_out<6> , \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , 
        \op0_out<1> , \op0_out<0> }), .Cout(Cout) );
  shifter shift ( .In({\op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> , 
        \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> , 
        \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> , \op0_A<1> , 
        \op0_A<0> }), .Cnt({\op1_A<3> , \op1_A<2> , \op1_A<1> , \op1_A<0> }), 
        .Op({n72, n74}), .Out({\op1_out<15> , \op1_out<14> , \op1_out<13> , 
        \op1_out<12> , \op1_out<11> , \op1_out<10> , \op1_out<9> , 
        \op1_out<8> , \op1_out<7> , \op1_out<6> , \op1_out<5> , \op1_out<4> , 
        \op1_out<3> , \op1_out<2> , \op1_out<1> , \op1_out<0> }) );
  XNOR2X1 U1 ( .A(\B<3> ), .B(n86), .Y(\B_real<3> ) );
  INVX1 U2 ( .A(\A<7> ), .Y(n5) );
  INVX1 U3 ( .A(\A<5> ), .Y(n1) );
  INVX1 U5 ( .A(\A<2> ), .Y(n4) );
  AND2X1 U6 ( .A(n112), .B(n98), .Y(n55) );
  INVX1 U7 ( .A(\A<3> ), .Y(n10) );
  INVX1 U8 ( .A(n11), .Y(\Out<6> ) );
  INVX1 U9 ( .A(n85), .Y(n12) );
  INVX1 U10 ( .A(n130), .Y(n18) );
  INVX1 U11 ( .A(\op1_out<12> ), .Y(n130) );
  INVX1 U12 ( .A(n97), .Y(n15) );
  INVX8 U13 ( .A(\Op<2> ), .Y(n107) );
  INVX1 U14 ( .A(n85), .Y(n16) );
  INVX1 U15 ( .A(n85), .Y(n13) );
  INVX1 U16 ( .A(n85), .Y(n14) );
  XNOR2X1 U17 ( .A(\B<0> ), .B(n86), .Y(\B_real<0> ) );
  INVX4 U18 ( .A(invB), .Y(n86) );
  XNOR2X1 U19 ( .A(n1), .B(n106), .Y(\A_real<5> ) );
  INVX2 U20 ( .A(n105), .Y(n2) );
  BUFX2 U21 ( .A(n65), .Y(n3) );
  XNOR2X1 U22 ( .A(\B<5> ), .B(n71), .Y(\B_real<5> ) );
  INVX4 U23 ( .A(n86), .Y(n87) );
  INVX2 U24 ( .A(invB), .Y(n71) );
  XNOR2X1 U25 ( .A(\B<8> ), .B(n71), .Y(\B_real<8> ) );
  XOR2X1 U26 ( .A(\B<7> ), .B(n87), .Y(\B_real<7> ) );
  XNOR2X1 U27 ( .A(\B<10> ), .B(n86), .Y(\B_real<10> ) );
  INVX8 U28 ( .A(n105), .Y(n106) );
  XNOR2X1 U29 ( .A(n4), .B(n106), .Y(\A_real<2> ) );
  XNOR2X1 U30 ( .A(invA), .B(n5), .Y(\A_real<7> ) );
  XNOR2X1 U31 ( .A(\B<12> ), .B(n71), .Y(\B_real<12> ) );
  XOR2X1 U32 ( .A(\B<1> ), .B(invB), .Y(\B_real<1> ) );
  XOR2X1 U33 ( .A(\B<6> ), .B(n87), .Y(\B_real<6> ) );
  MUX2X1 U34 ( .B(n67), .A(\op1_out<9> ), .S(n13), .Y(n102) );
  INVX1 U35 ( .A(n57), .Y(n6) );
  INVX1 U36 ( .A(n2), .Y(n93) );
  INVX1 U37 ( .A(n128), .Y(n7) );
  INVX1 U38 ( .A(n69), .Y(n8) );
  INVX1 U39 ( .A(n8), .Y(n9) );
  XNOR2X1 U40 ( .A(n10), .B(n106), .Y(\A_real<3> ) );
  MUX2X1 U41 ( .B(\op0_out<6> ), .A(\op1_out<6> ), .S(n12), .Y(n11) );
  INVX4 U42 ( .A(invA), .Y(n105) );
  XNOR2X1 U43 ( .A(\B<2> ), .B(n86), .Y(\B_real<2> ) );
  MUX2X1 U44 ( .B(n124), .A(n125), .S(n107), .Y(\Out<5> ) );
  MUX2X1 U45 ( .B(n61), .A(n18), .S(n13), .Y(n17) );
  BUFX2 U46 ( .A(\op0_out<8> ), .Y(n88) );
  XNOR2X1 U47 ( .A(\B<9> ), .B(n86), .Y(\B_real<9> ) );
  MUX2X1 U48 ( .B(n7), .A(\op1_out<10> ), .S(n14), .Y(n95) );
  INVX1 U49 ( .A(n57), .Y(n128) );
  XOR2X1 U50 ( .A(\B<11> ), .B(n15), .Y(\B_real<11> ) );
  MUX2X1 U51 ( .B(\op0_out<7> ), .A(\op1_out<7> ), .S(n16), .Y(n91) );
  AND2X2 U52 ( .A(n45), .B(n35), .Y(n52) );
  INVX1 U53 ( .A(n17), .Y(\Out<12> ) );
  AND2X2 U54 ( .A(n52), .B(n56), .Y(n19) );
  AND2X2 U55 ( .A(n90), .B(n55), .Y(n20) );
  BUFX4 U56 ( .A(\Op<1> ), .Y(n58) );
  OR2X2 U57 ( .A(\op1_out<2> ), .B(n73), .Y(n21) );
  INVX1 U58 ( .A(n21), .Y(n22) );
  AND2X2 U59 ( .A(n79), .B(n49), .Y(\Out<8> ) );
  OR2X2 U60 ( .A(\op1_out<8> ), .B(\op1_out<9> ), .Y(n24) );
  INVX1 U61 ( .A(n24), .Y(n25) );
  OR2X2 U62 ( .A(\op1_out<12> ), .B(\op1_out<13> ), .Y(n26) );
  INVX1 U63 ( .A(n26), .Y(n27) );
  AND2X2 U64 ( .A(n51), .B(n118), .Y(n28) );
  INVX1 U65 ( .A(n28), .Y(n29) );
  OR2X2 U66 ( .A(\op1_out<4> ), .B(\op1_out<5> ), .Y(n30) );
  INVX1 U67 ( .A(n30), .Y(n31) );
  OR2X2 U68 ( .A(n64), .B(n29), .Y(n32) );
  INVX1 U69 ( .A(n32), .Y(n33) );
  OR2X2 U70 ( .A(n65), .B(\op0_out<11> ), .Y(n34) );
  INVX1 U71 ( .A(n34), .Y(n35) );
  OR2X2 U72 ( .A(n54), .B(n67), .Y(n36) );
  INVX1 U73 ( .A(n36), .Y(n37) );
  OR2X1 U74 ( .A(\op1_out<10> ), .B(\op1_out<11> ), .Y(n38) );
  INVX1 U75 ( .A(n38), .Y(n39) );
  OR2X1 U77 ( .A(\op1_out<14> ), .B(\op1_out<15> ), .Y(n40) );
  INVX1 U78 ( .A(n40), .Y(n41) );
  OR2X2 U79 ( .A(\op1_out<6> ), .B(\op1_out<7> ), .Y(n42) );
  INVX1 U80 ( .A(n42), .Y(n43) );
  OR2X2 U81 ( .A(n69), .B(n68), .Y(n44) );
  INVX1 U82 ( .A(n44), .Y(n45) );
  AND2X2 U83 ( .A(n85), .B(n19), .Y(n46) );
  INVX1 U84 ( .A(n46), .Y(n47) );
  AND2X2 U85 ( .A(n100), .B(n126), .Y(n48) );
  INVX1 U86 ( .A(n48), .Y(n49) );
  OR2X2 U87 ( .A(\op0_out<1> ), .B(n70), .Y(n50) );
  INVX1 U88 ( .A(n50), .Y(n51) );
  AND2X2 U89 ( .A(n6), .B(n96), .Y(n53) );
  INVX1 U90 ( .A(n53), .Y(n54) );
  AND2X2 U91 ( .A(n37), .B(n20), .Y(n56) );
  BUFX2 U92 ( .A(\op0_out<10> ), .Y(n57) );
  BUFX2 U93 ( .A(\op0_out<12> ), .Y(n61) );
  BUFX2 U94 ( .A(\op0_out<1> ), .Y(n63) );
  BUFX2 U95 ( .A(\op0_out<4> ), .Y(n64) );
  BUFX2 U96 ( .A(\op0_out<14> ), .Y(n65) );
  BUFX2 U97 ( .A(\op0_out<3> ), .Y(n66) );
  BUFX2 U98 ( .A(\op0_out<9> ), .Y(n67) );
  BUFX2 U99 ( .A(\op0_out<13> ), .Y(n68) );
  BUFX2 U100 ( .A(\op0_out<15> ), .Y(n69) );
  INVX1 U101 ( .A(n114), .Y(n70) );
  XNOR2X1 U102 ( .A(\B<4> ), .B(n71), .Y(\B_real<4> ) );
  BUFX2 U103 ( .A(n58), .Y(n72) );
  INVX1 U104 ( .A(n121), .Y(n73) );
  BUFX2 U105 ( .A(\Op<0> ), .Y(n74) );
  INVX1 U106 ( .A(n106), .Y(n75) );
  XNOR2X1 U107 ( .A(\A<11> ), .B(n75), .Y(\A_real<11> ) );
  AND2X2 U108 ( .A(n129), .B(n107), .Y(n76) );
  INVX1 U109 ( .A(n76), .Y(n77) );
  AND2X2 U110 ( .A(n127), .B(n16), .Y(n78) );
  INVX1 U111 ( .A(n78), .Y(n79) );
  INVX1 U112 ( .A(n91), .Y(\Out<7> ) );
  INVX1 U113 ( .A(\op0_out<2> ), .Y(n118) );
  BUFX2 U114 ( .A(n59), .Y(n80) );
  INVX1 U115 ( .A(n80), .Y(Ofl) );
  AND2X2 U116 ( .A(n109), .B(n108), .Y(n81) );
  INVX1 U117 ( .A(n81), .Y(n82) );
  BUFX2 U118 ( .A(n113), .Y(n83) );
  BUFX2 U119 ( .A(n60), .Y(n84) );
  INVX1 U120 ( .A(\op0_out<0> ), .Y(n114) );
  INVX1 U121 ( .A(n63), .Y(n116) );
  OAI21X1 U122 ( .A(\op0_out<11> ), .B(n107), .C(n77), .Y(n94) );
  MUX2X1 U123 ( .B(\op1_out<13> ), .A(n68), .S(\Op<2> ), .Y(n103) );
  INVX8 U124 ( .A(n107), .Y(n85) );
  XNOR2X1 U125 ( .A(\A<8> ), .B(n93), .Y(\A_real<8> ) );
  INVX1 U126 ( .A(n92), .Y(\Out<15> ) );
  INVX1 U127 ( .A(\op0_out<8> ), .Y(n89) );
  INVX1 U128 ( .A(n64), .Y(n122) );
  INVX1 U129 ( .A(\op1_out<8> ), .Y(n127) );
  INVX1 U130 ( .A(n107), .Y(n100) );
  INVX1 U131 ( .A(n131), .Y(\A_real<15> ) );
  INVX1 U132 ( .A(\op1_out<1> ), .Y(n117) );
  INVX1 U133 ( .A(n61), .Y(n90) );
  MUX2X1 U134 ( .B(\op1_out<15> ), .A(n9), .S(n100), .Y(n92) );
  XOR2X1 U135 ( .A(n2), .B(\A<9> ), .Y(\A_real<9> ) );
  INVX1 U136 ( .A(n95), .Y(\Out<10> ) );
  INVX1 U137 ( .A(invB), .Y(n97) );
  INVX1 U138 ( .A(n94), .Y(\Out<11> ) );
  INVX1 U139 ( .A(\op1_out<11> ), .Y(n129) );
  INVX1 U140 ( .A(n88), .Y(n126) );
  AND2X2 U141 ( .A(n33), .B(n89), .Y(n96) );
  INVX1 U142 ( .A(\op0_out<7> ), .Y(n98) );
  INVX1 U143 ( .A(\op0_out<5> ), .Y(n124) );
  INVX8 U144 ( .A(n107), .Y(n99) );
  INVX8 U145 ( .A(n107), .Y(n101) );
  INVX1 U146 ( .A(n102), .Y(\Out<9> ) );
  INVX1 U147 ( .A(n103), .Y(\Out<13> ) );
  MUX2X1 U148 ( .B(n3), .A(\op1_out<14> ), .S(n14), .Y(n104) );
  INVX1 U149 ( .A(n66), .Y(n120) );
  INVX1 U150 ( .A(n104), .Y(\Out<14> ) );
  XNOR2X1 U151 ( .A(\B<15> ), .B(n87), .Y(n132) );
  INVX2 U152 ( .A(n132), .Y(\B_real<15> ) );
  XOR2X1 U153 ( .A(\B<14> ), .B(n87), .Y(\B_real<14> ) );
  XOR2X1 U154 ( .A(\B<13> ), .B(n87), .Y(\B_real<13> ) );
  XNOR2X1 U155 ( .A(\A<15> ), .B(n106), .Y(n131) );
  XOR2X1 U156 ( .A(\A<14> ), .B(n2), .Y(\A_real<14> ) );
  XOR2X1 U157 ( .A(\A<13> ), .B(n2), .Y(\A_real<13> ) );
  XOR2X1 U158 ( .A(\A<12> ), .B(n106), .Y(\A_real<12> ) );
  XOR2X1 U159 ( .A(\A<10> ), .B(n2), .Y(\A_real<10> ) );
  XOR2X1 U160 ( .A(\A<6> ), .B(n106), .Y(\A_real<6> ) );
  XOR2X1 U161 ( .A(\A<4> ), .B(n106), .Y(\A_real<4> ) );
  XOR2X1 U162 ( .A(\A<1> ), .B(n106), .Y(\A_real<1> ) );
  XOR2X1 U163 ( .A(\A<0> ), .B(n2), .Y(\A_real<0> ) );
  AND2X2 U164 ( .A(n25), .B(n39), .Y(n109) );
  AND2X2 U165 ( .A(n27), .B(n41), .Y(n108) );
  NOR3X1 U166 ( .A(\op1_out<1> ), .B(n85), .C(\op1_out<0> ), .Y(n111) );
  AND2X2 U167 ( .A(n31), .B(n43), .Y(n110) );
  NAND3X1 U168 ( .A(n111), .B(n22), .C(n110), .Y(n113) );
  NOR3X1 U169 ( .A(n66), .B(\op0_out<6> ), .C(\op0_out<5> ), .Y(n112) );
  OAI21X1 U170 ( .A(n82), .B(n83), .C(n47), .Y(Z) );
  INVX2 U171 ( .A(\op1_out<0> ), .Y(n115) );
  MUX2X1 U172 ( .B(n115), .A(n114), .S(n100), .Y(\Out<0> ) );
  MUX2X1 U173 ( .B(n117), .A(n116), .S(n85), .Y(\Out<1> ) );
  INVX2 U174 ( .A(\op1_out<2> ), .Y(n119) );
  MUX2X1 U175 ( .B(n119), .A(n118), .S(n100), .Y(\Out<2> ) );
  INVX2 U176 ( .A(\op1_out<3> ), .Y(n121) );
  MUX2X1 U177 ( .B(n121), .A(n120), .S(n85), .Y(\Out<3> ) );
  INVX2 U178 ( .A(\op1_out<4> ), .Y(n123) );
  MUX2X1 U179 ( .B(n123), .A(n122), .S(n100), .Y(\Out<4> ) );
  INVX2 U180 ( .A(\op1_out<5> ), .Y(n125) );
  XNOR2X1 U181 ( .A(n132), .B(n131), .Y(n133) );
  AOI21X1 U182 ( .A(sign), .B(n133), .C(n62), .Y(n60) );
endmodule


module mux4to1_16_5 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n83, n92, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151;

  BUFX2 U1 ( .A(n63), .Y(n119) );
  INVX1 U2 ( .A(n119), .Y(n144) );
  INVX1 U3 ( .A(n119), .Y(n137) );
  INVX1 U4 ( .A(n119), .Y(n139) );
  INVX1 U5 ( .A(n119), .Y(n146) );
  INVX1 U6 ( .A(n119), .Y(n123) );
  INVX1 U7 ( .A(n119), .Y(n142) );
  INVX1 U8 ( .A(n119), .Y(n133) );
  INVX1 U9 ( .A(n119), .Y(n135) );
  INVX1 U10 ( .A(n119), .Y(n129) );
  INVX1 U11 ( .A(n119), .Y(n131) );
  INVX1 U12 ( .A(n119), .Y(n126) );
  AND2X2 U13 ( .A(n68), .B(n3), .Y(n1) );
  INVX1 U14 ( .A(n1), .Y(\Out<13> ) );
  AND2X2 U15 ( .A(n27), .B(n35), .Y(n3) );
  AND2X2 U16 ( .A(\InC<1> ), .B(n66), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n5) );
  AND2X2 U18 ( .A(\InC<2> ), .B(n66), .Y(n6) );
  INVX1 U19 ( .A(n6), .Y(n7) );
  AND2X2 U20 ( .A(\InD<4> ), .B(n129), .Y(n8) );
  INVX1 U21 ( .A(n8), .Y(n9) );
  AND2X2 U22 ( .A(\InD<5> ), .B(n131), .Y(n10) );
  INVX1 U23 ( .A(n10), .Y(n11) );
  AND2X2 U24 ( .A(\InC<6> ), .B(n66), .Y(n12) );
  INVX1 U25 ( .A(n12), .Y(n13) );
  AND2X2 U26 ( .A(\InC<7> ), .B(n66), .Y(n14) );
  INVX1 U27 ( .A(n14), .Y(n15) );
  AND2X2 U28 ( .A(\InC<8> ), .B(n66), .Y(n16) );
  INVX1 U29 ( .A(n16), .Y(n17) );
  AND2X2 U30 ( .A(\InC<9> ), .B(n66), .Y(n18) );
  INVX1 U31 ( .A(n18), .Y(n19) );
  AND2X2 U32 ( .A(\InC<10> ), .B(n66), .Y(n20) );
  INVX1 U33 ( .A(n20), .Y(n21) );
  AND2X2 U34 ( .A(\InC<11> ), .B(n66), .Y(n22) );
  INVX1 U35 ( .A(n22), .Y(n23) );
  AND2X2 U36 ( .A(\InD<12> ), .B(n144), .Y(n24) );
  INVX1 U37 ( .A(n24), .Y(n25) );
  AND2X2 U38 ( .A(\InC<13> ), .B(n66), .Y(n26) );
  INVX1 U39 ( .A(n26), .Y(n27) );
  AND2X2 U40 ( .A(\InC<14> ), .B(n66), .Y(n28) );
  INVX1 U41 ( .A(n28), .Y(n29) );
  AND2X2 U42 ( .A(\InC<15> ), .B(n66), .Y(n30) );
  INVX1 U43 ( .A(n30), .Y(n31) );
  AND2X2 U44 ( .A(\InD<15> ), .B(n131), .Y(n32) );
  INVX1 U45 ( .A(n32), .Y(n33) );
  AND2X2 U46 ( .A(\InD<13> ), .B(n146), .Y(n34) );
  INVX1 U47 ( .A(n34), .Y(n35) );
  BUFX2 U48 ( .A(n122), .Y(n36) );
  AND2X2 U49 ( .A(\InD<1> ), .B(n123), .Y(n37) );
  INVX1 U50 ( .A(n37), .Y(n38) );
  AND2X2 U51 ( .A(\InD<2> ), .B(n126), .Y(n39) );
  INVX1 U52 ( .A(n39), .Y(n40) );
  AND2X2 U53 ( .A(\InC<3> ), .B(n66), .Y(n41) );
  INVX1 U54 ( .A(n41), .Y(n42) );
  AND2X2 U55 ( .A(\InD<6> ), .B(n133), .Y(n43) );
  INVX1 U56 ( .A(n43), .Y(n44) );
  AND2X2 U57 ( .A(\InD<7> ), .B(n135), .Y(n45) );
  INVX1 U58 ( .A(n45), .Y(n46) );
  AND2X2 U59 ( .A(\InD<8> ), .B(n137), .Y(n47) );
  INVX1 U60 ( .A(n47), .Y(n48) );
  AND2X2 U61 ( .A(\InD<9> ), .B(n139), .Y(n49) );
  INVX1 U62 ( .A(n49), .Y(n50) );
  AND2X2 U63 ( .A(\InD<10> ), .B(n131), .Y(n51) );
  INVX1 U64 ( .A(n51), .Y(n52) );
  AND2X2 U65 ( .A(\InD<11> ), .B(n142), .Y(n53) );
  INVX1 U66 ( .A(n53), .Y(n54) );
  AND2X2 U67 ( .A(\InD<14> ), .B(n131), .Y(n55) );
  INVX1 U68 ( .A(n55), .Y(n56) );
  AND2X2 U69 ( .A(n150), .B(\InB<0> ), .Y(n57) );
  INVX1 U70 ( .A(n57), .Y(n58) );
  BUFX2 U71 ( .A(n128), .Y(n59) );
  AND2X2 U72 ( .A(\InC<0> ), .B(n66), .Y(n60) );
  INVX1 U73 ( .A(n60), .Y(n61) );
  AND2X2 U74 ( .A(\S<0> ), .B(\S<1> ), .Y(n62) );
  INVX1 U75 ( .A(n62), .Y(n63) );
  AND2X2 U76 ( .A(\S<0> ), .B(n120), .Y(n64) );
  INVX1 U77 ( .A(n64), .Y(n65) );
  AND2X2 U78 ( .A(n121), .B(\S<1> ), .Y(n66) );
  INVX1 U79 ( .A(n147), .Y(n67) );
  INVX1 U80 ( .A(n67), .Y(n68) );
  INVX1 U81 ( .A(n130), .Y(n69) );
  INVX1 U82 ( .A(n69), .Y(n70) );
  AND2X2 U83 ( .A(\InC<4> ), .B(n66), .Y(n71) );
  INVX1 U84 ( .A(n71), .Y(n72) );
  AND2X2 U85 ( .A(\InC<5> ), .B(n66), .Y(n73) );
  INVX1 U86 ( .A(n73), .Y(n74) );
  INVX1 U87 ( .A(n132), .Y(n75) );
  INVX1 U88 ( .A(n75), .Y(n76) );
  INVX1 U89 ( .A(n145), .Y(n77) );
  INVX1 U90 ( .A(n77), .Y(n78) );
  BUFX2 U91 ( .A(n165), .Y(\Out<1> ) );
  BUFX2 U92 ( .A(n164), .Y(\Out<2> ) );
  BUFX2 U93 ( .A(n163), .Y(\Out<3> ) );
  BUFX2 U94 ( .A(n162), .Y(\Out<4> ) );
  INVX1 U95 ( .A(n161), .Y(n83) );
  INVX1 U96 ( .A(n83), .Y(\Out<5> ) );
  BUFX2 U97 ( .A(n160), .Y(\Out<6> ) );
  BUFX2 U98 ( .A(n159), .Y(\Out<7> ) );
  BUFX2 U99 ( .A(n157), .Y(\Out<9> ) );
  BUFX2 U100 ( .A(n156), .Y(\Out<10> ) );
  BUFX2 U101 ( .A(n152), .Y(\Out<15> ) );
  BUFX2 U102 ( .A(n158), .Y(\Out<8> ) );
  BUFX2 U103 ( .A(n155), .Y(\Out<11> ) );
  INVX1 U104 ( .A(n154), .Y(n92) );
  INVX1 U105 ( .A(n92), .Y(\Out<12> ) );
  BUFX2 U106 ( .A(n153), .Y(\Out<14> ) );
  AND2X2 U107 ( .A(\InC<12> ), .B(n66), .Y(n95) );
  INVX1 U108 ( .A(n95), .Y(n96) );
  AND2X2 U109 ( .A(\InD<3> ), .B(n126), .Y(n97) );
  INVX1 U110 ( .A(n97), .Y(n98) );
  INVX1 U111 ( .A(n125), .Y(n99) );
  INVX1 U112 ( .A(n99), .Y(n100) );
  INVX1 U113 ( .A(n127), .Y(n101) );
  INVX1 U114 ( .A(n101), .Y(n102) );
  INVX1 U115 ( .A(n134), .Y(n103) );
  INVX1 U116 ( .A(n103), .Y(n104) );
  INVX1 U117 ( .A(n136), .Y(n105) );
  INVX1 U118 ( .A(n105), .Y(n106) );
  INVX1 U119 ( .A(n138), .Y(n107) );
  INVX1 U120 ( .A(n107), .Y(n108) );
  INVX1 U121 ( .A(n140), .Y(n109) );
  INVX1 U122 ( .A(n109), .Y(n110) );
  INVX1 U123 ( .A(n141), .Y(n111) );
  INVX1 U124 ( .A(n111), .Y(n112) );
  INVX1 U125 ( .A(n143), .Y(n113) );
  INVX1 U126 ( .A(n113), .Y(n114) );
  INVX1 U127 ( .A(n148), .Y(n115) );
  INVX1 U128 ( .A(n115), .Y(n116) );
  INVX1 U129 ( .A(n151), .Y(n117) );
  INVX1 U130 ( .A(n117), .Y(n118) );
  AOI22X1 U131 ( .A(n126), .B(\InD<0> ), .C(n149), .D(\InA<0> ), .Y(n122) );
  INVX1 U132 ( .A(\S<1> ), .Y(n120) );
  INVX1 U133 ( .A(\S<0> ), .Y(n121) );
  INVX4 U134 ( .A(n65), .Y(n150) );
  INVX8 U135 ( .A(n124), .Y(n149) );
  OR2X2 U136 ( .A(\S<1> ), .B(\S<0> ), .Y(n124) );
  NAND3X1 U137 ( .A(n58), .B(n36), .C(n61), .Y(\Out<0> ) );
  AOI22X1 U138 ( .A(\InB<1> ), .B(n150), .C(\InA<1> ), .D(n149), .Y(n125) );
  NAND3X1 U139 ( .A(n38), .B(n5), .C(n100), .Y(n165) );
  AOI22X1 U140 ( .A(\InB<2> ), .B(n150), .C(\InA<2> ), .D(n149), .Y(n127) );
  NAND3X1 U141 ( .A(n40), .B(n7), .C(n102), .Y(n164) );
  AOI22X1 U142 ( .A(\InB<3> ), .B(n150), .C(\InA<3> ), .D(n149), .Y(n128) );
  NAND3X1 U143 ( .A(n42), .B(n98), .C(n59), .Y(n163) );
  AOI22X1 U144 ( .A(\InB<4> ), .B(n150), .C(\InA<4> ), .D(n149), .Y(n130) );
  NAND3X1 U145 ( .A(n72), .B(n9), .C(n70), .Y(n162) );
  AOI22X1 U146 ( .A(\InB<5> ), .B(n150), .C(\InA<5> ), .D(n149), .Y(n132) );
  NAND3X1 U147 ( .A(n74), .B(n11), .C(n76), .Y(n161) );
  AOI22X1 U148 ( .A(\InB<6> ), .B(n150), .C(\InA<6> ), .D(n149), .Y(n134) );
  NAND3X1 U149 ( .A(n44), .B(n13), .C(n104), .Y(n160) );
  AOI22X1 U150 ( .A(\InB<7> ), .B(n150), .C(\InA<7> ), .D(n149), .Y(n136) );
  NAND3X1 U151 ( .A(n46), .B(n15), .C(n106), .Y(n159) );
  AOI22X1 U152 ( .A(\InB<8> ), .B(n150), .C(\InA<8> ), .D(n149), .Y(n138) );
  NAND3X1 U153 ( .A(n48), .B(n17), .C(n108), .Y(n158) );
  AOI22X1 U154 ( .A(\InB<9> ), .B(n150), .C(\InA<9> ), .D(n149), .Y(n140) );
  NAND3X1 U155 ( .A(n50), .B(n19), .C(n110), .Y(n157) );
  AOI22X1 U156 ( .A(\InB<10> ), .B(n150), .C(\InA<10> ), .D(n149), .Y(n141) );
  NAND3X1 U157 ( .A(n52), .B(n21), .C(n112), .Y(n156) );
  AOI22X1 U158 ( .A(\InB<11> ), .B(n150), .C(\InA<11> ), .D(n149), .Y(n143) );
  NAND3X1 U159 ( .A(n54), .B(n23), .C(n114), .Y(n155) );
  AOI22X1 U160 ( .A(\InB<12> ), .B(n150), .C(\InA<12> ), .D(n149), .Y(n145) );
  NAND3X1 U161 ( .A(n96), .B(n25), .C(n78), .Y(n154) );
  AOI22X1 U162 ( .A(\InB<13> ), .B(n150), .C(\InA<13> ), .D(n149), .Y(n147) );
  AOI22X1 U163 ( .A(\InB<14> ), .B(n150), .C(\InA<14> ), .D(n149), .Y(n148) );
  NAND3X1 U164 ( .A(n56), .B(n29), .C(n116), .Y(n153) );
  AOI22X1 U165 ( .A(\InB<15> ), .B(n150), .C(\InA<15> ), .D(n149), .Y(n151) );
  NAND3X1 U166 ( .A(n31), .B(n33), .C(n118), .Y(n152) );
endmodule


module cla16_1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13;

  cla4_7 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_6 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n13), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_5 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n12), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_4 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n11), .S({\S<15> , \S<14> , \S<13> , \S<12> }), .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  INVX1 U1 ( .A(n3), .Y(n11) );
  INVX1 U2 ( .A(n11), .Y(n9) );
  BUFX2 U3 ( .A(n4), .Y(n1) );
  BUFX2 U4 ( .A(n5), .Y(n2) );
  BUFX2 U5 ( .A(n6), .Y(n3) );
  INVX1 U6 ( .A(\G<3> ), .Y(n7) );
  INVX1 U7 ( .A(\P<3> ), .Y(n8) );
  AOI21X1 U8 ( .A(Cin), .B(\P<0> ), .C(\G<0> ), .Y(n4) );
  INVX2 U9 ( .A(n1), .Y(n13) );
  AOI21X1 U10 ( .A(\P<1> ), .B(n13), .C(\G<1> ), .Y(n5) );
  INVX2 U11 ( .A(n2), .Y(n12) );
  AOI21X1 U12 ( .A(\P<2> ), .B(n12), .C(\G<2> ), .Y(n6) );
  OAI21X1 U13 ( .A(n9), .B(n8), .C(n7), .Y(Cout) );
endmodule


module mux4to1 ( InA, InB, InC, InD, .S({\S<1> , \S<0> }), Out );
  input InA, InB, InC, InD, \S<1> , \S<0> ;
  output Out;
  wire   n1, n2;

  MUX2X1 U1 ( .B(InA), .A(InC), .S(\S<1> ), .Y(n2) );
  MUX2X1 U2 ( .B(InB), .A(InD), .S(\S<1> ), .Y(n1) );
  MUX2X1 U3 ( .B(n2), .A(n1), .S(\S<0> ), .Y(Out) );
endmodule


module memory2c_0 ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, \mem<0><7> , \mem<0><6> ,
         \mem<0><5> , \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> ,
         \mem<0><0> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> ,
         \mem<2><6> , \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> ,
         \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> ,
         \mem<4><7> , \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> ,
         \mem<4><2> , \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> ,
         \mem<5><5> , \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> ,
         \mem<5><0> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> ,
         \mem<7><6> , \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> ,
         \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> ,
         \mem<9><7> , \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> ,
         \mem<9><2> , \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> ,
         \mem<10><5> , \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> ,
         \mem<10><0> , \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> ,
         \mem<11><3> , \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> ,
         \mem<12><6> , \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> ,
         \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> ,
         \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> ,
         \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> ,
         \mem<17><6> , \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> ,
         \mem<18><4> , \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> ,
         \mem<19><7> , \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> ,
         \mem<19><2> , \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> ,
         \mem<20><5> , \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> ,
         \mem<20><0> , \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> ,
         \mem<21><3> , \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> ,
         \mem<22><6> , \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> ,
         \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> ,
         \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> ,
         \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> ,
         \mem<27><6> , \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> ,
         \mem<28><4> , \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> ,
         \mem<29><7> , \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> ,
         \mem<29><2> , \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> ,
         \mem<30><5> , \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> ,
         \mem<30><0> , \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> ,
         \mem<31><3> , \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> ,
         \mem<32><6> , \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> ,
         \mem<32><1> , \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> ,
         \mem<33><4> , \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> ,
         \mem<34><7> , \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> ,
         \mem<34><2> , \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> ,
         \mem<35><5> , \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> ,
         \mem<35><0> , \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> ,
         \mem<36><3> , \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> ,
         \mem<37><6> , \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> ,
         \mem<37><1> , \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> ,
         \mem<38><4> , \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> ,
         \mem<39><7> , \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> ,
         \mem<39><2> , \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> ,
         \mem<40><5> , \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> ,
         \mem<40><0> , \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> ,
         \mem<41><3> , \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> ,
         \mem<42><6> , \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> ,
         \mem<42><1> , \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> ,
         \mem<43><4> , \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> ,
         \mem<44><7> , \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> ,
         \mem<44><2> , \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> ,
         \mem<45><5> , \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> ,
         \mem<45><0> , \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> ,
         \mem<46><3> , \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> ,
         \mem<47><6> , \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> ,
         \mem<47><1> , \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> ,
         \mem<48><4> , \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> ,
         \mem<49><7> , \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> ,
         \mem<49><2> , \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> ,
         \mem<50><5> , \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> ,
         \mem<50><0> , \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> ,
         \mem<51><3> , \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> ,
         \mem<52><6> , \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> ,
         \mem<52><1> , \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> ,
         \mem<53><4> , \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> ,
         \mem<54><7> , \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> ,
         \mem<54><2> , \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> ,
         \mem<55><5> , \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> ,
         \mem<55><0> , \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> ,
         \mem<56><3> , \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> ,
         \mem<57><6> , \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> ,
         \mem<57><1> , \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> ,
         \mem<58><4> , \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> ,
         \mem<59><7> , \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> ,
         \mem<59><2> , \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> ,
         \mem<60><5> , \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> ,
         \mem<60><0> , \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> ,
         \mem<61><3> , \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> ,
         \mem<62><6> , \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> ,
         \mem<62><1> , \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> ,
         \mem<63><4> , \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n769, n770, n771, n772,
         n773, n775, n776, n777, n778, n780, n782, n783, n784, n786, n787,
         n788, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n6429), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n6430), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n6431), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n6432), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n6433), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n6434), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n6435), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n6436), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n6437), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n6438), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n6439), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n6440), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n6441), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n6442), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n6443), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n6444), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n6445), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n6446), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n6447), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n6448), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n6449), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n6450), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n6451), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n6452), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n6453), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n6454), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n6455), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n6456), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n6457), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n6458), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n6459), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n6460), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n6461), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n6462), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n6463), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n6464), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n6465), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n6466), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n6467), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n6468), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n6469), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n6470), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n6471), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n6472), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n6473), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n6474), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n6475), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n6476), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n6477), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n6478), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n6479), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n6480), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n6481), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n6482), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n6483), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n6484), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n6485), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n6486), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n6487), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n6488), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n6489), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n6490), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n6491), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n6492), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n6493), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n6494), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n6495), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n6496), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n6497), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n6498), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n6499), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n6500), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n6501), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n6502), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n6503), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n6504), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n6505), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n6506), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n6507), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n6508), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n6509), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n6510), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n6511), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n6512), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n6513), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n6514), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n6515), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n6516), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n6517), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n6518), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n6519), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n6520), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n6521), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n6522), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n6523), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n6524), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n6525), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n6526), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n6527), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n6528), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n6529), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n6530), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n6531), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n6532), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n6533), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n6534), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n6535), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n6536), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n6537), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n6538), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n6539), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n6540), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n6541), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n6542), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n6543), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n6544), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n6545), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n6546), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n6547), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n6548), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n6549), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n6550), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n6551), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n6552), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n6553), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n6554), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n6555), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n6556), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n6557), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n6558), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n6559), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n6560), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n6561), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n6562), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n6563), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n6564), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n6565), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n6566), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n6567), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n6568), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n6569), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n6570), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n6571), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n6572), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n6573), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n6574), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n6575), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n6576), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n6577), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n6578), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n6579), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n6580), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n6581), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n6582), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n6583), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n6584), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n6585), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n6586), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n6587), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n6588), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n6589), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n6590), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n6591), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n6592), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n6593), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n6594), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n6595), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n6596), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n6597), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n6598), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n6599), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n6600), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n6601), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n6602), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n6603), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n6604), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n6605), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n6606), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n6607), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n6608), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n6609), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n6610), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n6611), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n6612), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n6613), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n6614), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n6615), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n6616), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n6617), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n6618), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n6619), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n6620), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n6621), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n6622), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n6623), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n6624), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n6625), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n6626), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n6627), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n6628), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n6629), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n6630), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n6631), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n6632), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n6633), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n6634), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n6635), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n6636), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n6637), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n6638), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n6639), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n6640), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n6641), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n6642), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n6643), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n6644), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n6645), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n6646), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n6647), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n6648), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n6649), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n6650), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n6651), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n6652), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n6653), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n6654), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n6655), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n6656), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n6657), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n6658), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n6659), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n6660), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n6661), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n6662), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n6663), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n6664), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n6665), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n6666), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n6667), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n6668), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n6669), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n6670), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n6671), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n6672), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n6673), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n6674), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n6675), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n6676), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n6677), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n6678), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n6679), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n6680), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n6681), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n6682), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n6683), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n6684), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n6685), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n6686), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n6687), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n6688), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n6689), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n6690), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n6691), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n6692), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n6693), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n6694), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n6695), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n6696), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n6697), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n6698), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n6699), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n6700), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n6701), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n6702), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n6703), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n6704), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n6705), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n6706), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n6707), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n6708), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n6709), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n6710), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n6711), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n6712), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n6713), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n6714), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n6715), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n6716), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n6717), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n6718), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n6719), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n6720), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n6721), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n6722), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n6723), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n6724), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n6725), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n6726), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n6727), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n6728), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n6729), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n6730), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n6731), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n6732), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n6733), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n6734), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n6735), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n6736), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n6737), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n6738), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n6739), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n6740), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n6741), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n6742), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n6743), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n6744), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n6745), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n6746), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n6747), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n6748), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n6749), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n6750), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n6751), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n6752), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n6753), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n6754), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n6755), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n6756), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n6757), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n6758), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n6759), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n6760), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n6761), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n6762), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n6763), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n6764), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n6765), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n6766), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n6767), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n6768), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n6769), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n6770), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n6771), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n6772), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n6773), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n6774), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n6775), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n6776), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n6777), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n6778), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n6779), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n6780), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n6781), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n6782), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n6783), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n6784), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n6785), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n6786), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n6787), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n6788), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n6789), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n6790), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n6791), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n6792), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n6793), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n6794), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n6795), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n6796), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n6797), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n6798), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n6799), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n6800), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n6801), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n6802), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n6803), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n6804), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n6805), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n6806), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n6807), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n6808), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n6809), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n6810), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n6811), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n6812), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n6813), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n6814), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n6815), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n6816), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n6817), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n6818), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n6819), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n6820), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n6821), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n6822), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n6823), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n6824), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n6825), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n6826), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n6827), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n6828), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n6829), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n6830), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n6831), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n6832), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n6833), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n6834), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n6835), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n6836), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n6837), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n6838), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n6839), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n6840), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n6841), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n6842), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n6843), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n6844), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n6845), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n6846), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n6847), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n6848), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n6849), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n6850), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n6851), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n6852), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n6853), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n6854), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n6855), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n6856), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n6857), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n6858), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n6859), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n6860), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n6861), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n6862), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n6863), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n6864), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n6865), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n6866), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n6867), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n6868), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n6869), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n6870), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n6871), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n6872), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n6873), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n6874), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n6875), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n6876), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n6877), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n6878), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n6879), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n6880), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n6881), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n6882), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n6883), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n6884), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n6885), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n6886), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n6887), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n6888), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n6889), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n6890), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n6891), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n6892), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n6893), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n6894), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n6895), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n6896), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n6897), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n6898), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n6899), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n6900), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n6901), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n6902), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n6903), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n6904), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n6905), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n6906), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n6907), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n6908), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n6909), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n6910), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n6911), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n6912), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n6913), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n6914), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n6915), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n6916), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n6917), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n6918), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n6919), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n6920), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n6921), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n6922), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n6923), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n6924), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n6925), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n6926), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n6927), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n6928), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n6929), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n6930), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n6931), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n6932), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n6933), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n6934), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n6935), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n6936), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n6937), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n6938), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n6939), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n6940), .CLK(clk), .Q(\mem<63><0> ) );
  INVX1 U3 ( .A(n4861), .Y(n1) );
  BUFX2 U4 ( .A(\addr<8> ), .Y(n2) );
  INVX1 U5 ( .A(n3660), .Y(n3) );
  INVX2 U6 ( .A(n3660), .Y(n3661) );
  INVX2 U7 ( .A(n3660), .Y(n4964) );
  INVX4 U8 ( .A(n3654), .Y(n4829) );
  INVX1 U9 ( .A(n4841), .Y(n3851) );
  OR2X2 U10 ( .A(n651), .B(n648), .Y(n647) );
  INVX2 U11 ( .A(N177), .Y(n4867) );
  INVX1 U12 ( .A(n3665), .Y(n4) );
  AND2X2 U13 ( .A(n87), .B(n4), .Y(n5) );
  INVX2 U14 ( .A(n44), .Y(n3873) );
  AND2X2 U15 ( .A(n6287), .B(n86), .Y(n6) );
  OR2X2 U16 ( .A(n3572), .B(n4978), .Y(n7) );
  INVX1 U17 ( .A(n6407), .Y(n8) );
  INVX1 U18 ( .A(n6337), .Y(n9) );
  INVX1 U19 ( .A(n6306), .Y(n10) );
  INVX1 U20 ( .A(n6341), .Y(n6340) );
  INVX1 U21 ( .A(n6412), .Y(n6411) );
  INVX1 U22 ( .A(n6310), .Y(n6309) );
  INVX1 U23 ( .A(n3631), .Y(n11) );
  INVX2 U24 ( .A(n3615), .Y(n3616) );
  INVX1 U25 ( .A(n4658), .Y(n12) );
  INVX2 U26 ( .A(n3585), .Y(n3586) );
  INVX1 U27 ( .A(n4856), .Y(n13) );
  INVX1 U28 ( .A(n4856), .Y(n4826) );
  INVX1 U29 ( .A(n97), .Y(n14) );
  INVX2 U30 ( .A(n3625), .Y(n3626) );
  INVX1 U31 ( .A(n4957), .Y(n15) );
  INVX1 U32 ( .A(n955), .Y(n16) );
  INVX2 U33 ( .A(n3637), .Y(n3638) );
  INVX1 U34 ( .A(n4812), .Y(n17) );
  INVX1 U35 ( .A(n6365), .Y(n18) );
  INVX1 U36 ( .A(n4632), .Y(n19) );
  INVX2 U37 ( .A(n3869), .Y(n6397) );
  AND2X2 U38 ( .A(n3856), .B(n3619), .Y(n20) );
  AND2X2 U39 ( .A(n4875), .B(n3585), .Y(n21) );
  INVX2 U40 ( .A(n3609), .Y(n3610) );
  INVX2 U41 ( .A(n3621), .Y(n3622) );
  INVX2 U42 ( .A(n3866), .Y(n6370) );
  INVX8 U43 ( .A(n4960), .Y(n4957) );
  INVX2 U44 ( .A(n3597), .Y(n3598) );
  INVX2 U45 ( .A(n574), .Y(n6330) );
  INVX1 U46 ( .A(n18), .Y(n22) );
  INVX1 U47 ( .A(n48), .Y(n23) );
  INVX1 U48 ( .A(n18), .Y(n49) );
  INVX1 U49 ( .A(n48), .Y(n24) );
  BUFX2 U50 ( .A(n6348), .Y(n4929) );
  INVX1 U51 ( .A(n6328), .Y(n25) );
  INVX1 U52 ( .A(n4629), .Y(n26) );
  INVX1 U53 ( .A(n1685), .Y(n27) );
  INVX2 U54 ( .A(n1685), .Y(n6329) );
  AND2X2 U55 ( .A(n4966), .B(n4858), .Y(n28) );
  INVX2 U56 ( .A(n29), .Y(n6359) );
  INVX1 U57 ( .A(n6354), .Y(n30) );
  OAI21X1 U58 ( .A(n4650), .B(n30), .C(n6417), .Y(n29) );
  BUFX2 U59 ( .A(n29), .Y(n4932) );
  INVX1 U60 ( .A(n3667), .Y(n31) );
  INVX1 U61 ( .A(n31), .Y(n32) );
  INVX1 U62 ( .A(n31), .Y(n33) );
  INVX1 U63 ( .A(n31), .Y(n34) );
  INVX1 U64 ( .A(n952), .Y(n35) );
  INVX1 U65 ( .A(n4917), .Y(n36) );
  INVX1 U66 ( .A(n3561), .Y(n37) );
  OR2X2 U67 ( .A(n39), .B(n6371), .Y(n38) );
  INVX8 U68 ( .A(\mem<22><0> ), .Y(n39) );
  AND2X2 U69 ( .A(n4680), .B(n3605), .Y(n40) );
  AND2X2 U70 ( .A(n4674), .B(n3587), .Y(n41) );
  INVX2 U71 ( .A(n3583), .Y(n3584) );
  INVX4 U72 ( .A(n3617), .Y(n3618) );
  AND2X2 U73 ( .A(n3873), .B(n3595), .Y(n42) );
  INVX2 U74 ( .A(n3623), .Y(n3624) );
  INVX1 U75 ( .A(n3660), .Y(n43) );
  INVX1 U76 ( .A(n43), .Y(n44) );
  INVX2 U77 ( .A(n3656), .Y(n3849) );
  INVX1 U78 ( .A(n4865), .Y(n45) );
  INVX1 U79 ( .A(n3674), .Y(n46) );
  AND2X2 U80 ( .A(n6366), .B(n3617), .Y(n47) );
  INVX1 U81 ( .A(n6365), .Y(n48) );
  AND2X2 U82 ( .A(n4674), .B(n6364), .Y(n50) );
  INVX1 U83 ( .A(n6365), .Y(n6364) );
  INVX2 U84 ( .A(n46), .Y(n4674) );
  INVX1 U85 ( .A(n6372), .Y(n51) );
  AND2X2 U86 ( .A(n3712), .B(n4853), .Y(n52) );
  AND2X2 U87 ( .A(n4674), .B(n3645), .Y(n53) );
  INVX1 U88 ( .A(n6373), .Y(n6371) );
  BUFX2 U89 ( .A(n6351), .Y(n4930) );
  INVX1 U90 ( .A(n4841), .Y(n54) );
  INVX1 U91 ( .A(n4841), .Y(n55) );
  INVX1 U92 ( .A(n2), .Y(n56) );
  INVX1 U93 ( .A(n56), .Y(n57) );
  INVX1 U94 ( .A(n4944), .Y(n58) );
  INVX1 U95 ( .A(n579), .Y(n59) );
  INVX8 U96 ( .A(n4945), .Y(n4944) );
  INVX1 U97 ( .A(n562), .Y(n60) );
  INVX1 U98 ( .A(n562), .Y(n61) );
  INVX1 U99 ( .A(n562), .Y(n4819) );
  AND2X2 U100 ( .A(n1049), .B(n1062), .Y(n1241) );
  OR2X2 U101 ( .A(n1257), .B(n1258), .Y(n62) );
  BUFX2 U102 ( .A(n3874), .Y(n4882) );
  INVX1 U103 ( .A(n4966), .Y(n63) );
  INVX1 U104 ( .A(n63), .Y(n64) );
  INVX1 U105 ( .A(n115), .Y(n65) );
  INVX1 U106 ( .A(n4980), .Y(n4817) );
  BUFX2 U107 ( .A(n3874), .Y(n4881) );
  MUX2X1 U108 ( .B(n6128), .A(n6127), .S(n4881), .Y(n6159) );
  INVX2 U109 ( .A(n4840), .Y(n4841) );
  AND2X2 U110 ( .A(n4778), .B(n4779), .Y(n5435) );
  INVX1 U111 ( .A(n745), .Y(n66) );
  INVX8 U112 ( .A(\data_in<8> ), .Y(n5076) );
  INVX4 U113 ( .A(n5063), .Y(n5060) );
  INVX8 U114 ( .A(\data_in<10> ), .Y(n5086) );
  INVX4 U115 ( .A(N180), .Y(n5009) );
  INVX8 U116 ( .A(n5130), .Y(n4946) );
  INVX2 U117 ( .A(n578), .Y(n4949) );
  INVX4 U118 ( .A(n5012), .Y(n5021) );
  OR2X2 U119 ( .A(n104), .B(n5748), .Y(n67) );
  INVX4 U120 ( .A(n3673), .Y(n4816) );
  INVX2 U121 ( .A(n4682), .Y(n4719) );
  INVX2 U122 ( .A(n814), .Y(n93) );
  INVX4 U123 ( .A(n3577), .Y(n3578) );
  INVX2 U124 ( .A(n3653), .Y(n3654) );
  OR2X2 U125 ( .A(n4750), .B(n6370), .Y(n68) );
  INVX4 U126 ( .A(n3668), .Y(n3669) );
  OR2X2 U127 ( .A(n6388), .B(n5634), .Y(n69) );
  OR2X2 U128 ( .A(n6388), .B(n5469), .Y(n70) );
  INVX2 U129 ( .A(n3613), .Y(n3614) );
  OR2X2 U130 ( .A(n4734), .B(n4850), .Y(n71) );
  AND2X1 U131 ( .A(n4944), .B(n5171), .Y(n1272) );
  AND2X1 U132 ( .A(n4944), .B(n5337), .Y(n1276) );
  AND2X1 U133 ( .A(n3880), .B(\mem<33><2> ), .Y(n1153) );
  INVX1 U134 ( .A(\mem<37><7> ), .Y(n5741) );
  INVX1 U135 ( .A(\mem<39><0> ), .Y(n5152) );
  INVX1 U136 ( .A(\mem<37><0> ), .Y(n5162) );
  INVX1 U137 ( .A(\mem<35><0> ), .Y(n5135) );
  INVX1 U138 ( .A(\mem<48><6> ), .Y(n5691) );
  INVX1 U139 ( .A(\mem<35><6> ), .Y(n5642) );
  INVX1 U140 ( .A(\mem<39><6> ), .Y(n5656) );
  INVX1 U141 ( .A(\mem<37><6> ), .Y(n5666) );
  INVX1 U142 ( .A(\mem<35><2> ), .Y(n5305) );
  INVX1 U143 ( .A(\mem<39><2> ), .Y(n5319) );
  INVX1 U144 ( .A(\mem<37><2> ), .Y(n5329) );
  INVX1 U145 ( .A(\mem<35><3> ), .Y(n5393) );
  INVX1 U146 ( .A(\mem<37><3> ), .Y(n5417) );
  INVX1 U147 ( .A(\mem<39><3> ), .Y(n5406) );
  INVX1 U148 ( .A(\mem<8><7> ), .Y(n5714) );
  INVX1 U149 ( .A(\mem<35><1> ), .Y(n5246) );
  INVX1 U150 ( .A(\mem<39><1> ), .Y(n5258) );
  INVX1 U151 ( .A(\mem<37><1> ), .Y(n5268) );
  INVX1 U152 ( .A(\mem<41><0> ), .Y(n5193) );
  INVX1 U153 ( .A(\mem<1><0> ), .Y(n5145) );
  INVX1 U154 ( .A(\mem<43><6> ), .Y(n5637) );
  INVX1 U155 ( .A(\mem<38><2> ), .Y(n5344) );
  INVX1 U156 ( .A(\mem<34><3> ), .Y(n5454) );
  INVX1 U157 ( .A(\mem<4><3> ), .Y(n5451) );
  INVX1 U158 ( .A(\mem<35><4> ), .Y(n5477) );
  INVX1 U159 ( .A(\mem<37><4> ), .Y(n5500) );
  INVX1 U160 ( .A(\mem<39><4> ), .Y(n5491) );
  INVX1 U161 ( .A(\mem<35><5> ), .Y(n5560) );
  INVX1 U162 ( .A(\mem<39><5> ), .Y(n5574) );
  INVX1 U163 ( .A(\mem<37><5> ), .Y(n5584) );
  INVX1 U164 ( .A(\mem<36><1> ), .Y(n5236) );
  INVX1 U165 ( .A(\mem<38><1> ), .Y(n5281) );
  INVX1 U166 ( .A(\mem<24><0> ), .Y(n5189) );
  INVX1 U167 ( .A(\mem<34><6> ), .Y(n5703) );
  INVX1 U168 ( .A(\mem<34><2> ), .Y(n5294) );
  INVX1 U169 ( .A(\mem<43><4> ), .Y(n5472) );
  INVX1 U170 ( .A(\mem<43><5> ), .Y(n5555) );
  INVX1 U171 ( .A(\mem<24><1> ), .Y(n5213) );
  INVX1 U172 ( .A(n5093), .Y(n5087) );
  INVX1 U173 ( .A(n5092), .Y(n5088) );
  INVX1 U174 ( .A(\data_in<9> ), .Y(n5081) );
  INVX1 U175 ( .A(\data_in<11> ), .Y(n5091) );
  INVX1 U176 ( .A(\data_in<14> ), .Y(n5106) );
  AND2X1 U177 ( .A(n4897), .B(n5149), .Y(n3896) );
  AND2X1 U178 ( .A(n4903), .B(n5159), .Y(n3900) );
  AND2X1 U179 ( .A(n4896), .B(n5653), .Y(n3942) );
  AND2X1 U180 ( .A(n4898), .B(n5663), .Y(n3944) );
  INVX1 U181 ( .A(\mem<46><6> ), .Y(n5674) );
  AND2X1 U182 ( .A(n4905), .B(n5326), .Y(n1151) );
  AND2X1 U183 ( .A(n4890), .B(n5389), .Y(n1157) );
  AND2X1 U184 ( .A(n121), .B(n5403), .Y(n1159) );
  INVX1 U185 ( .A(\mem<39><7> ), .Y(n5733) );
  AND2X1 U186 ( .A(n4892), .B(n5255), .Y(n1143) );
  INVX1 U187 ( .A(\mem<38><0> ), .Y(n5177) );
  INVX1 U188 ( .A(\mem<14><0> ), .Y(n5174) );
  INVX1 U189 ( .A(\mem<43><0> ), .Y(n5128) );
  INVX1 U190 ( .A(\mem<21><6> ), .Y(n564) );
  INVX1 U191 ( .A(\mem<41><2> ), .Y(n5356) );
  INVX1 U192 ( .A(\mem<25><2> ), .Y(n5357) );
  INVX1 U193 ( .A(\mem<56><2> ), .Y(n5354) );
  INVX1 U194 ( .A(\mem<46><3> ), .Y(n5426) );
  AND2X1 U195 ( .A(n4904), .B(n5474), .Y(n1165) );
  AND2X1 U196 ( .A(n4906), .B(n5557), .Y(n1175) );
  AND2X1 U197 ( .A(n812), .B(n5142), .Y(n5143) );
  AND2X1 U198 ( .A(n4892), .B(n5570), .Y(n1177) );
  AND2X1 U199 ( .A(n4905), .B(n5581), .Y(n1179) );
  INVX1 U200 ( .A(\mem<57><7> ), .Y(n5748) );
  INVX1 U201 ( .A(\mem<41><7> ), .Y(n5747) );
  INVX1 U202 ( .A(n5245), .Y(n559) );
  INVX1 U203 ( .A(\mem<19><1> ), .Y(n558) );
  INVX1 U204 ( .A(\mem<33><0> ), .Y(n4833) );
  INVX1 U205 ( .A(\mem<47><0> ), .Y(n5147) );
  INVX1 U206 ( .A(\mem<45><0> ), .Y(n5157) );
  INVX1 U207 ( .A(\mem<12><0> ), .Y(n5169) );
  INVX1 U208 ( .A(\mem<48><0> ), .Y(n5170) );
  INVX1 U209 ( .A(\mem<36><0> ), .Y(n5121) );
  INVX1 U210 ( .A(\mem<34><0> ), .Y(n5119) );
  INVX1 U211 ( .A(\mem<36><6> ), .Y(n5688) );
  INVX1 U212 ( .A(\mem<20><6> ), .Y(n5692) );
  INVX1 U213 ( .A(\mem<42><6> ), .Y(n5695) );
  INVX1 U214 ( .A(\mem<26><6> ), .Y(n5705) );
  INVX1 U215 ( .A(\mem<45><6> ), .Y(n5661) );
  INVX1 U216 ( .A(\mem<47><6> ), .Y(n5651) );
  INVX1 U217 ( .A(\mem<17><6> ), .Y(n5634) );
  INVX1 U218 ( .A(\mem<8><6> ), .Y(n5631) );
  INVX1 U219 ( .A(\mem<50><6> ), .Y(n5629) );
  INVX1 U220 ( .A(\mem<36><2> ), .Y(n5295) );
  INVX1 U221 ( .A(\mem<14><2> ), .Y(n5340) );
  INVX1 U222 ( .A(\mem<43><2> ), .Y(n5300) );
  INVX1 U223 ( .A(\mem<1><2> ), .Y(n5311) );
  INVX1 U224 ( .A(\mem<47><2> ), .Y(n5313) );
  INVX1 U225 ( .A(\mem<45><2> ), .Y(n5324) );
  INVX1 U226 ( .A(\mem<2><2> ), .Y(n5370) );
  INVX1 U227 ( .A(\mem<52><2> ), .Y(n5368) );
  INVX1 U228 ( .A(\mem<4><2> ), .Y(n4852) );
  INVX1 U229 ( .A(\mem<48><3> ), .Y(n5444) );
  INVX1 U230 ( .A(\mem<12><3> ), .Y(n567) );
  INVX1 U231 ( .A(\mem<43><3> ), .Y(n5387) );
  INVX1 U232 ( .A(\mem<1><3> ), .Y(n5399) );
  INVX1 U233 ( .A(\mem<45><3> ), .Y(n5411) );
  INVX1 U234 ( .A(\mem<47><3> ), .Y(n5401) );
  INVX1 U235 ( .A(\mem<8><3> ), .Y(n5384) );
  INVX1 U236 ( .A(\mem<46><4> ), .Y(n5509) );
  INVX1 U237 ( .A(\mem<23><4> ), .Y(n110) );
  INVX1 U238 ( .A(\mem<34><5> ), .Y(n5620) );
  INVX1 U239 ( .A(\mem<20><5> ), .Y(n5609) );
  INVX1 U240 ( .A(\mem<12><7> ), .Y(n4837) );
  INVX1 U241 ( .A(\mem<20><7> ), .Y(n5763) );
  INVX1 U242 ( .A(\mem<56><7> ), .Y(n4886) );
  INVX1 U243 ( .A(\mem<9><7> ), .Y(n5719) );
  INVX1 U244 ( .A(\mem<50><7> ), .Y(n5712) );
  INVX1 U245 ( .A(\mem<41><1> ), .Y(n5216) );
  INVX1 U246 ( .A(\mem<56><1> ), .Y(n5215) );
  INVX1 U247 ( .A(\mem<57><1> ), .Y(n5226) );
  INVX1 U248 ( .A(\mem<2><1> ), .Y(n5225) );
  INVX1 U249 ( .A(\mem<14><1> ), .Y(n5278) );
  INVX1 U250 ( .A(\mem<43><1> ), .Y(n5241) );
  INVX1 U251 ( .A(\mem<1><1> ), .Y(n5251) );
  INVX1 U252 ( .A(\mem<47><1> ), .Y(n5253) );
  INVX1 U253 ( .A(\mem<45><1> ), .Y(n5263) );
  INVX1 U254 ( .A(\mem<56><0> ), .Y(n5191) );
  INVX1 U255 ( .A(\mem<57><0> ), .Y(n5204) );
  INVX1 U256 ( .A(\mem<2><0> ), .Y(n5202) );
  INVX1 U257 ( .A(n5146), .Y(n556) );
  INVX1 U258 ( .A(\mem<60><0> ), .Y(n5117) );
  INVX1 U259 ( .A(\mem<4><6> ), .Y(n5700) );
  INVX1 U260 ( .A(\mem<1><6> ), .Y(n5648) );
  INVX1 U261 ( .A(\mem<9><6> ), .Y(n5627) );
  INVX1 U262 ( .A(\mem<60><2> ), .Y(n5292) );
  INVX1 U263 ( .A(\mem<12><2> ), .Y(n5335) );
  INVX1 U264 ( .A(\mem<48><2> ), .Y(n5336) );
  INVX1 U265 ( .A(\mem<50><2> ), .Y(n5365) );
  INVX1 U266 ( .A(\mem<26><2> ), .Y(n5363) );
  INVX1 U267 ( .A(\mem<36><3> ), .Y(n5440) );
  INVX1 U268 ( .A(\mem<16><3> ), .Y(n570) );
  INVX1 U269 ( .A(\mem<41><3> ), .Y(n5423) );
  INVX1 U270 ( .A(\mem<57><3> ), .Y(n5432) );
  INVX1 U271 ( .A(\mem<56><3> ), .Y(n5376) );
  INVX1 U272 ( .A(\mem<9><3> ), .Y(n5378) );
  INVX1 U273 ( .A(\mem<4><4> ), .Y(n5531) );
  INVX1 U274 ( .A(\mem<34><4> ), .Y(n5534) );
  INVX1 U275 ( .A(\mem<45><4> ), .Y(n5495) );
  INVX1 U276 ( .A(\mem<47><4> ), .Y(n5485) );
  INVX1 U277 ( .A(\mem<17><4> ), .Y(n5469) );
  INVX1 U278 ( .A(\mem<8><4> ), .Y(n5466) );
  INVX1 U279 ( .A(\mem<50><4> ), .Y(n5464) );
  INVX1 U280 ( .A(\mem<42><5> ), .Y(n5612) );
  INVX1 U281 ( .A(\mem<47><5> ), .Y(n5568) );
  INVX1 U282 ( .A(\mem<45><5> ), .Y(n5579) );
  INVX1 U283 ( .A(\mem<9><5> ), .Y(n5543) );
  INVX1 U284 ( .A(\mem<8><5> ), .Y(n5548) );
  INVX1 U285 ( .A(\mem<50><5> ), .Y(n5546) );
  INVX1 U286 ( .A(\mem<42><7> ), .Y(n106) );
  INVX1 U287 ( .A(n5766), .Y(n107) );
  INVX1 U288 ( .A(\mem<36><7> ), .Y(n5767) );
  INVX1 U289 ( .A(\mem<4><7> ), .Y(n5778) );
  INVX2 U290 ( .A(n6335), .Y(n4956) );
  INVX1 U291 ( .A(\mem<49><1> ), .Y(n5223) );
  INVX1 U292 ( .A(\mem<34><1> ), .Y(n5234) );
  INVX1 U293 ( .A(\mem<60><1> ), .Y(n5232) );
  INVX1 U294 ( .A(\mem<12><1> ), .Y(n5273) );
  INVX1 U295 ( .A(\mem<48><1> ), .Y(n5274) );
  INVX1 U296 ( .A(\mem<20><4> ), .Y(n5524) );
  INVX1 U297 ( .A(\mem<36><4> ), .Y(n5520) );
  INVX1 U298 ( .A(\mem<42><4> ), .Y(n5527) );
  INVX1 U299 ( .A(\mem<1><4> ), .Y(n5483) );
  INVX1 U300 ( .A(\mem<36><5> ), .Y(n5605) );
  INVX1 U301 ( .A(\mem<4><5> ), .Y(n5617) );
  INVX1 U302 ( .A(\mem<1><5> ), .Y(n5566) );
  INVX1 U303 ( .A(\mem<17><5> ), .Y(n5551) );
  INVX1 U304 ( .A(n6306), .Y(n6308) );
  INVX1 U305 ( .A(n6337), .Y(n6339) );
  INVX1 U306 ( .A(n6407), .Y(n6409) );
  INVX1 U307 ( .A(n4922), .Y(n6297) );
  INVX1 U308 ( .A(n84), .Y(n6302) );
  INVX1 U309 ( .A(n6348), .Y(n6346) );
  INVX1 U310 ( .A(n6351), .Y(n6349) );
  INVX1 U311 ( .A(n4935), .Y(n6375) );
  INVX1 U312 ( .A(n4937), .Y(n6395) );
  INVX1 U313 ( .A(n6392), .Y(n6394) );
  INVX2 U314 ( .A(n59), .Y(n6399) );
  INVX1 U315 ( .A(n5086), .Y(n5083) );
  INVX1 U316 ( .A(\mem<0><0> ), .Y(n6420) );
  INVX1 U317 ( .A(\mem<0><1> ), .Y(n6421) );
  INVX1 U318 ( .A(\mem<0><2> ), .Y(n6422) );
  INVX1 U319 ( .A(\mem<0><3> ), .Y(n6423) );
  INVX1 U320 ( .A(\mem<0><4> ), .Y(n6424) );
  INVX1 U321 ( .A(\mem<0><5> ), .Y(n6425) );
  INVX1 U322 ( .A(\mem<0><6> ), .Y(n6426) );
  INVX1 U323 ( .A(\mem<0><7> ), .Y(n6428) );
  INVX8 U324 ( .A(\data_in<12> ), .Y(n5097) );
  INVX8 U325 ( .A(\data_in<13> ), .Y(n5101) );
  INVX8 U326 ( .A(\data_in<7> ), .Y(n5071) );
  INVX8 U327 ( .A(\data_in<0> ), .Y(n5040) );
  INVX2 U328 ( .A(n5022), .Y(n5035) );
  INVX1 U329 ( .A(n5068), .Y(n5064) );
  INVX1 U330 ( .A(n5068), .Y(n5065) );
  INVX4 U331 ( .A(n4982), .Y(n4993) );
  INVX1 U332 ( .A(n5050), .Y(n5048) );
  INVX1 U333 ( .A(n5050), .Y(n5047) );
  INVX1 U334 ( .A(n5050), .Y(n5049) );
  INVX1 U335 ( .A(n5059), .Y(n5055) );
  INVX1 U336 ( .A(n5059), .Y(n5056) );
  INVX1 U337 ( .A(n4975), .Y(n3870) );
  INVX1 U338 ( .A(n5054), .Y(n5051) );
  INVX1 U339 ( .A(n5054), .Y(n5053) );
  INVX2 U340 ( .A(\data_in<9> ), .Y(n5080) );
  INVX1 U341 ( .A(n4982), .Y(n4996) );
  INVX2 U342 ( .A(n5022), .Y(n5034) );
  INVX2 U343 ( .A(n5062), .Y(n5061) );
  INVX2 U344 ( .A(n5067), .Y(n5066) );
  INVX1 U345 ( .A(\data_in<11> ), .Y(n5092) );
  INVX1 U346 ( .A(\data_in<11> ), .Y(n5093) );
  INVX2 U347 ( .A(\data_in<14> ), .Y(n5105) );
  INVX1 U348 ( .A(N178), .Y(n4983) );
  INVX1 U349 ( .A(n4983), .Y(n4982) );
  AND2X2 U350 ( .A(\mem<54><3> ), .B(n4948), .Y(n72) );
  AND2X2 U351 ( .A(\mem<54><5> ), .B(n4948), .Y(n73) );
  AND2X2 U352 ( .A(\mem<19><7> ), .B(n4957), .Y(n74) );
  AND2X2 U353 ( .A(\mem<51><7> ), .B(n4851), .Y(n75) );
  AND2X2 U354 ( .A(\mem<54><4> ), .B(n4948), .Y(n76) );
  AND2X2 U355 ( .A(\mem<54><6> ), .B(n4848), .Y(n77) );
  INVX1 U356 ( .A(\addr<15> ), .Y(n5134) );
  INVX1 U357 ( .A(n4889), .Y(n4893) );
  INVX1 U358 ( .A(n4627), .Y(n5192) );
  INVX2 U359 ( .A(n5115), .Y(n4853) );
  INVX1 U360 ( .A(n3650), .Y(n6389) );
  INVX1 U361 ( .A(n806), .Y(n4681) );
  INVX2 U362 ( .A(n5058), .Y(n5057) );
  INVX1 U363 ( .A(n5110), .Y(n5109) );
  INVX1 U364 ( .A(n5097), .Y(n5096) );
  INVX1 U365 ( .A(n5101), .Y(n5100) );
  INVX1 U366 ( .A(n5105), .Y(n5104) );
  INVX1 U367 ( .A(n5092), .Y(n5090) );
  INVX1 U368 ( .A(n5080), .Y(n5079) );
  INVX1 U369 ( .A(n5086), .Y(n5085) );
  INVX1 U370 ( .A(n5076), .Y(n5075) );
  INVX4 U371 ( .A(n7), .Y(n6427) );
  INVX2 U372 ( .A(n3593), .Y(n3594) );
  INVX2 U373 ( .A(n6418), .Y(n6419) );
  INVX2 U374 ( .A(n3579), .Y(n3580) );
  INVX1 U375 ( .A(n819), .Y(n78) );
  INVX1 U376 ( .A(n819), .Y(n4879) );
  AND2X2 U377 ( .A(n6287), .B(n79), .Y(n1688) );
  AND2X2 U378 ( .A(n4974), .B(n6289), .Y(n79) );
  BUFX2 U379 ( .A(n4775), .Y(n80) );
  INVX1 U380 ( .A(n80), .Y(n81) );
  INVX1 U381 ( .A(n80), .Y(n82) );
  INVX1 U382 ( .A(n80), .Y(n4972) );
  AND2X2 U383 ( .A(n122), .B(n52), .Y(n83) );
  AND2X2 U384 ( .A(n122), .B(n52), .Y(n84) );
  INVX2 U385 ( .A(n3619), .Y(n3620) );
  INVX2 U386 ( .A(n3591), .Y(n3592) );
  INVX1 U387 ( .A(n3631), .Y(n85) );
  INVX2 U388 ( .A(n4823), .Y(n4911) );
  INVX1 U389 ( .A(n3631), .Y(n3632) );
  INVX1 U390 ( .A(n6354), .Y(n6358) );
  AND2X2 U391 ( .A(n4974), .B(n3873), .Y(n86) );
  INVX1 U392 ( .A(n6324), .Y(n4952) );
  BUFX2 U393 ( .A(n6296), .Y(n4921) );
  INVX2 U394 ( .A(n6296), .Y(n87) );
  INVX1 U395 ( .A(n954), .Y(n88) );
  INVX1 U396 ( .A(n1031), .Y(n89) );
  INVX1 U397 ( .A(n4859), .Y(n90) );
  BUFX2 U398 ( .A(n3612), .Y(n91) );
  BUFX2 U399 ( .A(n3612), .Y(n92) );
  INVX1 U400 ( .A(n792), .Y(n94) );
  BUFX2 U401 ( .A(n6295), .Y(n4920) );
  INVX1 U402 ( .A(n93), .Y(n95) );
  INVX1 U403 ( .A(n95), .Y(n96) );
  INVX1 U404 ( .A(n3862), .Y(n97) );
  INVX2 U405 ( .A(n3595), .Y(n3596) );
  INVX1 U406 ( .A(n6372), .Y(n6374) );
  INVX2 U407 ( .A(n3627), .Y(n3628) );
  AND2X2 U408 ( .A(n6098), .B(n5846), .Y(\data_out<12> ) );
  BUFX2 U409 ( .A(n6307), .Y(n4924) );
  BUFX2 U410 ( .A(n6412), .Y(n4939) );
  BUFX2 U411 ( .A(n6341), .Y(n4928) );
  BUFX2 U412 ( .A(n6301), .Y(n4923) );
  BUFX2 U413 ( .A(n6408), .Y(n4938) );
  BUFX2 U414 ( .A(n6373), .Y(n4934) );
  BUFX2 U415 ( .A(n6338), .Y(n4927) );
  BUFX2 U416 ( .A(n6327), .Y(n4926) );
  BUFX2 U417 ( .A(n6393), .Y(n4936) );
  INVX1 U418 ( .A(n4694), .Y(n5846) );
  INVX1 U419 ( .A(n4981), .Y(n99) );
  INVX1 U420 ( .A(n4841), .Y(n114) );
  INVX1 U421 ( .A(n776), .Y(n100) );
  BUFX2 U422 ( .A(n6293), .Y(n4919) );
  INVX1 U423 ( .A(n4839), .Y(n101) );
  AND2X2 U424 ( .A(n4965), .B(n3633), .Y(n102) );
  INVX1 U425 ( .A(n4861), .Y(n103) );
  BUFX2 U426 ( .A(n3652), .Y(n104) );
  INVX8 U427 ( .A(n4846), .Y(n6342) );
  OAI21X1 U428 ( .A(n106), .B(n6332), .C(n107), .Y(n105) );
  INVX1 U429 ( .A(n78), .Y(n108) );
  INVX1 U430 ( .A(n6415), .Y(n555) );
  INVX1 U431 ( .A(n5489), .Y(n111) );
  OAI21X1 U432 ( .A(n110), .B(n4854), .C(n111), .Y(n109) );
  INVX4 U433 ( .A(n4957), .Y(n4854) );
  BUFX2 U434 ( .A(n6410), .Y(n112) );
  INVX4 U435 ( .A(n803), .Y(n804) );
  BUFX4 U436 ( .A(n4945), .Y(n113) );
  AND2X2 U437 ( .A(n4738), .B(n4739), .Y(n5683) );
  INVX1 U438 ( .A(n4840), .Y(n115) );
  INVX1 U439 ( .A(n44), .Y(n4965) );
  INVX4 U440 ( .A(n4883), .Y(n5037) );
  INVX8 U441 ( .A(n5037), .Y(n5031) );
  INVX8 U442 ( .A(n5037), .Y(n5032) );
  INVX1 U443 ( .A(n798), .Y(n116) );
  INVX1 U444 ( .A(n4839), .Y(n117) );
  INVX1 U445 ( .A(n4859), .Y(n118) );
  INVX1 U446 ( .A(n745), .Y(n119) );
  INVX1 U447 ( .A(n5112), .Y(n576) );
  INVX1 U448 ( .A(n3568), .Y(n120) );
  INVX1 U449 ( .A(n4816), .Y(n571) );
  INVX8 U450 ( .A(n3712), .Y(n4945) );
  INVX1 U451 ( .A(n4944), .Y(n4943) );
  INVX1 U452 ( .A(n5023), .Y(n5022) );
  INVX4 U453 ( .A(N182), .Y(n4885) );
  INVX1 U454 ( .A(n4889), .Y(n121) );
  AND2X2 U455 ( .A(n4865), .B(n5203), .Y(n122) );
  NOR3X1 U456 ( .A(n3854), .B(n800), .C(n101), .Y(n123) );
  INVX1 U457 ( .A(n123), .Y(n6335) );
  INVX1 U458 ( .A(n154), .Y(n124) );
  INVX1 U459 ( .A(n4956), .Y(n125) );
  INVX1 U460 ( .A(n4672), .Y(n126) );
  INVX1 U461 ( .A(n4888), .Y(n127) );
  INVX1 U462 ( .A(n6324), .Y(n128) );
  INVX1 U463 ( .A(n128), .Y(n129) );
  INVX1 U464 ( .A(n128), .Y(n130) );
  INVX1 U465 ( .A(n128), .Y(n131) );
  INVX1 U466 ( .A(n4859), .Y(n132) );
  INVX1 U467 ( .A(n132), .Y(n133) );
  INVX1 U468 ( .A(n132), .Y(n134) );
  INVX1 U469 ( .A(n132), .Y(n135) );
  INVX1 U470 ( .A(n3845), .Y(n136) );
  INVX1 U471 ( .A(n136), .Y(n137) );
  INVX1 U472 ( .A(n136), .Y(n138) );
  INVX1 U473 ( .A(n3845), .Y(n139) );
  INVX1 U474 ( .A(n139), .Y(n140) );
  INVX1 U475 ( .A(n139), .Y(n141) );
  INVX1 U476 ( .A(n151), .Y(n142) );
  INVX1 U477 ( .A(n90), .Y(n143) );
  INVX1 U478 ( .A(n118), .Y(n144) );
  INVX1 U479 ( .A(n118), .Y(n145) );
  INVX1 U480 ( .A(n143), .Y(n146) );
  INVX1 U481 ( .A(n143), .Y(n147) );
  INVX1 U482 ( .A(n144), .Y(n148) );
  INVX1 U483 ( .A(n144), .Y(n149) );
  INVX1 U484 ( .A(n145), .Y(n150) );
  INVX1 U485 ( .A(n145), .Y(n151) );
  INVX1 U486 ( .A(n4951), .Y(n152) );
  INVX1 U487 ( .A(n5751), .Y(n6324) );
  INVX1 U488 ( .A(n4952), .Y(n4951) );
  INVX1 U489 ( .A(n125), .Y(n153) );
  NOR3X1 U490 ( .A(n4981), .B(n580), .C(n15), .Y(n154) );
  INVX1 U491 ( .A(n154), .Y(n4823) );
  INVX1 U492 ( .A(n5203), .Y(n580) );
  INVX8 U493 ( .A(n4963), .Y(n4961) );
  AND2X2 U494 ( .A(n5134), .B(n2354), .Y(n155) );
  OR2X2 U495 ( .A(n4852), .B(n6414), .Y(n156) );
  AND2X2 U496 ( .A(\mem<38><3> ), .B(n4954), .Y(n157) );
  AND2X2 U497 ( .A(\mem<6><3> ), .B(n4838), .Y(n158) );
  AND2X2 U498 ( .A(\mem<38><4> ), .B(n4954), .Y(n159) );
  AND2X2 U499 ( .A(\mem<38><5> ), .B(n4954), .Y(n160) );
  AND2X2 U500 ( .A(\mem<38><6> ), .B(n4954), .Y(n161) );
  AND2X2 U501 ( .A(\mem<35><7> ), .B(n4954), .Y(n162) );
  AND2X2 U502 ( .A(\mem<3><7> ), .B(n4838), .Y(n163) );
  AND2X2 U503 ( .A(\mem<52><0> ), .B(n4877), .Y(n164) );
  INVX1 U504 ( .A(n164), .Y(n165) );
  AND2X2 U505 ( .A(\mem<50><0> ), .B(n3668), .Y(n166) );
  INVX1 U506 ( .A(n166), .Y(n167) );
  AND2X2 U507 ( .A(\mem<52><1> ), .B(n4877), .Y(n168) );
  INVX1 U508 ( .A(n168), .Y(n169) );
  AND2X2 U509 ( .A(\mem<50><1> ), .B(n3668), .Y(n170) );
  INVX1 U510 ( .A(n170), .Y(n171) );
  AND2X2 U511 ( .A(\mem<40><1> ), .B(n4680), .Y(n172) );
  INVX1 U512 ( .A(n172), .Y(n173) );
  AND2X2 U513 ( .A(\mem<44><2> ), .B(n574), .Y(n174) );
  INVX1 U514 ( .A(n174), .Y(n175) );
  AND2X2 U515 ( .A(\mem<18><2> ), .B(n577), .Y(n176) );
  INVX1 U516 ( .A(n176), .Y(n177) );
  AND2X2 U517 ( .A(\mem<53><7> ), .B(n4949), .Y(n178) );
  INVX1 U518 ( .A(n178), .Y(n179) );
  AND2X2 U519 ( .A(\mem<22><7> ), .B(n4959), .Y(n180) );
  INVX1 U520 ( .A(n180), .Y(n181) );
  AND2X2 U521 ( .A(\mem<63><0> ), .B(n4692), .Y(n182) );
  INVX1 U522 ( .A(n182), .Y(n183) );
  AND2X2 U523 ( .A(\mem<63><1> ), .B(n4693), .Y(n184) );
  INVX1 U524 ( .A(n184), .Y(n185) );
  AND2X2 U525 ( .A(\mem<63><3> ), .B(n4693), .Y(n186) );
  INVX1 U526 ( .A(n186), .Y(n187) );
  AND2X2 U527 ( .A(\mem<63><4> ), .B(n4692), .Y(n188) );
  INVX1 U528 ( .A(n188), .Y(n189) );
  AND2X2 U529 ( .A(\mem<63><6> ), .B(n4692), .Y(n190) );
  INVX1 U530 ( .A(n190), .Y(n191) );
  AND2X2 U531 ( .A(\mem<63><7> ), .B(n4693), .Y(n192) );
  INVX1 U532 ( .A(n192), .Y(n193) );
  AND2X2 U533 ( .A(\mem<60><0> ), .B(n4921), .Y(n194) );
  INVX1 U534 ( .A(n194), .Y(n195) );
  AND2X2 U535 ( .A(\mem<60><1> ), .B(n4921), .Y(n196) );
  INVX1 U536 ( .A(n196), .Y(n197) );
  AND2X2 U537 ( .A(\mem<60><2> ), .B(n4921), .Y(n198) );
  INVX1 U538 ( .A(n198), .Y(n199) );
  AND2X2 U539 ( .A(\mem<60><3> ), .B(n4921), .Y(n200) );
  INVX1 U540 ( .A(n200), .Y(n201) );
  AND2X2 U541 ( .A(\mem<60><4> ), .B(n4921), .Y(n202) );
  INVX1 U542 ( .A(n202), .Y(n203) );
  AND2X2 U543 ( .A(\mem<60><5> ), .B(n4921), .Y(n204) );
  INVX1 U544 ( .A(n204), .Y(n205) );
  AND2X2 U545 ( .A(\mem<60><6> ), .B(n4921), .Y(n206) );
  INVX1 U546 ( .A(n206), .Y(n207) );
  AND2X2 U547 ( .A(\mem<60><7> ), .B(n4921), .Y(n208) );
  INVX1 U548 ( .A(n208), .Y(n209) );
  AND2X2 U549 ( .A(\mem<59><0> ), .B(n4922), .Y(n210) );
  INVX1 U550 ( .A(n210), .Y(n211) );
  AND2X2 U551 ( .A(\mem<59><1> ), .B(n4922), .Y(n212) );
  INVX1 U552 ( .A(n212), .Y(n213) );
  AND2X2 U553 ( .A(\mem<59><2> ), .B(n4922), .Y(n214) );
  INVX1 U554 ( .A(n214), .Y(n215) );
  AND2X2 U555 ( .A(\mem<59><3> ), .B(n4922), .Y(n216) );
  INVX1 U556 ( .A(n216), .Y(n217) );
  AND2X2 U557 ( .A(\mem<59><4> ), .B(n4922), .Y(n218) );
  INVX1 U558 ( .A(n218), .Y(n219) );
  AND2X2 U559 ( .A(\mem<59><5> ), .B(n4922), .Y(n220) );
  INVX1 U560 ( .A(n220), .Y(n221) );
  AND2X2 U561 ( .A(\mem<59><6> ), .B(n4922), .Y(n222) );
  INVX1 U562 ( .A(n222), .Y(n223) );
  AND2X2 U563 ( .A(\mem<59><7> ), .B(n4922), .Y(n224) );
  INVX1 U564 ( .A(n224), .Y(n225) );
  AND2X2 U565 ( .A(\mem<56><4> ), .B(n3582), .Y(n226) );
  INVX1 U566 ( .A(n226), .Y(n227) );
  AND2X2 U567 ( .A(\mem<55><4> ), .B(n3584), .Y(n228) );
  INVX1 U568 ( .A(n228), .Y(n229) );
  AND2X2 U569 ( .A(\mem<52><4> ), .B(n3586), .Y(n230) );
  INVX1 U570 ( .A(n230), .Y(n231) );
  AND2X2 U571 ( .A(\mem<51><4> ), .B(n3588), .Y(n232) );
  INVX1 U572 ( .A(n232), .Y(n233) );
  AND2X2 U573 ( .A(\mem<49><0> ), .B(n3592), .Y(n234) );
  INVX1 U574 ( .A(n234), .Y(n235) );
  AND2X2 U575 ( .A(\mem<47><4> ), .B(n3596), .Y(n236) );
  INVX1 U576 ( .A(n236), .Y(n237) );
  AND2X2 U577 ( .A(\mem<41><4> ), .B(n3604), .Y(n238) );
  INVX1 U578 ( .A(n238), .Y(n239) );
  AND2X2 U579 ( .A(\mem<36><4> ), .B(n3610), .Y(n240) );
  INVX1 U580 ( .A(n240), .Y(n241) );
  AND2X2 U581 ( .A(\mem<35><4> ), .B(n92), .Y(n242) );
  INVX1 U582 ( .A(n242), .Y(n243) );
  AND2X2 U583 ( .A(\mem<33><4> ), .B(n3616), .Y(n244) );
  INVX1 U584 ( .A(n244), .Y(n245) );
  AND2X2 U585 ( .A(\mem<31><0> ), .B(n4930), .Y(n246) );
  INVX1 U586 ( .A(n246), .Y(n247) );
  AND2X2 U587 ( .A(\mem<31><1> ), .B(n4930), .Y(n248) );
  INVX1 U588 ( .A(n248), .Y(n249) );
  AND2X2 U589 ( .A(\mem<31><2> ), .B(n4930), .Y(n250) );
  INVX1 U590 ( .A(n250), .Y(n251) );
  AND2X2 U591 ( .A(\mem<31><3> ), .B(n4930), .Y(n252) );
  INVX1 U592 ( .A(n252), .Y(n253) );
  AND2X2 U593 ( .A(\mem<31><4> ), .B(n4930), .Y(n254) );
  INVX1 U594 ( .A(n254), .Y(n255) );
  AND2X2 U595 ( .A(\mem<31><5> ), .B(n4930), .Y(n256) );
  INVX1 U596 ( .A(n256), .Y(n257) );
  AND2X2 U597 ( .A(\mem<31><6> ), .B(n4930), .Y(n258) );
  INVX1 U598 ( .A(n258), .Y(n259) );
  AND2X2 U599 ( .A(\mem<31><7> ), .B(n4930), .Y(n260) );
  INVX1 U600 ( .A(n260), .Y(n261) );
  AND2X2 U601 ( .A(\mem<30><0> ), .B(n4931), .Y(n262) );
  INVX1 U602 ( .A(n262), .Y(n263) );
  AND2X2 U603 ( .A(\mem<30><1> ), .B(n4931), .Y(n264) );
  INVX1 U604 ( .A(n264), .Y(n265) );
  AND2X2 U605 ( .A(\mem<30><2> ), .B(n4931), .Y(n266) );
  INVX1 U606 ( .A(n266), .Y(n267) );
  AND2X2 U607 ( .A(\mem<30><3> ), .B(n4931), .Y(n268) );
  INVX1 U608 ( .A(n268), .Y(n269) );
  AND2X2 U609 ( .A(\mem<30><4> ), .B(n4931), .Y(n270) );
  INVX1 U610 ( .A(n270), .Y(n271) );
  AND2X2 U611 ( .A(\mem<30><5> ), .B(n4931), .Y(n272) );
  INVX1 U612 ( .A(n272), .Y(n273) );
  AND2X2 U613 ( .A(\mem<30><6> ), .B(n4931), .Y(n274) );
  INVX1 U614 ( .A(n274), .Y(n275) );
  AND2X2 U615 ( .A(\mem<30><7> ), .B(n4931), .Y(n276) );
  INVX1 U616 ( .A(n276), .Y(n277) );
  BUFX2 U617 ( .A(n6357), .Y(n4931) );
  AND2X2 U618 ( .A(\mem<29><4> ), .B(n29), .Y(n278) );
  INVX1 U619 ( .A(n278), .Y(n279) );
  AND2X2 U620 ( .A(\mem<26><4> ), .B(n3618), .Y(n280) );
  INVX1 U621 ( .A(n280), .Y(n281) );
  AND2X2 U622 ( .A(\mem<23><4> ), .B(n3624), .Y(n282) );
  INVX1 U623 ( .A(n282), .Y(n283) );
  AND2X2 U624 ( .A(\mem<20><4> ), .B(n3626), .Y(n284) );
  INVX1 U625 ( .A(n284), .Y(n285) );
  AND2X2 U626 ( .A(\mem<15><4> ), .B(n3634), .Y(n286) );
  INVX1 U627 ( .A(n286), .Y(n287) );
  AND2X2 U628 ( .A(\mem<12><4> ), .B(n6397), .Y(n288) );
  INVX1 U629 ( .A(n288), .Y(n289) );
  AND2X2 U630 ( .A(\mem<11><0> ), .B(n34), .Y(n290) );
  INVX1 U631 ( .A(n290), .Y(n291) );
  AND2X2 U632 ( .A(\mem<11><1> ), .B(n33), .Y(n292) );
  INVX1 U633 ( .A(n292), .Y(n293) );
  AND2X2 U634 ( .A(\mem<11><2> ), .B(n32), .Y(n294) );
  INVX1 U635 ( .A(n294), .Y(n295) );
  AND2X2 U636 ( .A(\mem<11><3> ), .B(n32), .Y(n296) );
  INVX1 U637 ( .A(n296), .Y(n297) );
  AND2X2 U638 ( .A(\mem<11><4> ), .B(n32), .Y(n298) );
  INVX1 U639 ( .A(n298), .Y(n299) );
  AND2X2 U640 ( .A(\mem<4><4> ), .B(n3644), .Y(n300) );
  INVX1 U641 ( .A(n300), .Y(n301) );
  AND2X2 U642 ( .A(\mem<3><4> ), .B(n3646), .Y(n302) );
  INVX1 U643 ( .A(n302), .Y(n303) );
  AND2X2 U644 ( .A(\mem<63><3> ), .B(n4946), .Y(n304) );
  INVX1 U645 ( .A(n304), .Y(n305) );
  AND2X2 U646 ( .A(\mem<59><6> ), .B(n4946), .Y(n306) );
  INVX1 U647 ( .A(n306), .Y(n307) );
  AND2X2 U648 ( .A(\mem<57><7> ), .B(n3580), .Y(n308) );
  INVX1 U649 ( .A(n308), .Y(n309) );
  AND2X2 U650 ( .A(\mem<56><0> ), .B(n3582), .Y(n310) );
  INVX1 U651 ( .A(n310), .Y(n311) );
  AND2X2 U652 ( .A(\mem<56><1> ), .B(n3582), .Y(n312) );
  INVX1 U653 ( .A(n312), .Y(n313) );
  AND2X2 U654 ( .A(\mem<56><2> ), .B(n3582), .Y(n314) );
  INVX1 U655 ( .A(n314), .Y(n315) );
  AND2X2 U656 ( .A(\mem<56><3> ), .B(n3582), .Y(n316) );
  INVX1 U657 ( .A(n316), .Y(n317) );
  AND2X2 U658 ( .A(\mem<56><5> ), .B(n3582), .Y(n318) );
  INVX1 U659 ( .A(n318), .Y(n319) );
  AND2X2 U660 ( .A(\mem<56><6> ), .B(n3582), .Y(n320) );
  INVX1 U661 ( .A(n320), .Y(n321) );
  AND2X2 U662 ( .A(\mem<56><7> ), .B(n3582), .Y(n322) );
  INVX1 U663 ( .A(n322), .Y(n323) );
  AND2X2 U664 ( .A(\mem<55><0> ), .B(n3584), .Y(n324) );
  INVX1 U665 ( .A(n324), .Y(n325) );
  AND2X2 U666 ( .A(\mem<55><1> ), .B(n3584), .Y(n326) );
  INVX1 U667 ( .A(n326), .Y(n327) );
  AND2X2 U668 ( .A(\mem<55><2> ), .B(n3584), .Y(n328) );
  INVX1 U669 ( .A(n328), .Y(n329) );
  AND2X2 U670 ( .A(\mem<55><3> ), .B(n3584), .Y(n330) );
  INVX1 U671 ( .A(n330), .Y(n331) );
  AND2X2 U672 ( .A(\mem<55><5> ), .B(n3584), .Y(n332) );
  INVX1 U673 ( .A(n332), .Y(n333) );
  AND2X2 U674 ( .A(\mem<55><6> ), .B(n3584), .Y(n334) );
  INVX1 U675 ( .A(n334), .Y(n335) );
  AND2X2 U676 ( .A(\mem<55><7> ), .B(n3584), .Y(n336) );
  INVX1 U677 ( .A(n336), .Y(n337) );
  AND2X2 U678 ( .A(\mem<52><0> ), .B(n3586), .Y(n338) );
  INVX1 U679 ( .A(n338), .Y(n339) );
  AND2X2 U680 ( .A(\mem<52><1> ), .B(n3586), .Y(n340) );
  INVX1 U681 ( .A(n340), .Y(n341) );
  AND2X2 U682 ( .A(\mem<52><2> ), .B(n3586), .Y(n342) );
  INVX1 U683 ( .A(n342), .Y(n343) );
  AND2X2 U684 ( .A(\mem<52><3> ), .B(n3586), .Y(n344) );
  INVX1 U685 ( .A(n344), .Y(n345) );
  AND2X2 U686 ( .A(\mem<52><5> ), .B(n3586), .Y(n346) );
  INVX1 U687 ( .A(n346), .Y(n347) );
  AND2X2 U688 ( .A(\mem<52><6> ), .B(n3586), .Y(n348) );
  INVX1 U689 ( .A(n348), .Y(n349) );
  AND2X2 U690 ( .A(\mem<52><7> ), .B(n3586), .Y(n350) );
  INVX1 U691 ( .A(n350), .Y(n351) );
  AND2X2 U692 ( .A(\mem<51><0> ), .B(n3588), .Y(n352) );
  INVX1 U693 ( .A(n352), .Y(n353) );
  AND2X2 U694 ( .A(\mem<51><1> ), .B(n3588), .Y(n354) );
  INVX1 U695 ( .A(n354), .Y(n355) );
  AND2X2 U696 ( .A(\mem<51><2> ), .B(n3588), .Y(n356) );
  INVX1 U697 ( .A(n356), .Y(n357) );
  AND2X2 U698 ( .A(\mem<51><3> ), .B(n3588), .Y(n358) );
  INVX1 U699 ( .A(n358), .Y(n359) );
  AND2X2 U700 ( .A(\mem<51><5> ), .B(n3588), .Y(n360) );
  INVX1 U701 ( .A(n360), .Y(n361) );
  AND2X2 U702 ( .A(\mem<51><6> ), .B(n3588), .Y(n362) );
  INVX1 U703 ( .A(n362), .Y(n363) );
  AND2X2 U704 ( .A(\mem<51><7> ), .B(n3588), .Y(n364) );
  INVX1 U705 ( .A(n364), .Y(n365) );
  AND2X2 U706 ( .A(\mem<47><0> ), .B(n3596), .Y(n366) );
  INVX1 U707 ( .A(n366), .Y(n367) );
  AND2X2 U708 ( .A(\mem<47><1> ), .B(n3596), .Y(n368) );
  INVX1 U709 ( .A(n368), .Y(n369) );
  AND2X2 U710 ( .A(\mem<47><2> ), .B(n3596), .Y(n370) );
  INVX1 U711 ( .A(n370), .Y(n371) );
  AND2X2 U712 ( .A(\mem<47><3> ), .B(n3596), .Y(n372) );
  INVX1 U713 ( .A(n372), .Y(n373) );
  AND2X2 U714 ( .A(\mem<47><5> ), .B(n3596), .Y(n374) );
  INVX1 U715 ( .A(n374), .Y(n375) );
  AND2X2 U716 ( .A(\mem<47><6> ), .B(n3596), .Y(n376) );
  INVX1 U717 ( .A(n376), .Y(n377) );
  AND2X2 U718 ( .A(\mem<47><7> ), .B(n3596), .Y(n378) );
  INVX1 U719 ( .A(n378), .Y(n379) );
  AND2X2 U720 ( .A(\mem<41><0> ), .B(n3604), .Y(n380) );
  INVX1 U721 ( .A(n380), .Y(n381) );
  AND2X2 U722 ( .A(\mem<41><1> ), .B(n3604), .Y(n382) );
  INVX1 U723 ( .A(n382), .Y(n383) );
  AND2X2 U724 ( .A(\mem<41><2> ), .B(n3604), .Y(n384) );
  INVX1 U725 ( .A(n384), .Y(n385) );
  AND2X2 U726 ( .A(\mem<41><3> ), .B(n3604), .Y(n386) );
  INVX1 U727 ( .A(n386), .Y(n387) );
  AND2X2 U728 ( .A(\mem<41><5> ), .B(n3604), .Y(n388) );
  INVX1 U729 ( .A(n388), .Y(n389) );
  AND2X2 U730 ( .A(\mem<41><6> ), .B(n3604), .Y(n390) );
  INVX1 U731 ( .A(n390), .Y(n391) );
  AND2X2 U732 ( .A(\mem<41><7> ), .B(n3604), .Y(n392) );
  INVX1 U733 ( .A(n392), .Y(n393) );
  AND2X2 U734 ( .A(\mem<36><0> ), .B(n3610), .Y(n394) );
  INVX1 U735 ( .A(n394), .Y(n395) );
  AND2X2 U736 ( .A(\mem<36><1> ), .B(n3610), .Y(n396) );
  INVX1 U737 ( .A(n396), .Y(n397) );
  AND2X2 U738 ( .A(\mem<36><2> ), .B(n3610), .Y(n398) );
  INVX1 U739 ( .A(n398), .Y(n399) );
  AND2X2 U740 ( .A(\mem<36><3> ), .B(n3610), .Y(n400) );
  INVX1 U741 ( .A(n400), .Y(n401) );
  AND2X2 U742 ( .A(\mem<36><5> ), .B(n3610), .Y(n402) );
  INVX1 U743 ( .A(n402), .Y(n403) );
  AND2X2 U744 ( .A(\mem<36><6> ), .B(n3610), .Y(n404) );
  INVX1 U745 ( .A(n404), .Y(n405) );
  AND2X2 U746 ( .A(\mem<36><7> ), .B(n3610), .Y(n406) );
  INVX1 U747 ( .A(n406), .Y(n407) );
  AND2X2 U748 ( .A(\mem<35><0> ), .B(n91), .Y(n408) );
  INVX1 U749 ( .A(n408), .Y(n409) );
  AND2X2 U750 ( .A(\mem<35><1> ), .B(n92), .Y(n410) );
  INVX1 U751 ( .A(n410), .Y(n411) );
  AND2X2 U752 ( .A(\mem<35><2> ), .B(n91), .Y(n412) );
  INVX1 U753 ( .A(n412), .Y(n413) );
  AND2X2 U754 ( .A(\mem<35><3> ), .B(n92), .Y(n414) );
  INVX1 U755 ( .A(n414), .Y(n415) );
  AND2X2 U756 ( .A(\mem<35><5> ), .B(n91), .Y(n416) );
  INVX1 U757 ( .A(n416), .Y(n417) );
  AND2X2 U758 ( .A(\mem<35><6> ), .B(n92), .Y(n418) );
  INVX1 U759 ( .A(n418), .Y(n419) );
  AND2X2 U760 ( .A(\mem<35><7> ), .B(n91), .Y(n420) );
  INVX1 U761 ( .A(n420), .Y(n421) );
  AND2X2 U762 ( .A(\mem<33><0> ), .B(n3616), .Y(n422) );
  INVX1 U763 ( .A(n422), .Y(n423) );
  AND2X2 U764 ( .A(\mem<33><1> ), .B(n3616), .Y(n424) );
  INVX1 U765 ( .A(n424), .Y(n425) );
  AND2X2 U766 ( .A(\mem<33><2> ), .B(n3616), .Y(n426) );
  INVX1 U767 ( .A(n426), .Y(n427) );
  AND2X2 U768 ( .A(\mem<33><3> ), .B(n3616), .Y(n428) );
  INVX1 U769 ( .A(n428), .Y(n429) );
  AND2X2 U770 ( .A(\mem<33><5> ), .B(n3616), .Y(n430) );
  INVX1 U771 ( .A(n430), .Y(n431) );
  AND2X2 U772 ( .A(\mem<33><6> ), .B(n3616), .Y(n432) );
  INVX1 U773 ( .A(n432), .Y(n433) );
  AND2X2 U774 ( .A(\mem<33><7> ), .B(n3616), .Y(n434) );
  INVX1 U775 ( .A(n434), .Y(n435) );
  AND2X2 U776 ( .A(\mem<29><0> ), .B(n29), .Y(n436) );
  INVX1 U777 ( .A(n436), .Y(n437) );
  AND2X2 U778 ( .A(\mem<29><1> ), .B(n29), .Y(n438) );
  INVX1 U779 ( .A(n438), .Y(n439) );
  AND2X2 U780 ( .A(\mem<29><2> ), .B(n4932), .Y(n440) );
  INVX1 U781 ( .A(n440), .Y(n441) );
  AND2X2 U782 ( .A(\mem<29><3> ), .B(n4932), .Y(n442) );
  INVX1 U783 ( .A(n442), .Y(n443) );
  AND2X2 U784 ( .A(\mem<29><5> ), .B(n4932), .Y(n444) );
  INVX1 U785 ( .A(n444), .Y(n445) );
  AND2X2 U786 ( .A(\mem<29><6> ), .B(n4932), .Y(n446) );
  INVX1 U787 ( .A(n446), .Y(n447) );
  AND2X2 U788 ( .A(\mem<29><7> ), .B(n4932), .Y(n448) );
  INVX1 U789 ( .A(n448), .Y(n449) );
  AND2X2 U790 ( .A(\mem<26><0> ), .B(n3618), .Y(n450) );
  INVX1 U791 ( .A(n450), .Y(n451) );
  AND2X2 U792 ( .A(\mem<26><1> ), .B(n3618), .Y(n452) );
  INVX1 U793 ( .A(n452), .Y(n453) );
  AND2X2 U794 ( .A(\mem<26><2> ), .B(n3618), .Y(n454) );
  INVX1 U795 ( .A(n454), .Y(n455) );
  AND2X2 U796 ( .A(\mem<26><3> ), .B(n3618), .Y(n456) );
  INVX1 U797 ( .A(n456), .Y(n457) );
  AND2X2 U798 ( .A(\mem<26><5> ), .B(n3618), .Y(n458) );
  INVX1 U799 ( .A(n458), .Y(n459) );
  AND2X2 U800 ( .A(\mem<26><6> ), .B(n3618), .Y(n460) );
  INVX1 U801 ( .A(n460), .Y(n461) );
  AND2X2 U802 ( .A(\mem<26><7> ), .B(n3618), .Y(n462) );
  INVX1 U803 ( .A(n462), .Y(n463) );
  AND2X2 U804 ( .A(\mem<23><0> ), .B(n3624), .Y(n464) );
  INVX1 U805 ( .A(n464), .Y(n465) );
  AND2X2 U806 ( .A(\mem<23><1> ), .B(n3624), .Y(n466) );
  INVX1 U807 ( .A(n466), .Y(n467) );
  AND2X2 U808 ( .A(\mem<23><2> ), .B(n3624), .Y(n468) );
  INVX1 U809 ( .A(n468), .Y(n469) );
  AND2X2 U810 ( .A(\mem<23><3> ), .B(n3624), .Y(n470) );
  INVX1 U811 ( .A(n470), .Y(n471) );
  AND2X2 U812 ( .A(\mem<23><5> ), .B(n3624), .Y(n472) );
  INVX1 U813 ( .A(n472), .Y(n473) );
  AND2X2 U814 ( .A(\mem<23><6> ), .B(n3624), .Y(n474) );
  INVX1 U815 ( .A(n474), .Y(n475) );
  AND2X2 U816 ( .A(\mem<23><7> ), .B(n3624), .Y(n476) );
  INVX1 U817 ( .A(n476), .Y(n477) );
  AND2X2 U818 ( .A(\mem<20><0> ), .B(n3626), .Y(n478) );
  INVX1 U819 ( .A(n478), .Y(n479) );
  AND2X2 U820 ( .A(\mem<20><1> ), .B(n3626), .Y(n480) );
  INVX1 U821 ( .A(n480), .Y(n481) );
  AND2X2 U822 ( .A(\mem<20><2> ), .B(n3626), .Y(n482) );
  INVX1 U823 ( .A(n482), .Y(n483) );
  AND2X2 U824 ( .A(\mem<20><3> ), .B(n3626), .Y(n484) );
  INVX1 U825 ( .A(n484), .Y(n485) );
  AND2X2 U826 ( .A(\mem<20><5> ), .B(n3626), .Y(n486) );
  INVX1 U827 ( .A(n486), .Y(n487) );
  AND2X2 U828 ( .A(\mem<20><6> ), .B(n3626), .Y(n488) );
  INVX1 U829 ( .A(n488), .Y(n489) );
  AND2X2 U830 ( .A(\mem<20><7> ), .B(n3626), .Y(n490) );
  INVX1 U831 ( .A(n490), .Y(n491) );
  AND2X2 U832 ( .A(\mem<15><0> ), .B(n3634), .Y(n492) );
  INVX1 U833 ( .A(n492), .Y(n493) );
  AND2X2 U834 ( .A(\mem<15><1> ), .B(n3634), .Y(n494) );
  INVX1 U835 ( .A(n494), .Y(n495) );
  AND2X2 U836 ( .A(\mem<15><2> ), .B(n3634), .Y(n496) );
  INVX1 U837 ( .A(n496), .Y(n497) );
  AND2X2 U838 ( .A(\mem<15><3> ), .B(n3634), .Y(n498) );
  INVX1 U839 ( .A(n498), .Y(n499) );
  AND2X2 U840 ( .A(\mem<15><5> ), .B(n3634), .Y(n500) );
  INVX1 U841 ( .A(n500), .Y(n501) );
  AND2X2 U842 ( .A(\mem<15><6> ), .B(n3634), .Y(n502) );
  INVX1 U843 ( .A(n502), .Y(n503) );
  AND2X2 U844 ( .A(\mem<15><7> ), .B(n3634), .Y(n504) );
  INVX1 U845 ( .A(n504), .Y(n505) );
  AND2X2 U846 ( .A(\mem<12><0> ), .B(n6397), .Y(n506) );
  INVX1 U847 ( .A(n506), .Y(n507) );
  AND2X2 U848 ( .A(\mem<12><1> ), .B(n6397), .Y(n508) );
  INVX1 U849 ( .A(n508), .Y(n509) );
  AND2X2 U850 ( .A(\mem<12><2> ), .B(n6397), .Y(n510) );
  INVX1 U851 ( .A(n510), .Y(n511) );
  AND2X2 U852 ( .A(\mem<12><3> ), .B(n6397), .Y(n512) );
  INVX1 U853 ( .A(n512), .Y(n513) );
  AND2X2 U854 ( .A(\mem<12><5> ), .B(n6397), .Y(n514) );
  INVX1 U855 ( .A(n514), .Y(n515) );
  AND2X2 U856 ( .A(\mem<12><6> ), .B(n6397), .Y(n516) );
  INVX1 U857 ( .A(n516), .Y(n517) );
  AND2X2 U858 ( .A(\mem<12><7> ), .B(n6397), .Y(n518) );
  INVX1 U859 ( .A(n518), .Y(n519) );
  AND2X2 U860 ( .A(\mem<11><5> ), .B(n33), .Y(n520) );
  INVX1 U861 ( .A(n520), .Y(n521) );
  AND2X2 U862 ( .A(\mem<11><6> ), .B(n34), .Y(n522) );
  INVX1 U863 ( .A(n522), .Y(n523) );
  AND2X2 U864 ( .A(\mem<11><7> ), .B(n33), .Y(n524) );
  INVX1 U865 ( .A(n524), .Y(n525) );
  AND2X2 U866 ( .A(\mem<4><0> ), .B(n3644), .Y(n526) );
  INVX1 U867 ( .A(n526), .Y(n527) );
  AND2X2 U868 ( .A(\mem<4><1> ), .B(n3644), .Y(n528) );
  INVX1 U869 ( .A(n528), .Y(n529) );
  AND2X2 U870 ( .A(\mem<4><2> ), .B(n3644), .Y(n530) );
  INVX1 U871 ( .A(n530), .Y(n531) );
  AND2X2 U872 ( .A(\mem<4><3> ), .B(n3644), .Y(n532) );
  INVX1 U873 ( .A(n532), .Y(n533) );
  AND2X2 U874 ( .A(\mem<4><5> ), .B(n3644), .Y(n534) );
  INVX1 U875 ( .A(n534), .Y(n535) );
  AND2X2 U876 ( .A(\mem<4><6> ), .B(n3644), .Y(n536) );
  INVX1 U877 ( .A(n536), .Y(n537) );
  AND2X2 U878 ( .A(\mem<4><7> ), .B(n3644), .Y(n538) );
  INVX1 U879 ( .A(n538), .Y(n539) );
  AND2X2 U880 ( .A(\mem<3><0> ), .B(n3646), .Y(n540) );
  INVX1 U881 ( .A(n540), .Y(n541) );
  AND2X2 U882 ( .A(\mem<3><1> ), .B(n3646), .Y(n542) );
  INVX1 U883 ( .A(n542), .Y(n543) );
  AND2X2 U884 ( .A(\mem<3><2> ), .B(n3646), .Y(n544) );
  INVX1 U885 ( .A(n544), .Y(n545) );
  AND2X2 U886 ( .A(\mem<3><3> ), .B(n3646), .Y(n546) );
  INVX1 U887 ( .A(n546), .Y(n547) );
  AND2X2 U888 ( .A(\mem<3><5> ), .B(n3646), .Y(n548) );
  INVX1 U889 ( .A(n548), .Y(n549) );
  AND2X2 U890 ( .A(\mem<3><6> ), .B(n3646), .Y(n550) );
  INVX1 U891 ( .A(n550), .Y(n551) );
  AND2X2 U892 ( .A(\mem<3><7> ), .B(n3646), .Y(n552) );
  INVX1 U893 ( .A(n552), .Y(n553) );
  AND2X2 U894 ( .A(n66), .B(\mem<42><3> ), .Y(n5442) );
  AND2X2 U895 ( .A(n4776), .B(n4777), .Y(n764) );
  OAI21X1 U896 ( .A(n555), .B(n594), .C(n556), .Y(n554) );
  INVX1 U897 ( .A(n554), .Y(n5185) );
  INVX1 U898 ( .A(n5664), .Y(n565) );
  OAI21X1 U899 ( .A(n558), .B(n4854), .C(n559), .Y(n557) );
  INVX1 U900 ( .A(n4861), .Y(n560) );
  INVX1 U901 ( .A(N177), .Y(n561) );
  AND2X2 U902 ( .A(n4866), .B(n5192), .Y(n562) );
  OAI21X1 U903 ( .A(n564), .B(n4854), .C(n565), .Y(n563) );
  INVX1 U904 ( .A(n4681), .Y(n566) );
  INVX1 U905 ( .A(n4681), .Y(n6304) );
  INVX1 U906 ( .A(n5452), .Y(n572) );
  OR2X2 U907 ( .A(n567), .B(n3653), .Y(n5443) );
  INVX2 U908 ( .A(n5036), .Y(n5030) );
  INVX1 U909 ( .A(n4883), .Y(n5036) );
  INVX1 U910 ( .A(N177), .Y(n568) );
  AND2X2 U911 ( .A(n3861), .B(n155), .Y(n6312) );
  INVX1 U912 ( .A(n805), .Y(n4839) );
  OAI21X1 U913 ( .A(n570), .B(n571), .C(n572), .Y(n569) );
  INVX1 U914 ( .A(n4754), .Y(n573) );
  INVX1 U915 ( .A(n4960), .Y(n4958) );
  INVX2 U916 ( .A(n4960), .Y(n4959) );
  NOR3X1 U917 ( .A(n130), .B(n5126), .C(n4841), .Y(n574) );
  NOR3X1 U918 ( .A(n576), .B(n2352), .C(n808), .Y(n575) );
  INVX1 U919 ( .A(n575), .Y(n4836) );
  INVX1 U920 ( .A(n124), .Y(n577) );
  AND2X2 U921 ( .A(n4789), .B(n614), .Y(n794) );
  INVX1 U922 ( .A(n6312), .Y(n578) );
  INVX4 U923 ( .A(n4950), .Y(n4873) );
  OR2X2 U924 ( .A(n4960), .B(n5126), .Y(n748) );
  INVX4 U925 ( .A(n4831), .Y(n4960) );
  INVX8 U926 ( .A(n4956), .Y(n4953) );
  NOR3X1 U927 ( .A(n4913), .B(n580), .C(n1687), .Y(n579) );
  INVX1 U928 ( .A(n579), .Y(n6400) );
  INVX2 U929 ( .A(n1687), .Y(n6398) );
  INVX1 U930 ( .A(n3665), .Y(n4887) );
  INVX4 U931 ( .A(n3664), .Y(n3665) );
  INVX2 U932 ( .A(n805), .Y(n3861) );
  INVX8 U933 ( .A(n6398), .Y(n4963) );
  INVX8 U934 ( .A(n3663), .Y(n6378) );
  INVX2 U935 ( .A(n3662), .Y(n3663) );
  INVX1 U936 ( .A(n3662), .Y(n6377) );
  OR2X2 U937 ( .A(n4847), .B(n5198), .Y(n581) );
  INVX1 U938 ( .A(n581), .Y(n582) );
  OR2X2 U939 ( .A(n587), .B(n584), .Y(n583) );
  OR2X2 U940 ( .A(n586), .B(n585), .Y(n584) );
  INVX1 U941 ( .A(n5219), .Y(n585) );
  INVX1 U942 ( .A(n5221), .Y(n586) );
  INVX1 U943 ( .A(n5220), .Y(n587) );
  OR2X2 U944 ( .A(n592), .B(n590), .Y(n588) );
  INVX1 U945 ( .A(n588), .Y(n589) );
  OR2X2 U946 ( .A(n591), .B(n105), .Y(n590) );
  INVX1 U947 ( .A(n5770), .Y(n591) );
  INVX1 U948 ( .A(n5769), .Y(n592) );
  OR2X2 U949 ( .A(n598), .B(n595), .Y(n593) );
  INVX1 U950 ( .A(n593), .Y(n594) );
  OR2X2 U951 ( .A(n596), .B(n597), .Y(n595) );
  INVX1 U952 ( .A(n5137), .Y(n596) );
  INVX1 U953 ( .A(n5138), .Y(n597) );
  INVX1 U954 ( .A(n5139), .Y(n598) );
  OR2X2 U955 ( .A(n603), .B(n600), .Y(n599) );
  OR2X2 U956 ( .A(n601), .B(n602), .Y(n600) );
  INVX1 U957 ( .A(n5164), .Y(n601) );
  INVX1 U958 ( .A(n5165), .Y(n602) );
  INVX1 U959 ( .A(n5166), .Y(n603) );
  OR2X2 U960 ( .A(n607), .B(n605), .Y(n604) );
  OR2X2 U961 ( .A(n816), .B(n606), .Y(n605) );
  INVX1 U962 ( .A(n5196), .Y(n606) );
  INVX1 U963 ( .A(n5197), .Y(n607) );
  OR2X2 U964 ( .A(n612), .B(n609), .Y(n608) );
  OR2X2 U965 ( .A(n611), .B(n610), .Y(n609) );
  INVX1 U966 ( .A(n5229), .Y(n610) );
  INVX1 U967 ( .A(n770), .Y(n611) );
  INVX1 U968 ( .A(n5230), .Y(n612) );
  OR2X2 U969 ( .A(n617), .B(n615), .Y(n613) );
  INVX1 U970 ( .A(n613), .Y(n614) );
  OR2X2 U971 ( .A(n3888), .B(n616), .Y(n615) );
  INVX1 U972 ( .A(n5239), .Y(n616) );
  INVX1 U973 ( .A(n5240), .Y(n617) );
  OR2X2 U974 ( .A(n621), .B(n619), .Y(n618) );
  OR2X2 U975 ( .A(n620), .B(n557), .Y(n619) );
  INVX1 U976 ( .A(n5248), .Y(n620) );
  INVX1 U977 ( .A(n5249), .Y(n621) );
  OR2X2 U978 ( .A(n626), .B(n623), .Y(n622) );
  OR2X2 U979 ( .A(n625), .B(n624), .Y(n623) );
  INVX1 U980 ( .A(n5260), .Y(n624) );
  INVX1 U981 ( .A(n5261), .Y(n625) );
  INVX1 U982 ( .A(n5262), .Y(n626) );
  OR2X2 U983 ( .A(n631), .B(n628), .Y(n627) );
  OR2X2 U984 ( .A(n629), .B(n630), .Y(n628) );
  INVX1 U985 ( .A(n5270), .Y(n629) );
  INVX1 U986 ( .A(n5271), .Y(n630) );
  INVX1 U987 ( .A(n5272), .Y(n631) );
  OR2X2 U988 ( .A(n636), .B(n634), .Y(n632) );
  INVX1 U989 ( .A(n632), .Y(n633) );
  OR2X2 U990 ( .A(n3889), .B(n635), .Y(n634) );
  INVX1 U991 ( .A(n5298), .Y(n635) );
  INVX1 U992 ( .A(n5299), .Y(n636) );
  OR2X2 U993 ( .A(n641), .B(n638), .Y(n637) );
  OR2X2 U994 ( .A(n640), .B(n639), .Y(n638) );
  INVX1 U995 ( .A(n5331), .Y(n639) );
  INVX1 U996 ( .A(n5332), .Y(n640) );
  INVX1 U997 ( .A(n5333), .Y(n641) );
  OR2X2 U998 ( .A(n646), .B(n643), .Y(n642) );
  OR2X2 U999 ( .A(n644), .B(n645), .Y(n643) );
  INVX1 U1000 ( .A(n5395), .Y(n644) );
  INVX1 U1001 ( .A(n5396), .Y(n645) );
  INVX1 U1002 ( .A(n5397), .Y(n646) );
  OR2X2 U1003 ( .A(n649), .B(n650), .Y(n648) );
  INVX1 U1004 ( .A(n5408), .Y(n649) );
  INVX1 U1005 ( .A(n5409), .Y(n650) );
  INVX1 U1006 ( .A(n5410), .Y(n651) );
  OR2X2 U1007 ( .A(n656), .B(n653), .Y(n652) );
  OR2X2 U1008 ( .A(n654), .B(n655), .Y(n653) );
  INVX1 U1009 ( .A(n5419), .Y(n654) );
  INVX1 U1010 ( .A(n5420), .Y(n655) );
  INVX1 U1011 ( .A(n5421), .Y(n656) );
  OR2X2 U1012 ( .A(n157), .B(n659), .Y(n657) );
  INVX1 U1013 ( .A(n657), .Y(n658) );
  OR2X2 U1014 ( .A(n158), .B(n72), .Y(n659) );
  OR2X2 U1015 ( .A(n664), .B(n661), .Y(n660) );
  OR2X2 U1016 ( .A(n662), .B(n663), .Y(n661) );
  INVX1 U1017 ( .A(n5479), .Y(n662) );
  INVX1 U1018 ( .A(n5480), .Y(n663) );
  INVX1 U1019 ( .A(n5481), .Y(n664) );
  OR2X2 U1020 ( .A(n669), .B(n666), .Y(n665) );
  OR2X2 U1021 ( .A(n667), .B(n668), .Y(n666) );
  INVX1 U1022 ( .A(n5502), .Y(n667) );
  INVX1 U1023 ( .A(n5503), .Y(n668) );
  INVX1 U1024 ( .A(n5504), .Y(n669) );
  OR2X2 U1025 ( .A(n159), .B(n672), .Y(n670) );
  INVX1 U1026 ( .A(n670), .Y(n671) );
  OR2X2 U1027 ( .A(n76), .B(n4123), .Y(n672) );
  OR2X2 U1028 ( .A(n677), .B(n675), .Y(n673) );
  INVX1 U1029 ( .A(n673), .Y(n674) );
  OR2X2 U1030 ( .A(n4066), .B(n676), .Y(n675) );
  INVX1 U1031 ( .A(n5530), .Y(n676) );
  INVX1 U1032 ( .A(n5529), .Y(n677) );
  OR2X2 U1033 ( .A(n682), .B(n679), .Y(n678) );
  OR2X2 U1034 ( .A(n680), .B(n681), .Y(n679) );
  INVX1 U1035 ( .A(n5562), .Y(n680) );
  INVX1 U1036 ( .A(n5563), .Y(n681) );
  INVX1 U1037 ( .A(n5564), .Y(n682) );
  OR2X2 U1038 ( .A(n687), .B(n684), .Y(n683) );
  OR2X2 U1039 ( .A(n685), .B(n686), .Y(n684) );
  INVX1 U1040 ( .A(n5586), .Y(n685) );
  INVX1 U1041 ( .A(n5587), .Y(n686) );
  INVX1 U1042 ( .A(n5588), .Y(n687) );
  OR2X2 U1043 ( .A(n4124), .B(n690), .Y(n688) );
  INVX1 U1044 ( .A(n688), .Y(n689) );
  OR2X2 U1045 ( .A(n160), .B(n73), .Y(n690) );
  OR2X2 U1046 ( .A(n695), .B(n692), .Y(n691) );
  OR2X2 U1047 ( .A(n693), .B(n694), .Y(n692) );
  INVX1 U1048 ( .A(n5644), .Y(n693) );
  INVX1 U1049 ( .A(n5645), .Y(n694) );
  INVX1 U1050 ( .A(n5646), .Y(n695) );
  OR2X2 U1051 ( .A(n699), .B(n697), .Y(n696) );
  OR2X2 U1052 ( .A(n698), .B(n563), .Y(n697) );
  INVX1 U1053 ( .A(n5668), .Y(n698) );
  INVX1 U1054 ( .A(n5669), .Y(n699) );
  OR2X2 U1055 ( .A(n161), .B(n702), .Y(n700) );
  INVX1 U1056 ( .A(n700), .Y(n701) );
  OR2X2 U1057 ( .A(n77), .B(n4125), .Y(n702) );
  OR2X2 U1058 ( .A(n707), .B(n705), .Y(n703) );
  INVX1 U1059 ( .A(n703), .Y(n704) );
  OR2X2 U1060 ( .A(n4067), .B(n706), .Y(n705) );
  INVX1 U1061 ( .A(n5697), .Y(n706) );
  INVX1 U1062 ( .A(n5698), .Y(n707) );
  OR2X2 U1063 ( .A(n712), .B(n710), .Y(n708) );
  INVX1 U1064 ( .A(n708), .Y(n709) );
  OR2X2 U1065 ( .A(n711), .B(n828), .Y(n710) );
  INVX1 U1066 ( .A(n5721), .Y(n711) );
  INVX1 U1067 ( .A(n5722), .Y(n712) );
  OR2X2 U1068 ( .A(n75), .B(n714), .Y(n713) );
  OR2X2 U1069 ( .A(n163), .B(n162), .Y(n714) );
  OR2X2 U1070 ( .A(n787), .B(n717), .Y(n715) );
  INVX1 U1071 ( .A(n715), .Y(n716) );
  OR2X2 U1072 ( .A(n718), .B(n719), .Y(n717) );
  INVX1 U1073 ( .A(n5780), .Y(n718) );
  INVX1 U1074 ( .A(n5781), .Y(n719) );
  OR2X2 U1075 ( .A(n1058), .B(n721), .Y(n720) );
  OR2X2 U1076 ( .A(n1056), .B(n1057), .Y(n721) );
  OR2X2 U1077 ( .A(n1246), .B(n723), .Y(n722) );
  OR2X2 U1078 ( .A(n3887), .B(n1245), .Y(n723) );
  OR2X2 U1079 ( .A(n1250), .B(n725), .Y(n724) );
  OR2X2 U1080 ( .A(n3780), .B(n569), .Y(n725) );
  OR2X2 U1081 ( .A(n1252), .B(n727), .Y(n726) );
  OR2X2 U1082 ( .A(n766), .B(n1251), .Y(n727) );
  OR2X2 U1083 ( .A(n1255), .B(n729), .Y(n728) );
  OR2X2 U1084 ( .A(n4122), .B(n1254), .Y(n729) );
  OR2X2 U1085 ( .A(n1256), .B(n62), .Y(n730) );
  OR2X2 U1086 ( .A(n1806), .B(n732), .Y(n731) );
  OR2X2 U1087 ( .A(n1804), .B(n1805), .Y(n732) );
  OR2X2 U1088 ( .A(n2335), .B(n734), .Y(n733) );
  OR2X2 U1089 ( .A(n2333), .B(n2334), .Y(n734) );
  OR2X2 U1090 ( .A(n2338), .B(n736), .Y(n735) );
  OR2X2 U1091 ( .A(n2336), .B(n2337), .Y(n736) );
  OR2X2 U1092 ( .A(n2340), .B(n738), .Y(n737) );
  OR2X2 U1093 ( .A(n2339), .B(n109), .Y(n738) );
  OR2X2 U1094 ( .A(n2343), .B(n740), .Y(n739) );
  OR2X2 U1095 ( .A(n2341), .B(n2342), .Y(n740) );
  OR2X2 U1096 ( .A(n2346), .B(n742), .Y(n741) );
  OR2X2 U1097 ( .A(n2345), .B(n2344), .Y(n742) );
  OR2X2 U1098 ( .A(n3558), .B(n744), .Y(n743) );
  OR2X2 U1099 ( .A(n74), .B(n3557), .Y(n744) );
  OR2X2 U1100 ( .A(n746), .B(n129), .Y(n745) );
  OR2X2 U1101 ( .A(n4867), .B(n3844), .Y(n746) );
  AND2X2 U1102 ( .A(n5167), .B(n146), .Y(n747) );
  OR2X2 U1103 ( .A(n126), .B(n4915), .Y(n749) );
  OR2X2 U1104 ( .A(n568), .B(n5126), .Y(n750) );
  AND2X2 U1105 ( .A(n1214), .B(n1200), .Y(n751) );
  AND2X2 U1106 ( .A(n1218), .B(n1202), .Y(n752) );
  AND2X2 U1107 ( .A(n1222), .B(n1204), .Y(n753) );
  AND2X2 U1108 ( .A(n1226), .B(n1206), .Y(n754) );
  AND2X2 U1109 ( .A(n1208), .B(n1230), .Y(n755) );
  AND2X2 U1110 ( .A(n1234), .B(n1210), .Y(n756) );
  AND2X2 U1111 ( .A(n1238), .B(n1212), .Y(n757) );
  AND2X2 U1112 ( .A(n5745), .B(n5744), .Y(n758) );
  OR2X2 U1113 ( .A(n4914), .B(n760), .Y(n759) );
  OR2X2 U1114 ( .A(n3952), .B(n3953), .Y(n760) );
  OR2X2 U1115 ( .A(n4684), .B(n762), .Y(n761) );
  OR2X2 U1116 ( .A(rst), .B(n4683), .Y(n762) );
  AND2X2 U1117 ( .A(n716), .B(n589), .Y(n763) );
  AND2X2 U1118 ( .A(n4709), .B(n4710), .Y(n765) );
  INVX1 U1119 ( .A(n765), .Y(n766) );
  OR2X2 U1120 ( .A(n4711), .B(n4695), .Y(n767) );
  INVX1 U1121 ( .A(n767), .Y(\data_out<11> ) );
  AND2X2 U1122 ( .A(n4728), .B(n4729), .Y(n769) );
  AND2X2 U1123 ( .A(n4795), .B(n4794), .Y(n770) );
  OR2X2 U1124 ( .A(n3876), .B(n4735), .Y(n771) );
  AND2X2 U1125 ( .A(n4755), .B(n4756), .Y(n772) );
  OR2X2 U1126 ( .A(n4730), .B(n4696), .Y(n773) );
  INVX1 U1127 ( .A(n773), .Y(\data_out<14> ) );
  AND2X2 U1128 ( .A(n52), .B(n6410), .Y(n775) );
  OR2X2 U1129 ( .A(n3676), .B(n4735), .Y(n776) );
  INVX1 U1130 ( .A(n776), .Y(n777) );
  OR2X2 U1131 ( .A(n4740), .B(n4696), .Y(n778) );
  INVX1 U1132 ( .A(n778), .Y(\data_out<15> ) );
  OR2X2 U1133 ( .A(n4741), .B(n4695), .Y(n780) );
  INVX1 U1134 ( .A(n780), .Y(\data_out<9> ) );
  OR2X2 U1135 ( .A(n3875), .B(n6352), .Y(n782) );
  INVX1 U1136 ( .A(n782), .Y(n783) );
  OR2X2 U1137 ( .A(n4744), .B(n4694), .Y(n784) );
  INVX1 U1138 ( .A(n784), .Y(\data_out<13> ) );
  AND2X2 U1139 ( .A(n4746), .B(n4747), .Y(n786) );
  INVX1 U1140 ( .A(n786), .Y(n787) );
  OR2X2 U1141 ( .A(n4748), .B(n4695), .Y(n788) );
  INVX1 U1142 ( .A(n788), .Y(\data_out<10> ) );
  AND2X2 U1143 ( .A(n4761), .B(n4762), .Y(n790) );
  AND2X2 U1144 ( .A(n4771), .B(n4772), .Y(n791) );
  OR2X2 U1145 ( .A(n6357), .B(n6404), .Y(n792) );
  AND2X2 U1146 ( .A(n4780), .B(n4781), .Y(n793) );
  AND2X2 U1147 ( .A(n633), .B(n4786), .Y(n795) );
  OR2X2 U1148 ( .A(n4801), .B(n4735), .Y(n796) );
  OR2X2 U1149 ( .A(n1), .B(n4963), .Y(n797) );
  OR2X2 U1150 ( .A(n4819), .B(n125), .Y(n798) );
  OR2X2 U1151 ( .A(n5037), .B(n5008), .Y(n799) );
  OR2X2 U1152 ( .A(n5017), .B(n799), .Y(n800) );
  AND2X2 U1153 ( .A(n3949), .B(n1198), .Y(n801) );
  AND2X2 U1154 ( .A(n5709), .B(n5708), .Y(n802) );
  OR2X2 U1155 ( .A(n61), .B(n6352), .Y(n803) );
  OR2X2 U1156 ( .A(n1242), .B(n4836), .Y(n805) );
  OR2X2 U1157 ( .A(n61), .B(n4909), .Y(n806) );
  OR2X2 U1158 ( .A(n5019), .B(n4885), .Y(n807) );
  OR2X2 U1159 ( .A(\addr<11> ), .B(\addr<13> ), .Y(n808) );
  OR2X2 U1160 ( .A(n759), .B(n1260), .Y(n809) );
  INVX1 U1161 ( .A(n809), .Y(n810) );
  OR2X2 U1162 ( .A(n1244), .B(n3955), .Y(n811) );
  INVX1 U1163 ( .A(n811), .Y(n812) );
  AND2X2 U1164 ( .A(n4996), .B(n5002), .Y(n813) );
  AND2X2 U1165 ( .A(n562), .B(n147), .Y(n814) );
  INVX1 U1166 ( .A(n814), .Y(n815) );
  OR2X2 U1167 ( .A(n5194), .B(n5195), .Y(n816) );
  OR2X2 U1168 ( .A(n4953), .B(n5198), .Y(n817) );
  INVX1 U1169 ( .A(n817), .Y(n818) );
  AND2X2 U1170 ( .A(n122), .B(n80), .Y(n819) );
  OR2X2 U1171 ( .A(n5424), .B(n4907), .Y(n820) );
  INVX1 U1172 ( .A(n820), .Y(n821) );
  OR2X2 U1173 ( .A(n5507), .B(n4902), .Y(n822) );
  INVX1 U1174 ( .A(n822), .Y(n823) );
  OR2X2 U1175 ( .A(n5591), .B(n4908), .Y(n824) );
  INVX1 U1176 ( .A(n824), .Y(n825) );
  OR2X2 U1177 ( .A(n5672), .B(n4907), .Y(n826) );
  INVX1 U1178 ( .A(n826), .Y(n827) );
  OR2X2 U1179 ( .A(n5715), .B(n5716), .Y(n828) );
  AND2X2 U1180 ( .A(n5723), .B(n3685), .Y(n829) );
  INVX1 U1181 ( .A(n829), .Y(n830) );
  AND2X2 U1182 ( .A(n6287), .B(n4974), .Y(n831) );
  AND2X2 U1183 ( .A(n5072), .B(n6292), .Y(n832) );
  INVX1 U1184 ( .A(n832), .Y(n833) );
  AND2X2 U1185 ( .A(n5078), .B(n6292), .Y(n834) );
  INVX1 U1186 ( .A(n834), .Y(n835) );
  AND2X2 U1187 ( .A(n5085), .B(n6292), .Y(n836) );
  INVX1 U1188 ( .A(n836), .Y(n837) );
  AND2X2 U1189 ( .A(n5090), .B(n6292), .Y(n838) );
  INVX1 U1190 ( .A(n838), .Y(n839) );
  AND2X2 U1191 ( .A(n5095), .B(n6292), .Y(n840) );
  INVX1 U1192 ( .A(n840), .Y(n841) );
  AND2X2 U1193 ( .A(n5099), .B(n6292), .Y(n842) );
  INVX1 U1194 ( .A(n842), .Y(n843) );
  AND2X2 U1195 ( .A(n5104), .B(n6292), .Y(n844) );
  INVX1 U1196 ( .A(n844), .Y(n845) );
  AND2X2 U1197 ( .A(n5107), .B(n6292), .Y(n846) );
  INVX1 U1198 ( .A(n846), .Y(n847) );
  AND2X2 U1199 ( .A(n1692), .B(n5047), .Y(n848) );
  INVX1 U1200 ( .A(n848), .Y(n849) );
  AND2X2 U1201 ( .A(n1692), .B(n5061), .Y(n850) );
  INVX1 U1202 ( .A(n850), .Y(n851) );
  AND2X2 U1203 ( .A(n5039), .B(n1694), .Y(n852) );
  INVX1 U1204 ( .A(n852), .Y(n853) );
  AND2X2 U1205 ( .A(n5072), .B(n1695), .Y(n854) );
  INVX1 U1206 ( .A(n854), .Y(n855) );
  AND2X2 U1207 ( .A(n5045), .B(n1694), .Y(n856) );
  INVX1 U1208 ( .A(n856), .Y(n857) );
  AND2X2 U1209 ( .A(n5078), .B(n1695), .Y(n858) );
  INVX1 U1210 ( .A(n858), .Y(n859) );
  AND2X2 U1211 ( .A(n5048), .B(n1694), .Y(n860) );
  INVX1 U1212 ( .A(n860), .Y(n861) );
  AND2X2 U1213 ( .A(n5084), .B(n1695), .Y(n862) );
  INVX1 U1214 ( .A(n862), .Y(n863) );
  AND2X2 U1215 ( .A(n5052), .B(n1694), .Y(n864) );
  INVX1 U1216 ( .A(n864), .Y(n865) );
  AND2X2 U1217 ( .A(n5089), .B(n1695), .Y(n866) );
  INVX1 U1218 ( .A(n866), .Y(n867) );
  AND2X2 U1219 ( .A(n5057), .B(n1694), .Y(n868) );
  INVX1 U1220 ( .A(n868), .Y(n869) );
  AND2X2 U1221 ( .A(n5095), .B(n1695), .Y(n870) );
  INVX1 U1222 ( .A(n870), .Y(n871) );
  AND2X2 U1223 ( .A(n5061), .B(n1694), .Y(n872) );
  INVX1 U1224 ( .A(n872), .Y(n873) );
  AND2X2 U1225 ( .A(n5099), .B(n1695), .Y(n874) );
  INVX1 U1226 ( .A(n874), .Y(n875) );
  AND2X2 U1227 ( .A(n5066), .B(n1694), .Y(n876) );
  AND2X2 U1228 ( .A(n5103), .B(n1695), .Y(n877) );
  INVX1 U1229 ( .A(n877), .Y(n878) );
  AND2X2 U1230 ( .A(n5070), .B(n1694), .Y(n879) );
  INVX1 U1231 ( .A(n879), .Y(n880) );
  AND2X2 U1232 ( .A(n5108), .B(n1695), .Y(n881) );
  INVX1 U1233 ( .A(n881), .Y(n882) );
  AND2X2 U1234 ( .A(n5072), .B(n1699), .Y(n883) );
  INVX1 U1235 ( .A(n883), .Y(n884) );
  AND2X2 U1236 ( .A(n5078), .B(n1699), .Y(n885) );
  INVX1 U1237 ( .A(n885), .Y(n886) );
  AND2X2 U1238 ( .A(n5084), .B(n1699), .Y(n887) );
  INVX1 U1239 ( .A(n887), .Y(n888) );
  AND2X2 U1240 ( .A(n5089), .B(n1699), .Y(n889) );
  INVX1 U1241 ( .A(n889), .Y(n890) );
  AND2X2 U1242 ( .A(n5095), .B(n1699), .Y(n891) );
  INVX1 U1243 ( .A(n891), .Y(n892) );
  AND2X2 U1244 ( .A(n5099), .B(n1699), .Y(n893) );
  INVX1 U1245 ( .A(n893), .Y(n894) );
  AND2X2 U1246 ( .A(n5103), .B(n1699), .Y(n895) );
  INVX1 U1247 ( .A(n895), .Y(n896) );
  AND2X2 U1248 ( .A(n5039), .B(n1700), .Y(n897) );
  INVX1 U1249 ( .A(n897), .Y(n898) );
  AND2X2 U1250 ( .A(n5045), .B(n1700), .Y(n899) );
  INVX1 U1251 ( .A(n899), .Y(n900) );
  AND2X2 U1252 ( .A(n5048), .B(n1700), .Y(n901) );
  INVX1 U1253 ( .A(n901), .Y(n902) );
  AND2X2 U1254 ( .A(n5052), .B(n1700), .Y(n903) );
  INVX1 U1255 ( .A(n903), .Y(n904) );
  AND2X2 U1256 ( .A(n5057), .B(n1700), .Y(n905) );
  INVX1 U1257 ( .A(n905), .Y(n906) );
  AND2X2 U1258 ( .A(n5061), .B(n1700), .Y(n907) );
  INVX1 U1259 ( .A(n907), .Y(n908) );
  AND2X2 U1260 ( .A(n5066), .B(n1700), .Y(n909) );
  AND2X2 U1261 ( .A(n5070), .B(n1700), .Y(n910) );
  INVX1 U1262 ( .A(n910), .Y(n911) );
  AND2X2 U1263 ( .A(n5047), .B(n1706), .Y(n912) );
  INVX1 U1264 ( .A(n912), .Y(n913) );
  AND2X2 U1265 ( .A(n5057), .B(n1706), .Y(n914) );
  INVX1 U1266 ( .A(n914), .Y(n915) );
  AND2X2 U1267 ( .A(n5061), .B(n1706), .Y(n916) );
  INVX1 U1268 ( .A(n916), .Y(n917) );
  AND2X2 U1269 ( .A(n5066), .B(n1706), .Y(n918) );
  INVX1 U1270 ( .A(n918), .Y(n919) );
  AND2X2 U1271 ( .A(n5039), .B(n1714), .Y(n920) );
  INVX1 U1272 ( .A(n920), .Y(n921) );
  AND2X2 U1273 ( .A(n5072), .B(n1715), .Y(n922) );
  INVX1 U1274 ( .A(n922), .Y(n923) );
  AND2X2 U1275 ( .A(n5044), .B(n1714), .Y(n924) );
  INVX1 U1276 ( .A(n924), .Y(n925) );
  AND2X2 U1277 ( .A(n5077), .B(n1715), .Y(n926) );
  INVX1 U1278 ( .A(n926), .Y(n927) );
  AND2X2 U1279 ( .A(\data_in<2> ), .B(n1714), .Y(n928) );
  INVX1 U1280 ( .A(n928), .Y(n929) );
  AND2X2 U1281 ( .A(n5082), .B(n1715), .Y(n930) );
  INVX1 U1282 ( .A(n930), .Y(n931) );
  AND2X2 U1283 ( .A(n5052), .B(n1714), .Y(n932) );
  INVX1 U1284 ( .A(n932), .Y(n933) );
  AND2X2 U1285 ( .A(n5089), .B(n1715), .Y(n934) );
  INVX1 U1286 ( .A(n934), .Y(n935) );
  AND2X2 U1287 ( .A(n5057), .B(n1714), .Y(n936) );
  INVX1 U1288 ( .A(n936), .Y(n937) );
  AND2X2 U1289 ( .A(n5094), .B(n1715), .Y(n938) );
  INVX1 U1290 ( .A(n938), .Y(n939) );
  AND2X2 U1291 ( .A(n5061), .B(n1714), .Y(n940) );
  INVX1 U1292 ( .A(n940), .Y(n941) );
  AND2X2 U1293 ( .A(n5098), .B(n1715), .Y(n942) );
  INVX1 U1294 ( .A(n942), .Y(n943) );
  AND2X2 U1295 ( .A(n5066), .B(n1714), .Y(n944) );
  INVX1 U1296 ( .A(n944), .Y(n945) );
  AND2X2 U1297 ( .A(n5102), .B(n1715), .Y(n946) );
  INVX1 U1298 ( .A(n946), .Y(n947) );
  AND2X2 U1299 ( .A(n5070), .B(n1714), .Y(n948) );
  INVX1 U1300 ( .A(n948), .Y(n949) );
  AND2X2 U1301 ( .A(n5108), .B(n1715), .Y(n950) );
  INVX1 U1302 ( .A(n950), .Y(n951) );
  AND2X2 U1303 ( .A(n147), .B(n3), .Y(n952) );
  AND2X2 U1304 ( .A(n148), .B(n4967), .Y(n953) );
  AND2X2 U1305 ( .A(n4818), .B(n3), .Y(n954) );
  AND2X2 U1306 ( .A(n4818), .B(n4967), .Y(n955) );
  AND2X2 U1307 ( .A(n5049), .B(n1746), .Y(n956) );
  INVX1 U1308 ( .A(n956), .Y(n957) );
  AND2X2 U1309 ( .A(n5055), .B(n1746), .Y(n958) );
  INVX1 U1310 ( .A(n958), .Y(n959) );
  AND2X2 U1311 ( .A(n5060), .B(n1746), .Y(n960) );
  INVX1 U1312 ( .A(n960), .Y(n961) );
  AND2X2 U1313 ( .A(n5064), .B(n1746), .Y(n962) );
  INVX1 U1314 ( .A(n962), .Y(n963) );
  AND2X2 U1315 ( .A(n5073), .B(n6356), .Y(n964) );
  INVX1 U1316 ( .A(n964), .Y(n965) );
  AND2X2 U1317 ( .A(n5078), .B(n6356), .Y(n966) );
  INVX1 U1318 ( .A(n966), .Y(n967) );
  AND2X2 U1319 ( .A(n5082), .B(n6356), .Y(n968) );
  INVX1 U1320 ( .A(n968), .Y(n969) );
  AND2X2 U1321 ( .A(n5087), .B(n6356), .Y(n970) );
  INVX1 U1322 ( .A(n970), .Y(n971) );
  AND2X2 U1323 ( .A(n5095), .B(n6356), .Y(n972) );
  INVX1 U1324 ( .A(n972), .Y(n973) );
  AND2X2 U1325 ( .A(n5099), .B(n6356), .Y(n974) );
  INVX1 U1326 ( .A(n974), .Y(n975) );
  AND2X2 U1327 ( .A(n5103), .B(n6356), .Y(n976) );
  INVX1 U1328 ( .A(n976), .Y(n977) );
  AND2X2 U1329 ( .A(n5107), .B(n6356), .Y(n978) );
  INVX1 U1330 ( .A(n978), .Y(n979) );
  AND2X2 U1331 ( .A(n5075), .B(n3716), .Y(n980) );
  INVX1 U1332 ( .A(n980), .Y(n981) );
  AND2X2 U1333 ( .A(n5079), .B(n3716), .Y(n982) );
  INVX1 U1334 ( .A(n982), .Y(n983) );
  AND2X2 U1335 ( .A(n5083), .B(n3716), .Y(n984) );
  INVX1 U1336 ( .A(n984), .Y(n985) );
  AND2X2 U1337 ( .A(n5088), .B(n3716), .Y(n986) );
  INVX1 U1338 ( .A(n986), .Y(n987) );
  AND2X2 U1339 ( .A(n5095), .B(n3716), .Y(n988) );
  INVX1 U1340 ( .A(n988), .Y(n989) );
  AND2X2 U1341 ( .A(n5100), .B(n3716), .Y(n990) );
  INVX1 U1342 ( .A(n990), .Y(n991) );
  AND2X2 U1343 ( .A(n5103), .B(n3716), .Y(n992) );
  INVX1 U1344 ( .A(n992), .Y(n993) );
  AND2X2 U1345 ( .A(n5109), .B(n3716), .Y(n994) );
  INVX1 U1346 ( .A(n994), .Y(n995) );
  AND2X2 U1347 ( .A(n5072), .B(n1773), .Y(n996) );
  INVX1 U1348 ( .A(n996), .Y(n997) );
  AND2X2 U1349 ( .A(n5078), .B(n1773), .Y(n998) );
  INVX1 U1350 ( .A(n998), .Y(n999) );
  AND2X2 U1351 ( .A(n5083), .B(n1773), .Y(n1000) );
  INVX1 U1352 ( .A(n1000), .Y(n1001) );
  AND2X2 U1353 ( .A(n5088), .B(n1773), .Y(n1002) );
  INVX1 U1354 ( .A(n1002), .Y(n1003) );
  AND2X2 U1355 ( .A(n5056), .B(n1772), .Y(n1004) );
  INVX1 U1356 ( .A(n1004), .Y(n1005) );
  AND2X2 U1357 ( .A(n5095), .B(n1773), .Y(n1006) );
  INVX1 U1358 ( .A(n1006), .Y(n1007) );
  AND2X2 U1359 ( .A(n5060), .B(n1772), .Y(n1008) );
  AND2X2 U1360 ( .A(n5099), .B(n1773), .Y(n1009) );
  INVX1 U1361 ( .A(n1009), .Y(n1010) );
  AND2X2 U1362 ( .A(n5065), .B(n1772), .Y(n1011) );
  INVX1 U1363 ( .A(n1011), .Y(n1012) );
  AND2X2 U1364 ( .A(n5103), .B(n1773), .Y(n1013) );
  INVX1 U1365 ( .A(n1013), .Y(n1014) );
  AND2X2 U1366 ( .A(n5108), .B(n1773), .Y(n1015) );
  INVX1 U1367 ( .A(n1015), .Y(n1016) );
  AND2X2 U1368 ( .A(n5074), .B(n3877), .Y(n1017) );
  AND2X2 U1369 ( .A(n5078), .B(n3878), .Y(n1018) );
  AND2X2 U1370 ( .A(n5083), .B(n3877), .Y(n1019) );
  INVX1 U1371 ( .A(n1019), .Y(n1020) );
  AND2X2 U1372 ( .A(n5088), .B(n3878), .Y(n1021) );
  INVX1 U1373 ( .A(n1021), .Y(n1022) );
  AND2X2 U1374 ( .A(n5095), .B(n3877), .Y(n1023) );
  INVX1 U1375 ( .A(n1023), .Y(n1024) );
  AND2X2 U1376 ( .A(n5100), .B(n3878), .Y(n1025) );
  INVX1 U1377 ( .A(n1025), .Y(n1026) );
  AND2X2 U1378 ( .A(n5103), .B(n3877), .Y(n1027) );
  INVX1 U1379 ( .A(n1027), .Y(n1028) );
  AND2X2 U1380 ( .A(n5109), .B(n3878), .Y(n1029) );
  INVX1 U1381 ( .A(n1029), .Y(n1030) );
  AND2X2 U1382 ( .A(n4969), .B(n4967), .Y(n1031) );
  AND2X2 U1383 ( .A(n5038), .B(n1803), .Y(n1032) );
  INVX1 U1384 ( .A(n1032), .Y(n1033) );
  AND2X2 U1385 ( .A(n5041), .B(n1803), .Y(n1034) );
  INVX1 U1386 ( .A(n1034), .Y(n1035) );
  AND2X2 U1387 ( .A(n5047), .B(n1803), .Y(n1036) );
  INVX1 U1388 ( .A(n1036), .Y(n1037) );
  AND2X2 U1389 ( .A(n5051), .B(n1803), .Y(n1038) );
  INVX1 U1390 ( .A(n1038), .Y(n1039) );
  AND2X2 U1391 ( .A(n5055), .B(n1803), .Y(n1040) );
  INVX1 U1392 ( .A(n1040), .Y(n1041) );
  AND2X2 U1393 ( .A(n1803), .B(n5060), .Y(n1042) );
  INVX1 U1394 ( .A(n1042), .Y(n1043) );
  AND2X2 U1395 ( .A(n5064), .B(n1803), .Y(n1044) );
  INVX1 U1396 ( .A(n1044), .Y(n1045) );
  AND2X2 U1397 ( .A(n5069), .B(n1803), .Y(n1046) );
  INVX1 U1398 ( .A(n1046), .Y(n1047) );
  OR2X2 U1399 ( .A(\addr<12> ), .B(\addr<10> ), .Y(n1048) );
  INVX1 U1400 ( .A(n1048), .Y(n1049) );
  OR2X2 U1401 ( .A(n5008), .B(n5033), .Y(n1050) );
  INVX1 U1402 ( .A(n1050), .Y(n1051) );
  AND2X2 U1403 ( .A(n4830), .B(n4622), .Y(n1052) );
  INVX1 U1404 ( .A(n1052), .Y(n1053) );
  AND2X2 U1405 ( .A(n4829), .B(n4643), .Y(n1054) );
  INVX1 U1406 ( .A(n1054), .Y(n1055) );
  INVX1 U1407 ( .A(n5735), .Y(n1056) );
  INVX1 U1408 ( .A(n5736), .Y(n1057) );
  INVX1 U1409 ( .A(n5737), .Y(n1058) );
  AND2X2 U1410 ( .A(n758), .B(n5743), .Y(n1059) );
  INVX1 U1411 ( .A(n1059), .Y(n1060) );
  OR2X2 U1412 ( .A(\addr<9> ), .B(\addr<6> ), .Y(n1061) );
  INVX1 U1413 ( .A(n1061), .Y(n1062) );
  AND2X2 U1414 ( .A(n6302), .B(n3652), .Y(n1063) );
  INVX1 U1415 ( .A(n1063), .Y(n1064) );
  AND2X2 U1416 ( .A(n104), .B(n566), .Y(n1065) );
  INVX1 U1417 ( .A(n1065), .Y(n1066) );
  AND2X2 U1418 ( .A(n4719), .B(n4653), .Y(n1067) );
  INVX1 U1419 ( .A(n1067), .Y(n1068) );
  AND2X2 U1420 ( .A(n6313), .B(n4631), .Y(n1069) );
  INVX1 U1421 ( .A(n1069), .Y(n1070) );
  AND2X2 U1422 ( .A(n3669), .B(n4630), .Y(n1071) );
  INVX1 U1423 ( .A(n1071), .Y(n1072) );
  AND2X2 U1424 ( .A(n6314), .B(n3669), .Y(n1073) );
  INVX1 U1425 ( .A(n1073), .Y(n1074) );
  AND2X2 U1426 ( .A(n93), .B(n4812), .Y(n1075) );
  INVX1 U1427 ( .A(n1075), .Y(n1076) );
  AND2X2 U1428 ( .A(n96), .B(n35), .Y(n1077) );
  INVX1 U1429 ( .A(n1077), .Y(n1078) );
  AND2X2 U1430 ( .A(n6330), .B(n3860), .Y(n1079) );
  INVX1 U1431 ( .A(n1079), .Y(n1080) );
  AND2X2 U1432 ( .A(n6330), .B(n4633), .Y(n1081) );
  INVX1 U1433 ( .A(n1081), .Y(n1082) );
  AND2X2 U1434 ( .A(n1684), .B(n4634), .Y(n1083) );
  INVX1 U1435 ( .A(n1083), .Y(n1084) );
  AND2X2 U1436 ( .A(n1684), .B(n3677), .Y(n1085) );
  INVX1 U1437 ( .A(n1085), .Y(n1086) );
  AND2X2 U1438 ( .A(n4649), .B(n3677), .Y(n1087) );
  INVX1 U1439 ( .A(n1087), .Y(n1088) );
  AND2X2 U1440 ( .A(n88), .B(n4649), .Y(n1089) );
  INVX1 U1441 ( .A(n1089), .Y(n1090) );
  AND2X2 U1442 ( .A(n6342), .B(n16), .Y(n1091) );
  INVX1 U1443 ( .A(n1091), .Y(n1092) );
  AND2X2 U1444 ( .A(n6342), .B(n4636), .Y(n1093) );
  INVX1 U1445 ( .A(n1093), .Y(n1094) );
  AND2X2 U1446 ( .A(n6344), .B(n4637), .Y(n1095) );
  INVX1 U1447 ( .A(n1095), .Y(n1096) );
  AND2X2 U1448 ( .A(n6344), .B(n6345), .Y(n1097) );
  INVX1 U1449 ( .A(n1097), .Y(n1098) );
  AND2X2 U1450 ( .A(n4918), .B(n4664), .Y(n1099) );
  INVX1 U1451 ( .A(n1099), .Y(n1100) );
  AND2X2 U1452 ( .A(n3575), .B(n3850), .Y(n1101) );
  INVX1 U1453 ( .A(n1101), .Y(n1102) );
  AND2X2 U1454 ( .A(n3575), .B(n6370), .Y(n1103) );
  INVX1 U1455 ( .A(n1103), .Y(n1104) );
  AND2X2 U1456 ( .A(n3560), .B(n4751), .Y(n1105) );
  INVX1 U1457 ( .A(n1105), .Y(n1106) );
  AND2X2 U1458 ( .A(n6378), .B(n3846), .Y(n1107) );
  INVX1 U1459 ( .A(n1107), .Y(n1108) );
  AND2X2 U1460 ( .A(n4639), .B(n6378), .Y(n1109) );
  INVX1 U1461 ( .A(n1109), .Y(n1110) );
  AND2X2 U1462 ( .A(n4823), .B(n4640), .Y(n1111) );
  INVX1 U1463 ( .A(n1111), .Y(n1112) );
  AND2X2 U1464 ( .A(n4823), .B(n6388), .Y(n1113) );
  INVX1 U1465 ( .A(n1113), .Y(n1114) );
  AND2X2 U1466 ( .A(n3673), .B(n4660), .Y(n1115) );
  INVX1 U1467 ( .A(n1115), .Y(n1116) );
  AND2X2 U1468 ( .A(n4828), .B(n4644), .Y(n1117) );
  INVX1 U1469 ( .A(n1117), .Y(n1118) );
  AND2X2 U1470 ( .A(n4828), .B(n4821), .Y(n1119) );
  INVX1 U1471 ( .A(n1119), .Y(n1120) );
  AND2X2 U1472 ( .A(n4678), .B(n3578), .Y(n1121) );
  INVX1 U1473 ( .A(n1121), .Y(n1122) );
  AND2X2 U1474 ( .A(n4870), .B(n37), .Y(n1123) );
  INVX1 U1475 ( .A(n1123), .Y(n1124) );
  AND2X2 U1476 ( .A(n6414), .B(n89), .Y(n1125) );
  INVX1 U1477 ( .A(n1125), .Y(n1126) );
  AND2X2 U1478 ( .A(n6414), .B(n4647), .Y(n1127) );
  INVX1 U1479 ( .A(n1127), .Y(n1128) );
  AND2X2 U1480 ( .A(n4879), .B(n4648), .Y(n1129) );
  INVX1 U1481 ( .A(n1129), .Y(n1130) );
  AND2X2 U1482 ( .A(n5187), .B(n4860), .Y(n1131) );
  INVX1 U1483 ( .A(n1131), .Y(n1132) );
  AND2X2 U1484 ( .A(\mem<44><0> ), .B(n4868), .Y(n1133) );
  INVX1 U1485 ( .A(n1133), .Y(n1134) );
  AND2X2 U1486 ( .A(\mem<53><0> ), .B(n4873), .Y(n1135) );
  INVX1 U1487 ( .A(n1135), .Y(n1136) );
  AND2X2 U1488 ( .A(\mem<54><0> ), .B(n4873), .Y(n1137) );
  INVX1 U1489 ( .A(n1137), .Y(n1138) );
  AND2X2 U1490 ( .A(\mem<44><1> ), .B(n4868), .Y(n1139) );
  INVX1 U1491 ( .A(n1139), .Y(n1140) );
  AND2X2 U1492 ( .A(n4893), .B(n5243), .Y(n1141) );
  INVX1 U1493 ( .A(n1141), .Y(n1142) );
  INVX1 U1494 ( .A(n1143), .Y(n1144) );
  AND2X2 U1495 ( .A(n127), .B(n5265), .Y(n1145) );
  INVX1 U1496 ( .A(n1145), .Y(n1146) );
  AND2X2 U1497 ( .A(n4899), .B(n5302), .Y(n1147) );
  INVX1 U1498 ( .A(n1147), .Y(n1148) );
  AND2X2 U1499 ( .A(n4893), .B(n5315), .Y(n1149) );
  INVX1 U1500 ( .A(n1149), .Y(n1150) );
  INVX1 U1501 ( .A(n1151), .Y(n1152) );
  INVX1 U1502 ( .A(n1153), .Y(n1154) );
  AND2X2 U1503 ( .A(\mem<24><2> ), .B(n3867), .Y(n1155) );
  INVX1 U1504 ( .A(n1155), .Y(n1156) );
  INVX1 U1505 ( .A(n1157), .Y(n1158) );
  INVX1 U1506 ( .A(n1159), .Y(n1160) );
  AND2X2 U1507 ( .A(n4941), .B(n5413), .Y(n1161) );
  INVX1 U1508 ( .A(n1161), .Y(n1162) );
  AND2X2 U1509 ( .A(\mem<58><3> ), .B(n83), .Y(n1163) );
  INVX1 U1510 ( .A(n1163), .Y(n1164) );
  INVX1 U1511 ( .A(n1165), .Y(n1166) );
  AND2X2 U1512 ( .A(n4891), .B(n5487), .Y(n1167) );
  INVX1 U1513 ( .A(n1167), .Y(n1168) );
  AND2X2 U1514 ( .A(n4903), .B(n5497), .Y(n1169) );
  INVX1 U1515 ( .A(n1169), .Y(n1170) );
  AND2X2 U1516 ( .A(\mem<58><4> ), .B(n84), .Y(n1171) );
  INVX1 U1517 ( .A(n1171), .Y(n1172) );
  AND2X2 U1518 ( .A(\mem<44><4> ), .B(n4868), .Y(n1173) );
  INVX1 U1519 ( .A(n1173), .Y(n1174) );
  INVX1 U1520 ( .A(n1175), .Y(n1176) );
  INVX1 U1521 ( .A(n1177), .Y(n1178) );
  INVX1 U1522 ( .A(n1179), .Y(n1180) );
  AND2X2 U1523 ( .A(\mem<58><5> ), .B(n83), .Y(n1181) );
  INVX1 U1524 ( .A(n1181), .Y(n1182) );
  AND2X2 U1525 ( .A(\mem<40><5> ), .B(n116), .Y(n1183) );
  INVX1 U1526 ( .A(n1183), .Y(n1184) );
  AND2X2 U1527 ( .A(\mem<44><5> ), .B(n4868), .Y(n1185) );
  INVX1 U1528 ( .A(n1185), .Y(n1186) );
  AND2X2 U1529 ( .A(\mem<52><6> ), .B(n4877), .Y(n1187) );
  INVX1 U1530 ( .A(n1187), .Y(n1188) );
  AND2X2 U1531 ( .A(n4899), .B(n5639), .Y(n1189) );
  INVX1 U1532 ( .A(n1189), .Y(n1190) );
  AND2X2 U1533 ( .A(\mem<58><6> ), .B(n84), .Y(n1191) );
  INVX1 U1534 ( .A(n1191), .Y(n1192) );
  AND2X2 U1535 ( .A(\mem<40><6> ), .B(n116), .Y(n1193) );
  INVX1 U1536 ( .A(n1193), .Y(n1194) );
  AND2X2 U1537 ( .A(\mem<58><7> ), .B(n3864), .Y(n1195) );
  INVX1 U1538 ( .A(n1195), .Y(n1196) );
  AND2X2 U1539 ( .A(n6158), .B(n4841), .Y(n1197) );
  INVX1 U1540 ( .A(n1197), .Y(n1198) );
  AND2X2 U1541 ( .A(n5077), .B(n3714), .Y(n1199) );
  INVX1 U1542 ( .A(n1199), .Y(n1200) );
  AND2X2 U1543 ( .A(\data_in<10> ), .B(n3714), .Y(n1201) );
  INVX1 U1544 ( .A(n1201), .Y(n1202) );
  AND2X2 U1545 ( .A(\data_in<11> ), .B(n3714), .Y(n1203) );
  INVX1 U1546 ( .A(n1203), .Y(n1204) );
  AND2X2 U1547 ( .A(n5094), .B(n3714), .Y(n1205) );
  INVX1 U1548 ( .A(n1205), .Y(n1206) );
  AND2X2 U1549 ( .A(n5098), .B(n3714), .Y(n1207) );
  INVX1 U1550 ( .A(n1207), .Y(n1208) );
  AND2X2 U1551 ( .A(n5102), .B(n3714), .Y(n1209) );
  INVX1 U1552 ( .A(n1209), .Y(n1210) );
  AND2X2 U1553 ( .A(\data_in<15> ), .B(n3714), .Y(n1211) );
  INVX1 U1554 ( .A(n1211), .Y(n1212) );
  AND2X2 U1555 ( .A(n5045), .B(n1713), .Y(n1213) );
  INVX1 U1556 ( .A(n1213), .Y(n1214) );
  AND2X2 U1557 ( .A(\mem<49><1> ), .B(n3592), .Y(n1215) );
  INVX1 U1558 ( .A(n1215), .Y(n1216) );
  AND2X2 U1559 ( .A(\data_in<2> ), .B(n1713), .Y(n1217) );
  INVX1 U1560 ( .A(n1217), .Y(n1218) );
  AND2X2 U1561 ( .A(\mem<49><2> ), .B(n3592), .Y(n1219) );
  INVX1 U1562 ( .A(n1219), .Y(n1220) );
  AND2X2 U1563 ( .A(n5052), .B(n1713), .Y(n1221) );
  INVX1 U1564 ( .A(n1221), .Y(n1222) );
  AND2X2 U1565 ( .A(\mem<49><3> ), .B(n3592), .Y(n1223) );
  INVX1 U1566 ( .A(n1223), .Y(n1224) );
  AND2X2 U1567 ( .A(n5057), .B(n1713), .Y(n1225) );
  INVX1 U1568 ( .A(n1225), .Y(n1226) );
  AND2X2 U1569 ( .A(\mem<49><4> ), .B(n3592), .Y(n1227) );
  INVX1 U1570 ( .A(n1227), .Y(n1228) );
  AND2X2 U1571 ( .A(n5061), .B(n1713), .Y(n1229) );
  INVX1 U1572 ( .A(n1229), .Y(n1230) );
  AND2X2 U1573 ( .A(\mem<49><5> ), .B(n3592), .Y(n1231) );
  INVX1 U1574 ( .A(n1231), .Y(n1232) );
  AND2X2 U1575 ( .A(n5066), .B(n1713), .Y(n1233) );
  INVX1 U1576 ( .A(n1233), .Y(n1234) );
  AND2X2 U1577 ( .A(\mem<49><6> ), .B(n3592), .Y(n1235) );
  INVX1 U1578 ( .A(n1235), .Y(n1236) );
  AND2X2 U1579 ( .A(\data_in<7> ), .B(n1713), .Y(n1237) );
  INVX1 U1580 ( .A(n1237), .Y(n1238) );
  AND2X2 U1581 ( .A(\mem<49><7> ), .B(n3592), .Y(n1239) );
  INVX1 U1582 ( .A(n1239), .Y(n1240) );
  INVX1 U1583 ( .A(n1241), .Y(n1242) );
  AND2X2 U1584 ( .A(\addr<6> ), .B(n5033), .Y(n1243) );
  INVX1 U1585 ( .A(n1243), .Y(n1244) );
  INVX1 U1586 ( .A(n5124), .Y(n1245) );
  INVX1 U1587 ( .A(n5125), .Y(n1246) );
  BUFX2 U1588 ( .A(n5176), .Y(n1247) );
  BUFX2 U1589 ( .A(n5280), .Y(n1248) );
  BUFX2 U1590 ( .A(n5342), .Y(n1249) );
  INVX1 U1591 ( .A(n5459), .Y(n1250) );
  INVX1 U1592 ( .A(n5614), .Y(n1251) );
  INVX1 U1593 ( .A(n5615), .Y(n1252) );
  BUFX2 U1594 ( .A(n5186), .Y(n1253) );
  INVX1 U1595 ( .A(n5448), .Y(n1254) );
  INVX1 U1596 ( .A(n5449), .Y(n1255) );
  INVX1 U1597 ( .A(n5625), .Y(n1256) );
  INVX1 U1598 ( .A(n5624), .Y(n1257) );
  INVX1 U1599 ( .A(n5626), .Y(n1258) );
  BUFX2 U1600 ( .A(n5752), .Y(n1259) );
  BUFX2 U1601 ( .A(n5141), .Y(n1260) );
  BUFX2 U1602 ( .A(n4803), .Y(n1261) );
  AND2X2 U1603 ( .A(n5754), .B(n3951), .Y(n1262) );
  INVX1 U1604 ( .A(n1262), .Y(n1263) );
  BUFX2 U1605 ( .A(n5351), .Y(n1264) );
  BUFX2 U1606 ( .A(n5516), .Y(n1265) );
  BUFX2 U1607 ( .A(n5429), .Y(n1266) );
  BUFX2 U1608 ( .A(n5512), .Y(n1267) );
  BUFX2 U1609 ( .A(n5602), .Y(n1268) );
  BUFX2 U1610 ( .A(n5594), .Y(n1269) );
  BUFX2 U1611 ( .A(n5685), .Y(n1270) );
  BUFX2 U1612 ( .A(n5677), .Y(n1271) );
  INVX1 U1613 ( .A(n1272), .Y(n1273) );
  AND2X2 U1614 ( .A(n4944), .B(n5275), .Y(n1274) );
  INVX1 U1615 ( .A(n1274), .Y(n1275) );
  INVX1 U1616 ( .A(n1276), .Y(n1277) );
  OR2X2 U1617 ( .A(n5467), .B(n5468), .Y(n1278) );
  INVX1 U1618 ( .A(n1278), .Y(n1279) );
  OR2X2 U1619 ( .A(n5549), .B(n5550), .Y(n1280) );
  INVX1 U1620 ( .A(n1280), .Y(n1281) );
  OR2X2 U1621 ( .A(n5633), .B(n5632), .Y(n1282) );
  INVX1 U1622 ( .A(n1282), .Y(n1283) );
  OR2X2 U1623 ( .A(n5707), .B(n5706), .Y(n1284) );
  INVX1 U1624 ( .A(n1284), .Y(n1285) );
  AND2X2 U1625 ( .A(n5039), .B(n6), .Y(n1286) );
  INVX1 U1626 ( .A(n1286), .Y(n1287) );
  AND2X2 U1627 ( .A(n5044), .B(n6), .Y(n1288) );
  INVX1 U1628 ( .A(n1288), .Y(n1289) );
  AND2X2 U1629 ( .A(n5047), .B(n6), .Y(n1290) );
  INVX1 U1630 ( .A(n1290), .Y(n1291) );
  AND2X2 U1631 ( .A(n5052), .B(n6), .Y(n1292) );
  INVX1 U1632 ( .A(n1292), .Y(n1293) );
  AND2X2 U1633 ( .A(n5057), .B(n6), .Y(n1294) );
  INVX1 U1634 ( .A(n1294), .Y(n1295) );
  AND2X2 U1635 ( .A(n5061), .B(n6), .Y(n1296) );
  INVX1 U1636 ( .A(n1296), .Y(n1297) );
  AND2X2 U1637 ( .A(n5066), .B(n6), .Y(n1298) );
  INVX1 U1638 ( .A(n1298), .Y(n1299) );
  AND2X2 U1639 ( .A(n5070), .B(n6), .Y(n1300) );
  INVX1 U1640 ( .A(n1300), .Y(n1301) );
  AND2X2 U1641 ( .A(n5039), .B(n1698), .Y(n1302) );
  INVX1 U1642 ( .A(n1302), .Y(n1303) );
  AND2X2 U1643 ( .A(n5045), .B(n1698), .Y(n1304) );
  INVX1 U1644 ( .A(n1304), .Y(n1305) );
  AND2X2 U1645 ( .A(n5047), .B(n1698), .Y(n1306) );
  INVX1 U1646 ( .A(n1306), .Y(n1307) );
  AND2X2 U1647 ( .A(n5052), .B(n1698), .Y(n1308) );
  INVX1 U1648 ( .A(n1308), .Y(n1309) );
  AND2X2 U1649 ( .A(n5057), .B(n1698), .Y(n1310) );
  INVX1 U1650 ( .A(n1310), .Y(n1311) );
  AND2X2 U1651 ( .A(n5061), .B(n1698), .Y(n1312) );
  INVX1 U1652 ( .A(n1312), .Y(n1313) );
  AND2X2 U1653 ( .A(n5066), .B(n1698), .Y(n1314) );
  INVX1 U1654 ( .A(n1314), .Y(n1315) );
  AND2X2 U1655 ( .A(n5070), .B(n1698), .Y(n1316) );
  INVX1 U1656 ( .A(n1316), .Y(n1317) );
  AND2X2 U1657 ( .A(n5039), .B(n1702), .Y(n1318) );
  INVX1 U1658 ( .A(n1318), .Y(n1319) );
  AND2X2 U1659 ( .A(n5045), .B(n1702), .Y(n1320) );
  INVX1 U1660 ( .A(n1320), .Y(n1321) );
  AND2X2 U1661 ( .A(n5048), .B(n1702), .Y(n1322) );
  INVX1 U1662 ( .A(n1322), .Y(n1323) );
  AND2X2 U1663 ( .A(n5052), .B(n1702), .Y(n1324) );
  INVX1 U1664 ( .A(n1324), .Y(n1325) );
  AND2X2 U1665 ( .A(n5057), .B(n1702), .Y(n1326) );
  INVX1 U1666 ( .A(n1326), .Y(n1327) );
  AND2X2 U1667 ( .A(n5061), .B(n1702), .Y(n1328) );
  INVX1 U1668 ( .A(n1328), .Y(n1329) );
  AND2X2 U1669 ( .A(n5066), .B(n1702), .Y(n1330) );
  INVX1 U1670 ( .A(n1330), .Y(n1331) );
  AND2X2 U1671 ( .A(n5070), .B(n1702), .Y(n1332) );
  INVX1 U1672 ( .A(n1332), .Y(n1333) );
  AND2X2 U1673 ( .A(n5039), .B(n21), .Y(n1334) );
  INVX1 U1674 ( .A(n1334), .Y(n1335) );
  AND2X2 U1675 ( .A(n5045), .B(n1707), .Y(n1336) );
  INVX1 U1676 ( .A(n1336), .Y(n1337) );
  AND2X2 U1677 ( .A(n5047), .B(n1707), .Y(n1338) );
  INVX1 U1678 ( .A(n1338), .Y(n1339) );
  AND2X2 U1679 ( .A(n5052), .B(n21), .Y(n1340) );
  INVX1 U1680 ( .A(n1340), .Y(n1341) );
  AND2X2 U1681 ( .A(n5057), .B(n21), .Y(n1342) );
  INVX1 U1682 ( .A(n1342), .Y(n1343) );
  AND2X2 U1683 ( .A(n5061), .B(n1707), .Y(n1344) );
  INVX1 U1684 ( .A(n1344), .Y(n1345) );
  AND2X2 U1685 ( .A(n5066), .B(n21), .Y(n1346) );
  INVX1 U1686 ( .A(n1346), .Y(n1347) );
  AND2X2 U1687 ( .A(n5070), .B(n1707), .Y(n1348) );
  INVX1 U1688 ( .A(n1348), .Y(n1349) );
  AND2X2 U1689 ( .A(n5039), .B(n41), .Y(n1350) );
  INVX1 U1690 ( .A(n1350), .Y(n1351) );
  AND2X2 U1691 ( .A(n5045), .B(n1709), .Y(n1352) );
  INVX1 U1692 ( .A(n1352), .Y(n1353) );
  AND2X2 U1693 ( .A(n5048), .B(n1709), .Y(n1354) );
  INVX1 U1694 ( .A(n1354), .Y(n1355) );
  AND2X2 U1695 ( .A(n5051), .B(n41), .Y(n1356) );
  INVX1 U1696 ( .A(n1356), .Y(n1357) );
  AND2X2 U1697 ( .A(n5057), .B(n41), .Y(n1358) );
  INVX1 U1698 ( .A(n1358), .Y(n1359) );
  AND2X2 U1699 ( .A(n5061), .B(n41), .Y(n1360) );
  INVX1 U1700 ( .A(n1360), .Y(n1361) );
  AND2X2 U1701 ( .A(n5066), .B(n1709), .Y(n1362) );
  INVX1 U1702 ( .A(n1362), .Y(n1363) );
  AND2X2 U1703 ( .A(n5070), .B(n1709), .Y(n1364) );
  INVX1 U1704 ( .A(n1364), .Y(n1365) );
  AND2X2 U1705 ( .A(n5039), .B(n1716), .Y(n1366) );
  INVX1 U1706 ( .A(n1366), .Y(n1367) );
  AND2X2 U1707 ( .A(n5044), .B(n1716), .Y(n1368) );
  INVX1 U1708 ( .A(n1368), .Y(n1369) );
  AND2X2 U1709 ( .A(n5048), .B(n1716), .Y(n1370) );
  INVX1 U1710 ( .A(n1370), .Y(n1371) );
  AND2X2 U1711 ( .A(n5052), .B(n42), .Y(n1372) );
  INVX1 U1712 ( .A(n1372), .Y(n1373) );
  AND2X2 U1713 ( .A(n5057), .B(n42), .Y(n1374) );
  INVX1 U1714 ( .A(n1374), .Y(n1375) );
  AND2X2 U1715 ( .A(n5061), .B(n42), .Y(n1376) );
  INVX1 U1716 ( .A(n1376), .Y(n1377) );
  AND2X2 U1717 ( .A(n5066), .B(n1716), .Y(n1378) );
  INVX1 U1718 ( .A(n1378), .Y(n1379) );
  AND2X2 U1719 ( .A(n5070), .B(n42), .Y(n1380) );
  INVX1 U1720 ( .A(n1380), .Y(n1381) );
  AND2X2 U1721 ( .A(n5039), .B(n1728), .Y(n1382) );
  INVX1 U1722 ( .A(n1382), .Y(n1383) );
  AND2X2 U1723 ( .A(n5044), .B(n1728), .Y(n1384) );
  INVX1 U1724 ( .A(n1384), .Y(n1385) );
  AND2X2 U1725 ( .A(n5047), .B(n1728), .Y(n1386) );
  INVX1 U1726 ( .A(n1386), .Y(n1387) );
  AND2X2 U1727 ( .A(n5052), .B(n1728), .Y(n1388) );
  INVX1 U1728 ( .A(n1388), .Y(n1389) );
  AND2X2 U1729 ( .A(n5057), .B(n1728), .Y(n1390) );
  INVX1 U1730 ( .A(n1390), .Y(n1391) );
  AND2X2 U1731 ( .A(n5061), .B(n1728), .Y(n1392) );
  INVX1 U1732 ( .A(n1392), .Y(n1393) );
  AND2X2 U1733 ( .A(n5066), .B(n1728), .Y(n1394) );
  INVX1 U1734 ( .A(n1394), .Y(n1395) );
  AND2X2 U1735 ( .A(n5070), .B(n1728), .Y(n1396) );
  INVX1 U1736 ( .A(n1396), .Y(n1397) );
  AND2X2 U1737 ( .A(n5039), .B(n40), .Y(n1398) );
  INVX1 U1738 ( .A(n1398), .Y(n1399) );
  AND2X2 U1739 ( .A(n5044), .B(n1730), .Y(n1400) );
  INVX1 U1740 ( .A(n1400), .Y(n1401) );
  AND2X2 U1741 ( .A(n5048), .B(n1730), .Y(n1402) );
  INVX1 U1742 ( .A(n1402), .Y(n1403) );
  AND2X2 U1743 ( .A(n5052), .B(n40), .Y(n1404) );
  INVX1 U1744 ( .A(n1404), .Y(n1405) );
  AND2X2 U1745 ( .A(n5057), .B(n1730), .Y(n1406) );
  INVX1 U1746 ( .A(n1406), .Y(n1407) );
  AND2X2 U1747 ( .A(n5061), .B(n40), .Y(n1408) );
  INVX1 U1748 ( .A(n1408), .Y(n1409) );
  AND2X2 U1749 ( .A(n5066), .B(n40), .Y(n1410) );
  INVX1 U1750 ( .A(n1410), .Y(n1411) );
  AND2X2 U1751 ( .A(n5070), .B(n1730), .Y(n1412) );
  INVX1 U1752 ( .A(n1412), .Y(n1413) );
  AND2X2 U1753 ( .A(n5038), .B(n1738), .Y(n1414) );
  INVX1 U1754 ( .A(n1414), .Y(n1415) );
  AND2X2 U1755 ( .A(n5043), .B(n1738), .Y(n1416) );
  INVX1 U1756 ( .A(n1416), .Y(n1417) );
  AND2X2 U1757 ( .A(n1738), .B(n5049), .Y(n1418) );
  INVX1 U1758 ( .A(n1418), .Y(n1419) );
  AND2X2 U1759 ( .A(n5053), .B(n1738), .Y(n1420) );
  INVX1 U1760 ( .A(n1420), .Y(n1421) );
  AND2X2 U1761 ( .A(n5055), .B(n1738), .Y(n1422) );
  INVX1 U1762 ( .A(n1422), .Y(n1423) );
  AND2X2 U1763 ( .A(n5060), .B(n1738), .Y(n1424) );
  INVX1 U1764 ( .A(n1424), .Y(n1425) );
  AND2X2 U1765 ( .A(n5064), .B(n1738), .Y(n1426) );
  INVX1 U1766 ( .A(n1426), .Y(n1427) );
  AND2X2 U1767 ( .A(n5069), .B(n1738), .Y(n1428) );
  INVX1 U1768 ( .A(n1428), .Y(n1429) );
  AND2X2 U1769 ( .A(n5038), .B(n1740), .Y(n1430) );
  INVX1 U1770 ( .A(n1430), .Y(n1431) );
  AND2X2 U1771 ( .A(n5043), .B(n1740), .Y(n1432) );
  INVX1 U1772 ( .A(n1432), .Y(n1433) );
  AND2X2 U1773 ( .A(n5049), .B(n1740), .Y(n1434) );
  INVX1 U1774 ( .A(n1434), .Y(n1435) );
  AND2X2 U1775 ( .A(n5053), .B(n1740), .Y(n1436) );
  INVX1 U1776 ( .A(n1436), .Y(n1437) );
  AND2X2 U1777 ( .A(n5056), .B(n1740), .Y(n1438) );
  INVX1 U1778 ( .A(n1438), .Y(n1439) );
  AND2X2 U1779 ( .A(n5060), .B(n1740), .Y(n1440) );
  INVX1 U1780 ( .A(n1440), .Y(n1441) );
  AND2X2 U1781 ( .A(n5065), .B(n1740), .Y(n1442) );
  INVX1 U1782 ( .A(n1442), .Y(n1443) );
  AND2X2 U1783 ( .A(n5069), .B(n1740), .Y(n1444) );
  INVX1 U1784 ( .A(n1444), .Y(n1445) );
  AND2X2 U1785 ( .A(n5038), .B(n1744), .Y(n1446) );
  INVX1 U1786 ( .A(n1446), .Y(n1447) );
  AND2X2 U1787 ( .A(n5043), .B(n1744), .Y(n1448) );
  INVX1 U1788 ( .A(n1448), .Y(n1449) );
  AND2X2 U1789 ( .A(n5049), .B(n1744), .Y(n1450) );
  INVX1 U1790 ( .A(n1450), .Y(n1451) );
  AND2X2 U1791 ( .A(n5053), .B(n1744), .Y(n1452) );
  INVX1 U1792 ( .A(n1452), .Y(n1453) );
  AND2X2 U1793 ( .A(n5055), .B(n1744), .Y(n1454) );
  INVX1 U1794 ( .A(n1454), .Y(n1455) );
  AND2X2 U1795 ( .A(n5060), .B(n1744), .Y(n1456) );
  INVX1 U1796 ( .A(n1456), .Y(n1457) );
  AND2X2 U1797 ( .A(n5064), .B(n1744), .Y(n1458) );
  INVX1 U1798 ( .A(n1458), .Y(n1459) );
  AND2X2 U1799 ( .A(n5069), .B(n1744), .Y(n1460) );
  INVX1 U1800 ( .A(n1460), .Y(n1461) );
  AND2X2 U1801 ( .A(n5038), .B(n1747), .Y(n1462) );
  INVX1 U1802 ( .A(n1462), .Y(n1463) );
  AND2X2 U1803 ( .A(n5043), .B(n1747), .Y(n1464) );
  INVX1 U1804 ( .A(n1464), .Y(n1465) );
  AND2X2 U1805 ( .A(n5049), .B(n1747), .Y(n1466) );
  INVX1 U1806 ( .A(n1466), .Y(n1467) );
  AND2X2 U1807 ( .A(n5053), .B(n1747), .Y(n1468) );
  INVX1 U1808 ( .A(n1468), .Y(n1469) );
  AND2X2 U1809 ( .A(n5056), .B(n1747), .Y(n1470) );
  INVX1 U1810 ( .A(n1470), .Y(n1471) );
  AND2X2 U1811 ( .A(n5060), .B(n1747), .Y(n1472) );
  INVX1 U1812 ( .A(n1472), .Y(n1473) );
  AND2X2 U1813 ( .A(n5065), .B(n1747), .Y(n1474) );
  INVX1 U1814 ( .A(n1474), .Y(n1475) );
  AND2X2 U1815 ( .A(n5069), .B(n1747), .Y(n1476) );
  INVX1 U1816 ( .A(n1476), .Y(n1477) );
  AND2X2 U1817 ( .A(n5038), .B(n1749), .Y(n1478) );
  INVX1 U1818 ( .A(n1478), .Y(n1479) );
  AND2X2 U1819 ( .A(n5043), .B(n1749), .Y(n1480) );
  INVX1 U1820 ( .A(n1480), .Y(n1481) );
  AND2X2 U1821 ( .A(n5049), .B(n1749), .Y(n1482) );
  INVX1 U1822 ( .A(n1482), .Y(n1483) );
  AND2X2 U1823 ( .A(n5053), .B(n1749), .Y(n1484) );
  INVX1 U1824 ( .A(n1484), .Y(n1485) );
  AND2X2 U1825 ( .A(n5055), .B(n1749), .Y(n1486) );
  INVX1 U1826 ( .A(n1486), .Y(n1487) );
  AND2X2 U1827 ( .A(n5060), .B(n1749), .Y(n1488) );
  INVX1 U1828 ( .A(n1488), .Y(n1489) );
  AND2X2 U1829 ( .A(n5065), .B(n1749), .Y(n1490) );
  INVX1 U1830 ( .A(n1490), .Y(n1491) );
  AND2X2 U1831 ( .A(n5069), .B(n1749), .Y(n1492) );
  INVX1 U1832 ( .A(n1492), .Y(n1493) );
  AND2X2 U1833 ( .A(n5038), .B(n47), .Y(n1494) );
  INVX1 U1834 ( .A(n1494), .Y(n1495) );
  AND2X2 U1835 ( .A(n5043), .B(n47), .Y(n1496) );
  INVX1 U1836 ( .A(n1496), .Y(n1497) );
  AND2X2 U1837 ( .A(n5049), .B(n1755), .Y(n1498) );
  INVX1 U1838 ( .A(n1498), .Y(n1499) );
  AND2X2 U1839 ( .A(n5053), .B(n47), .Y(n1500) );
  INVX1 U1840 ( .A(n1500), .Y(n1501) );
  AND2X2 U1841 ( .A(n5056), .B(n47), .Y(n1502) );
  INVX1 U1842 ( .A(n1502), .Y(n1503) );
  AND2X2 U1843 ( .A(n5060), .B(n1755), .Y(n1504) );
  INVX1 U1844 ( .A(n1504), .Y(n1505) );
  AND2X2 U1845 ( .A(n5064), .B(n1755), .Y(n1506) );
  INVX1 U1846 ( .A(n1506), .Y(n1507) );
  AND2X2 U1847 ( .A(n5069), .B(n1755), .Y(n1508) );
  INVX1 U1848 ( .A(n1508), .Y(n1509) );
  AND2X2 U1849 ( .A(\mem<25><4> ), .B(n3620), .Y(n1510) );
  INVX1 U1850 ( .A(n1510), .Y(n1511) );
  AND2X2 U1851 ( .A(\mem<24><4> ), .B(n3622), .Y(n1512) );
  INVX1 U1852 ( .A(n1512), .Y(n1513) );
  AND2X2 U1853 ( .A(n5038), .B(n1760), .Y(n1514) );
  INVX1 U1854 ( .A(n1514), .Y(n1515) );
  AND2X2 U1855 ( .A(n5042), .B(n1760), .Y(n1516) );
  INVX1 U1856 ( .A(n1516), .Y(n1517) );
  AND2X2 U1857 ( .A(n5048), .B(n1760), .Y(n1518) );
  INVX1 U1858 ( .A(n1518), .Y(n1519) );
  AND2X2 U1859 ( .A(n5052), .B(n1760), .Y(n1520) );
  INVX1 U1860 ( .A(n1520), .Y(n1521) );
  AND2X2 U1861 ( .A(n5056), .B(n1760), .Y(n1522) );
  INVX1 U1862 ( .A(n1522), .Y(n1523) );
  AND2X2 U1863 ( .A(n5060), .B(n1760), .Y(n1524) );
  INVX1 U1864 ( .A(n1524), .Y(n1525) );
  AND2X2 U1865 ( .A(n5065), .B(n1760), .Y(n1526) );
  INVX1 U1866 ( .A(n1526), .Y(n1527) );
  AND2X2 U1867 ( .A(n5069), .B(n1760), .Y(n1528) );
  INVX1 U1868 ( .A(n1528), .Y(n1529) );
  AND2X2 U1869 ( .A(n5038), .B(n1766), .Y(n1530) );
  INVX1 U1870 ( .A(n1530), .Y(n1531) );
  AND2X2 U1871 ( .A(n5042), .B(n1766), .Y(n1532) );
  INVX1 U1872 ( .A(n1532), .Y(n1533) );
  AND2X2 U1873 ( .A(n5048), .B(n1766), .Y(n1534) );
  INVX1 U1874 ( .A(n1534), .Y(n1535) );
  AND2X2 U1875 ( .A(n5052), .B(n1766), .Y(n1536) );
  INVX1 U1876 ( .A(n1536), .Y(n1537) );
  AND2X2 U1877 ( .A(n5056), .B(n1766), .Y(n1538) );
  INVX1 U1878 ( .A(n1538), .Y(n1539) );
  AND2X2 U1879 ( .A(n5060), .B(n1766), .Y(n1540) );
  INVX1 U1880 ( .A(n1540), .Y(n1541) );
  AND2X2 U1881 ( .A(n5065), .B(n1766), .Y(n1542) );
  INVX1 U1882 ( .A(n1542), .Y(n1543) );
  AND2X2 U1883 ( .A(n5069), .B(n1766), .Y(n1544) );
  INVX1 U1884 ( .A(n1544), .Y(n1545) );
  AND2X2 U1885 ( .A(n5038), .B(n1768), .Y(n1546) );
  INVX1 U1886 ( .A(n1546), .Y(n1547) );
  AND2X2 U1887 ( .A(n5042), .B(n1768), .Y(n1548) );
  INVX1 U1888 ( .A(n1548), .Y(n1549) );
  AND2X2 U1889 ( .A(n5048), .B(n1768), .Y(n1550) );
  INVX1 U1890 ( .A(n1550), .Y(n1551) );
  AND2X2 U1891 ( .A(n5052), .B(n1768), .Y(n1552) );
  INVX1 U1892 ( .A(n1552), .Y(n1553) );
  AND2X2 U1893 ( .A(n5056), .B(n1768), .Y(n1554) );
  INVX1 U1894 ( .A(n1554), .Y(n1555) );
  AND2X2 U1895 ( .A(n5060), .B(n1768), .Y(n1556) );
  INVX1 U1896 ( .A(n1556), .Y(n1557) );
  AND2X2 U1897 ( .A(n5065), .B(n1768), .Y(n1558) );
  INVX1 U1898 ( .A(n1558), .Y(n1559) );
  AND2X2 U1899 ( .A(n5069), .B(n1768), .Y(n1560) );
  INVX1 U1900 ( .A(n1560), .Y(n1561) );
  AND2X2 U1901 ( .A(n5052), .B(n1774), .Y(n1562) );
  INVX1 U1902 ( .A(n1562), .Y(n1563) );
  AND2X2 U1903 ( .A(n5056), .B(n1774), .Y(n1564) );
  INVX1 U1904 ( .A(n1564), .Y(n1565) );
  AND2X2 U1905 ( .A(n5060), .B(n1774), .Y(n1566) );
  INVX1 U1906 ( .A(n1566), .Y(n1567) );
  AND2X2 U1907 ( .A(n5065), .B(n1774), .Y(n1568) );
  INVX1 U1908 ( .A(n1568), .Y(n1569) );
  AND2X2 U1909 ( .A(n5069), .B(n1774), .Y(n1570) );
  INVX1 U1910 ( .A(n1570), .Y(n1571) );
  AND2X2 U1911 ( .A(n5038), .B(n1775), .Y(n1572) );
  INVX1 U1912 ( .A(n1572), .Y(n1573) );
  AND2X2 U1913 ( .A(n5042), .B(n102), .Y(n1574) );
  INVX1 U1914 ( .A(n1574), .Y(n1575) );
  AND2X2 U1915 ( .A(n5048), .B(n1775), .Y(n1576) );
  INVX1 U1916 ( .A(n1576), .Y(n1577) );
  AND2X2 U1917 ( .A(n5052), .B(n102), .Y(n1578) );
  INVX1 U1918 ( .A(n1578), .Y(n1579) );
  AND2X2 U1919 ( .A(n5056), .B(n102), .Y(n1580) );
  INVX1 U1920 ( .A(n1580), .Y(n1581) );
  AND2X2 U1921 ( .A(n5060), .B(n102), .Y(n1582) );
  INVX1 U1922 ( .A(n1582), .Y(n1583) );
  AND2X2 U1923 ( .A(n5065), .B(n1775), .Y(n1584) );
  INVX1 U1924 ( .A(n1584), .Y(n1585) );
  AND2X2 U1925 ( .A(n5069), .B(n1775), .Y(n1586) );
  INVX1 U1926 ( .A(n1586), .Y(n1587) );
  AND2X2 U1927 ( .A(n5038), .B(n1781), .Y(n1588) );
  INVX1 U1928 ( .A(n1588), .Y(n1589) );
  AND2X2 U1929 ( .A(n5041), .B(n1781), .Y(n1590) );
  INVX1 U1930 ( .A(n1590), .Y(n1591) );
  AND2X2 U1931 ( .A(n5047), .B(n1781), .Y(n1592) );
  INVX1 U1932 ( .A(n1592), .Y(n1593) );
  AND2X2 U1933 ( .A(n5051), .B(n1781), .Y(n1594) );
  INVX1 U1934 ( .A(n1594), .Y(n1595) );
  AND2X2 U1935 ( .A(n5055), .B(n1781), .Y(n1596) );
  INVX1 U1936 ( .A(n1596), .Y(n1597) );
  AND2X2 U1937 ( .A(n5060), .B(n1781), .Y(n1598) );
  INVX1 U1938 ( .A(n1598), .Y(n1599) );
  AND2X2 U1939 ( .A(n5064), .B(n1781), .Y(n1600) );
  INVX1 U1940 ( .A(n1600), .Y(n1601) );
  AND2X2 U1941 ( .A(n5069), .B(n1781), .Y(n1602) );
  INVX1 U1942 ( .A(n1602), .Y(n1603) );
  AND2X2 U1943 ( .A(n5038), .B(n1783), .Y(n1604) );
  INVX1 U1944 ( .A(n1604), .Y(n1605) );
  AND2X2 U1945 ( .A(n5041), .B(n1783), .Y(n1606) );
  INVX1 U1946 ( .A(n1606), .Y(n1607) );
  AND2X2 U1947 ( .A(n5047), .B(n1783), .Y(n1608) );
  INVX1 U1948 ( .A(n1608), .Y(n1609) );
  AND2X2 U1949 ( .A(n5051), .B(n1783), .Y(n1610) );
  INVX1 U1950 ( .A(n1610), .Y(n1611) );
  AND2X2 U1951 ( .A(n5055), .B(n1783), .Y(n1612) );
  INVX1 U1952 ( .A(n1612), .Y(n1613) );
  AND2X2 U1953 ( .A(n5060), .B(n1783), .Y(n1614) );
  INVX1 U1954 ( .A(n1614), .Y(n1615) );
  AND2X2 U1955 ( .A(n5064), .B(n1783), .Y(n1616) );
  INVX1 U1956 ( .A(n1616), .Y(n1617) );
  AND2X2 U1957 ( .A(n5069), .B(n1783), .Y(n1618) );
  INVX1 U1958 ( .A(n1618), .Y(n1619) );
  AND2X2 U1959 ( .A(n5038), .B(n1789), .Y(n1620) );
  INVX1 U1960 ( .A(n1620), .Y(n1621) );
  AND2X2 U1961 ( .A(n5041), .B(n1789), .Y(n1622) );
  INVX1 U1962 ( .A(n1622), .Y(n1623) );
  AND2X2 U1963 ( .A(n5047), .B(n1789), .Y(n1624) );
  INVX1 U1964 ( .A(n1624), .Y(n1625) );
  AND2X2 U1965 ( .A(n5051), .B(n1789), .Y(n1626) );
  INVX1 U1966 ( .A(n1626), .Y(n1627) );
  AND2X2 U1967 ( .A(n5055), .B(n1789), .Y(n1628) );
  INVX1 U1968 ( .A(n1628), .Y(n1629) );
  AND2X2 U1969 ( .A(n5060), .B(n1789), .Y(n1630) );
  INVX1 U1970 ( .A(n1630), .Y(n1631) );
  AND2X2 U1971 ( .A(n5064), .B(n1789), .Y(n1632) );
  INVX1 U1972 ( .A(n1632), .Y(n1633) );
  AND2X2 U1973 ( .A(n5108), .B(n1790), .Y(n1634) );
  INVX1 U1974 ( .A(n1634), .Y(n1635) );
  AND2X2 U1975 ( .A(n5038), .B(n1797), .Y(n1636) );
  INVX1 U1976 ( .A(n1636), .Y(n1637) );
  AND2X2 U1977 ( .A(n5041), .B(n1797), .Y(n1638) );
  INVX1 U1978 ( .A(n1638), .Y(n1639) );
  AND2X2 U1979 ( .A(n5047), .B(n1797), .Y(n1640) );
  INVX1 U1980 ( .A(n1640), .Y(n1641) );
  AND2X2 U1981 ( .A(n5051), .B(n1797), .Y(n1642) );
  INVX1 U1982 ( .A(n1642), .Y(n1643) );
  AND2X2 U1983 ( .A(n5055), .B(n1797), .Y(n1644) );
  INVX1 U1984 ( .A(n1644), .Y(n1645) );
  AND2X2 U1985 ( .A(n5060), .B(n1797), .Y(n1646) );
  INVX1 U1986 ( .A(n1646), .Y(n1647) );
  AND2X2 U1987 ( .A(n5064), .B(n1797), .Y(n1648) );
  INVX1 U1988 ( .A(n1648), .Y(n1649) );
  AND2X2 U1989 ( .A(n5069), .B(n1797), .Y(n1650) );
  INVX1 U1990 ( .A(n1650), .Y(n1651) );
  AND2X2 U1991 ( .A(n5038), .B(n53), .Y(n1652) );
  INVX1 U1992 ( .A(n1652), .Y(n1653) );
  AND2X2 U1993 ( .A(n5041), .B(n1799), .Y(n1654) );
  INVX1 U1994 ( .A(n1654), .Y(n1655) );
  AND2X2 U1995 ( .A(n5047), .B(n1799), .Y(n1656) );
  INVX1 U1996 ( .A(n1656), .Y(n1657) );
  AND2X2 U1997 ( .A(n5051), .B(n1799), .Y(n1658) );
  INVX1 U1998 ( .A(n1658), .Y(n1659) );
  AND2X2 U1999 ( .A(n5055), .B(n53), .Y(n1660) );
  INVX1 U2000 ( .A(n1660), .Y(n1661) );
  AND2X2 U2001 ( .A(n5060), .B(n1799), .Y(n1662) );
  INVX1 U2002 ( .A(n1662), .Y(n1663) );
  AND2X2 U2003 ( .A(n5064), .B(n53), .Y(n1664) );
  INVX1 U2004 ( .A(n1664), .Y(n1665) );
  AND2X2 U2005 ( .A(n5069), .B(n53), .Y(n1666) );
  INVX1 U2006 ( .A(n1666), .Y(n1667) );
  AND2X2 U2007 ( .A(\mem<1><0> ), .B(n6419), .Y(n1668) );
  INVX1 U2008 ( .A(n1668), .Y(n1669) );
  AND2X2 U2009 ( .A(\mem<1><1> ), .B(n6419), .Y(n1670) );
  INVX1 U2010 ( .A(n1670), .Y(n1671) );
  AND2X2 U2011 ( .A(\mem<1><2> ), .B(n6419), .Y(n1672) );
  INVX1 U2012 ( .A(n1672), .Y(n1673) );
  AND2X2 U2013 ( .A(\mem<1><3> ), .B(n6419), .Y(n1674) );
  INVX1 U2014 ( .A(n1674), .Y(n1675) );
  AND2X2 U2015 ( .A(\mem<1><4> ), .B(n6419), .Y(n1676) );
  INVX1 U2016 ( .A(n1676), .Y(n1677) );
  AND2X2 U2017 ( .A(\mem<1><5> ), .B(n6419), .Y(n1678) );
  INVX1 U2018 ( .A(n1678), .Y(n1679) );
  AND2X2 U2019 ( .A(\mem<1><6> ), .B(n6419), .Y(n1680) );
  INVX1 U2020 ( .A(n1680), .Y(n1681) );
  AND2X2 U2021 ( .A(\mem<1><7> ), .B(n6419), .Y(n1682) );
  INVX1 U2022 ( .A(n1682), .Y(n1683) );
  BUFX2 U2023 ( .A(n3852), .Y(n1684) );
  BUFX2 U2024 ( .A(n3859), .Y(n1685) );
  BUFX2 U2025 ( .A(n6291), .Y(n1686) );
  BUFX2 U2026 ( .A(n6390), .Y(n1687) );
  AND2X2 U2027 ( .A(n6290), .B(n6405), .Y(n1689) );
  AND2X2 U2028 ( .A(n112), .B(n6294), .Y(n1690) );
  AND2X2 U2029 ( .A(n4624), .B(n6294), .Y(n1691) );
  AND2X2 U2030 ( .A(n3665), .B(n87), .Y(n1692) );
  AND2X2 U2031 ( .A(n87), .B(n4), .Y(n1693) );
  AND2X2 U2032 ( .A(n4674), .B(n6297), .Y(n1694) );
  AND2X2 U2033 ( .A(n6297), .B(n6298), .Y(n1695) );
  AND2X2 U2034 ( .A(n6300), .B(n3864), .Y(n1696) );
  AND2X2 U2035 ( .A(n6300), .B(n6302), .Y(n1697) );
  AND2X2 U2036 ( .A(n6303), .B(n3579), .Y(n1698) );
  AND2X2 U2037 ( .A(n3652), .B(n3579), .Y(n1699) );
  AND2X2 U2038 ( .A(n4682), .B(n3581), .Y(n1700) );
  AND2X2 U2039 ( .A(n4719), .B(n3581), .Y(n1701) );
  AND2X2 U2040 ( .A(n3583), .B(n3873), .Y(n1702) );
  AND2X2 U2041 ( .A(n4653), .B(n3583), .Y(n1703) );
  AND2X2 U2042 ( .A(n6405), .B(n6305), .Y(n1704) );
  AND2X2 U2043 ( .A(n6306), .B(n6305), .Y(n1705) );
  AND2X2 U2044 ( .A(n6309), .B(n112), .Y(n1706) );
  AND2X2 U2045 ( .A(n4875), .B(n3585), .Y(n1707) );
  AND2X2 U2046 ( .A(n6313), .B(n3585), .Y(n1708) );
  AND2X2 U2047 ( .A(n4674), .B(n3587), .Y(n1709) );
  AND2X2 U2048 ( .A(n26), .B(n3587), .Y(n1710) );
  AND2X2 U2049 ( .A(n3668), .B(n3589), .Y(n1711) );
  AND2X2 U2050 ( .A(n3669), .B(n3589), .Y(n1712) );
  AND2X2 U2051 ( .A(n4824), .B(n3591), .Y(n1713) );
  AND2X2 U2052 ( .A(n6315), .B(n3593), .Y(n1714) );
  AND2X2 U2053 ( .A(n3593), .B(n96), .Y(n1715) );
  AND2X2 U2054 ( .A(n3873), .B(n3595), .Y(n1716) );
  AND2X2 U2055 ( .A(n4654), .B(n3595), .Y(n1717) );
  AND2X2 U2056 ( .A(n6325), .B(n6405), .Y(n1718) );
  AND2X2 U2057 ( .A(n6325), .B(n25), .Y(n1719) );
  AND2X2 U2058 ( .A(n112), .B(n1685), .Y(n1720) );
  AND2X2 U2059 ( .A(n4655), .B(n1685), .Y(n1721) );
  AND2X2 U2060 ( .A(n574), .B(n3597), .Y(n1722) );
  AND2X2 U2061 ( .A(n6330), .B(n3597), .Y(n1723) );
  AND2X2 U2062 ( .A(n3599), .B(n4674), .Y(n1724) );
  AND2X2 U2063 ( .A(n3599), .B(n19), .Y(n1725) );
  AND2X2 U2064 ( .A(n6331), .B(n3601), .Y(n1726) );
  AND2X2 U2065 ( .A(n1684), .B(n3601), .Y(n1727) );
  AND2X2 U2066 ( .A(n36), .B(n3603), .Y(n1728) );
  AND2X2 U2067 ( .A(n3881), .B(n3603), .Y(n1729) );
  AND2X2 U2068 ( .A(n4680), .B(n3605), .Y(n1730) );
  AND2X2 U2069 ( .A(n4649), .B(n3605), .Y(n1731) );
  AND2X2 U2070 ( .A(n4965), .B(n3607), .Y(n1732) );
  AND2X2 U2071 ( .A(n3607), .B(n4656), .Y(n1733) );
  AND2X2 U2072 ( .A(n6405), .B(n6336), .Y(n1734) );
  AND2X2 U2073 ( .A(n6336), .B(n6337), .Y(n1735) );
  AND2X2 U2074 ( .A(n6340), .B(n64), .Y(n1736) );
  AND2X2 U2075 ( .A(n6340), .B(n4657), .Y(n1737) );
  AND2X2 U2076 ( .A(n4846), .B(n3609), .Y(n1738) );
  AND2X2 U2077 ( .A(n6342), .B(n3609), .Y(n1739) );
  AND2X2 U2078 ( .A(n4674), .B(n3611), .Y(n1740) );
  AND2X2 U2079 ( .A(n4636), .B(n3611), .Y(n1741) );
  AND2X2 U2080 ( .A(n6343), .B(n3613), .Y(n1742) );
  AND2X2 U2081 ( .A(n6344), .B(n3613), .Y(n1743) );
  AND2X2 U2082 ( .A(n3615), .B(n4822), .Y(n1744) );
  AND2X2 U2083 ( .A(n6345), .B(n3615), .Y(n1745) );
  AND2X2 U2084 ( .A(n6346), .B(n804), .Y(n1746) );
  AND2X2 U2085 ( .A(n6349), .B(n3873), .Y(n1747) );
  AND2X2 U2086 ( .A(n6350), .B(n6349), .Y(n1748) );
  AND2X2 U2087 ( .A(n6359), .B(n4966), .Y(n1749) );
  AND2X2 U2088 ( .A(n4651), .B(n6359), .Y(n1750) );
  AND2X2 U2089 ( .A(n6363), .B(n6360), .Y(n1751) );
  AND2X2 U2090 ( .A(n6360), .B(n4857), .Y(n1752) );
  AND2X2 U2091 ( .A(n4674), .B(n6364), .Y(n1753) );
  AND2X2 U2092 ( .A(n4664), .B(n6364), .Y(n1754) );
  AND2X2 U2093 ( .A(n6366), .B(n3617), .Y(n1755) );
  AND2X2 U2094 ( .A(n4918), .B(n3617), .Y(n1756) );
  AND2X2 U2095 ( .A(n3856), .B(n3619), .Y(n1757) );
  AND2X2 U2096 ( .A(n4849), .B(n3619), .Y(n1758) );
  AND2X2 U2097 ( .A(n3867), .B(n3621), .Y(n1759) );
  AND2X2 U2098 ( .A(n4965), .B(n3623), .Y(n1760) );
  AND2X2 U2099 ( .A(n3560), .B(n3623), .Y(n1761) );
  AND2X2 U2100 ( .A(n6405), .B(n6371), .Y(n1762) );
  AND2X2 U2101 ( .A(n6372), .B(n6371), .Y(n1763) );
  AND2X2 U2102 ( .A(n64), .B(n6375), .Y(n1764) );
  AND2X2 U2103 ( .A(n4658), .B(n6375), .Y(n1765) );
  AND2X2 U2104 ( .A(n6377), .B(n3625), .Y(n1766) );
  AND2X2 U2105 ( .A(n6378), .B(n3625), .Y(n1767) );
  AND2X2 U2106 ( .A(n4674), .B(n3627), .Y(n1768) );
  AND2X2 U2107 ( .A(n4641), .B(n3627), .Y(n1769) );
  AND2X2 U2108 ( .A(n4911), .B(n3629), .Y(n1770) );
  AND2X2 U2109 ( .A(n4823), .B(n3629), .Y(n1771) );
  AND2X2 U2110 ( .A(n6387), .B(n3631), .Y(n1772) );
  AND2X2 U2111 ( .A(n13), .B(n3631), .Y(n1773) );
  AND2X2 U2112 ( .A(n4816), .B(n3651), .Y(n1774) );
  AND2X2 U2113 ( .A(n4965), .B(n3633), .Y(n1775) );
  AND2X2 U2114 ( .A(n4661), .B(n3633), .Y(n1776) );
  AND2X2 U2115 ( .A(n6405), .B(n6391), .Y(n1777) );
  AND2X2 U2116 ( .A(n6392), .B(n6391), .Y(n1778) );
  AND2X2 U2117 ( .A(n64), .B(n6395), .Y(n1779) );
  AND2X2 U2118 ( .A(n4662), .B(n6395), .Y(n1780) );
  AND2X2 U2119 ( .A(n3654), .B(n3869), .Y(n1781) );
  AND2X2 U2120 ( .A(n4829), .B(n3869), .Y(n1782) );
  AND2X2 U2121 ( .A(n4674), .B(n3666), .Y(n1783) );
  AND2X2 U2122 ( .A(n4645), .B(n3666), .Y(n1784) );
  AND2X2 U2123 ( .A(n3635), .B(n6399), .Y(n1785) );
  AND2X2 U2124 ( .A(n4828), .B(n3635), .Y(n1786) );
  AND2X2 U2125 ( .A(n3863), .B(n3637), .Y(n1787) );
  AND2X2 U2126 ( .A(n3637), .B(n14), .Y(n1788) );
  AND2X2 U2127 ( .A(n6402), .B(n3639), .Y(n1789) );
  AND2X2 U2128 ( .A(n4870), .B(n3639), .Y(n1790) );
  AND2X2 U2129 ( .A(n3641), .B(n3873), .Y(n1791) );
  AND2X2 U2130 ( .A(n3562), .B(n3641), .Y(n1792) );
  AND2X2 U2131 ( .A(n6405), .B(n6406), .Y(n1793) );
  AND2X2 U2132 ( .A(n6407), .B(n6406), .Y(n1794) );
  AND2X2 U2133 ( .A(n4966), .B(n6411), .Y(n1795) );
  AND2X2 U2134 ( .A(n6411), .B(n4663), .Y(n1796) );
  AND2X2 U2135 ( .A(n6413), .B(n3643), .Y(n1797) );
  AND2X2 U2136 ( .A(n6414), .B(n3643), .Y(n1798) );
  AND2X2 U2137 ( .A(n4674), .B(n3645), .Y(n1799) );
  AND2X2 U2138 ( .A(n4647), .B(n3645), .Y(n1800) );
  AND2X2 U2139 ( .A(n108), .B(n3647), .Y(n1801) );
  AND2X2 U2140 ( .A(n78), .B(n3647), .Y(n1802) );
  AND2X2 U2141 ( .A(n4810), .B(n6418), .Y(n1803) );
  INVX1 U2142 ( .A(n5307), .Y(n1804) );
  INVX1 U2143 ( .A(n5308), .Y(n1805) );
  INVX1 U2144 ( .A(n5309), .Y(n1806) );
  OR2X2 U2145 ( .A(n1253), .B(n722), .Y(n1807) );
  INVX1 U2146 ( .A(n1807), .Y(n1808) );
  OR2X2 U2147 ( .A(n724), .B(n728), .Y(n1809) );
  INVX1 U2148 ( .A(n1809), .Y(n1810) );
  OR2X2 U2149 ( .A(n726), .B(n730), .Y(n1811) );
  INVX1 U2150 ( .A(n1811), .Y(n1812) );
  OR2X2 U2151 ( .A(n5753), .B(n1259), .Y(n1813) );
  INVX1 U2152 ( .A(n1813), .Y(n1814) );
  AND2X2 U2153 ( .A(\mem<59><0> ), .B(n4946), .Y(n1815) );
  INVX1 U2154 ( .A(n1815), .Y(n2328) );
  AND2X2 U2155 ( .A(\mem<63><6> ), .B(n4946), .Y(n2329) );
  INVX1 U2156 ( .A(n2329), .Y(n2330) );
  AND2X2 U2157 ( .A(\mem<61><6> ), .B(n4946), .Y(n2331) );
  INVX1 U2158 ( .A(n2331), .Y(n2332) );
  INVX1 U2159 ( .A(n5154), .Y(n2333) );
  INVX1 U2160 ( .A(n5155), .Y(n2334) );
  INVX1 U2161 ( .A(n5156), .Y(n2335) );
  INVX1 U2162 ( .A(n5321), .Y(n2336) );
  INVX1 U2163 ( .A(n5322), .Y(n2337) );
  INVX1 U2164 ( .A(n5323), .Y(n2338) );
  INVX1 U2165 ( .A(n5493), .Y(n2339) );
  INVX1 U2166 ( .A(n5494), .Y(n2340) );
  INVX1 U2167 ( .A(n5576), .Y(n2341) );
  INVX1 U2168 ( .A(n5577), .Y(n2342) );
  INVX1 U2169 ( .A(n5578), .Y(n2343) );
  INVX1 U2170 ( .A(n5658), .Y(n2344) );
  INVX1 U2171 ( .A(n5659), .Y(n2345) );
  INVX1 U2172 ( .A(n5660), .Y(n2346) );
  BUFX2 U2173 ( .A(n5436), .Y(n2347) );
  BUFX2 U2174 ( .A(n5601), .Y(n2348) );
  BUFX2 U2175 ( .A(n5684), .Y(n2349) );
  BUFX2 U2176 ( .A(n5289), .Y(n2350) );
  BUFX2 U2177 ( .A(n5517), .Y(n2351) );
  OR2X2 U2178 ( .A(\addr<8> ), .B(\addr<7> ), .Y(n2352) );
  OR2X2 U2179 ( .A(n807), .B(n5008), .Y(n2353) );
  INVX1 U2180 ( .A(n2353), .Y(n2354) );
  AND2X2 U2181 ( .A(\mem<22><0> ), .B(n4957), .Y(n2355) );
  INVX1 U2182 ( .A(n2355), .Y(n2356) );
  AND2X2 U2183 ( .A(n4891), .B(n5276), .Y(n2357) );
  INVX1 U2184 ( .A(n2357), .Y(n2358) );
  AND2X2 U2185 ( .A(\mem<22><2> ), .B(n4957), .Y(n2359) );
  INVX1 U2186 ( .A(n2359), .Y(n2360) );
  AND2X2 U2187 ( .A(n5072), .B(n1688), .Y(n2361) );
  INVX1 U2188 ( .A(n2361), .Y(n2362) );
  AND2X2 U2189 ( .A(n5078), .B(n1688), .Y(n2363) );
  INVX1 U2190 ( .A(n2363), .Y(n2364) );
  AND2X2 U2191 ( .A(n5084), .B(n1688), .Y(n2365) );
  INVX1 U2192 ( .A(n2365), .Y(n2366) );
  AND2X2 U2193 ( .A(n5089), .B(n1688), .Y(n2367) );
  INVX1 U2194 ( .A(n2367), .Y(n2368) );
  AND2X2 U2195 ( .A(n5095), .B(n1688), .Y(n2369) );
  INVX1 U2196 ( .A(n2369), .Y(n2370) );
  AND2X2 U2197 ( .A(n5099), .B(n1688), .Y(n2371) );
  INVX1 U2198 ( .A(n2371), .Y(n2372) );
  AND2X2 U2199 ( .A(n5103), .B(n1688), .Y(n2373) );
  INVX1 U2200 ( .A(n2373), .Y(n2374) );
  AND2X2 U2201 ( .A(n5108), .B(n1688), .Y(n2375) );
  INVX1 U2202 ( .A(n2375), .Y(n2376) );
  AND2X2 U2203 ( .A(n5072), .B(n1691), .Y(n2377) );
  INVX1 U2204 ( .A(n2377), .Y(n2378) );
  AND2X2 U2205 ( .A(n5078), .B(n1691), .Y(n2379) );
  INVX1 U2206 ( .A(n2379), .Y(n2380) );
  AND2X2 U2207 ( .A(n5084), .B(n1691), .Y(n2381) );
  INVX1 U2208 ( .A(n2381), .Y(n2382) );
  AND2X2 U2209 ( .A(n5089), .B(n1691), .Y(n2383) );
  INVX1 U2210 ( .A(n2383), .Y(n2384) );
  AND2X2 U2211 ( .A(n5095), .B(n1691), .Y(n2385) );
  INVX1 U2212 ( .A(n2385), .Y(n2386) );
  AND2X2 U2213 ( .A(n5099), .B(n1691), .Y(n2387) );
  INVX1 U2214 ( .A(n2387), .Y(n2388) );
  AND2X2 U2215 ( .A(n5103), .B(n1691), .Y(n2389) );
  INVX1 U2216 ( .A(n2389), .Y(n2390) );
  AND2X2 U2217 ( .A(n5108), .B(n1691), .Y(n2391) );
  INVX1 U2218 ( .A(n2391), .Y(n2392) );
  AND2X2 U2219 ( .A(n5072), .B(n1697), .Y(n2393) );
  INVX1 U2220 ( .A(n2393), .Y(n2394) );
  AND2X2 U2221 ( .A(n5078), .B(n1697), .Y(n2395) );
  INVX1 U2222 ( .A(n2395), .Y(n2396) );
  AND2X2 U2223 ( .A(n5084), .B(n1697), .Y(n2397) );
  INVX1 U2224 ( .A(n2397), .Y(n2398) );
  AND2X2 U2225 ( .A(n5089), .B(n1697), .Y(n2399) );
  INVX1 U2226 ( .A(n2399), .Y(n2400) );
  AND2X2 U2227 ( .A(n5095), .B(n1697), .Y(n2401) );
  INVX1 U2228 ( .A(n2401), .Y(n2402) );
  AND2X2 U2229 ( .A(n5099), .B(n1697), .Y(n2403) );
  INVX1 U2230 ( .A(n2403), .Y(n2404) );
  AND2X2 U2231 ( .A(n5103), .B(n1697), .Y(n2405) );
  INVX1 U2232 ( .A(n2405), .Y(n2406) );
  AND2X2 U2233 ( .A(n5107), .B(n1697), .Y(n2407) );
  INVX1 U2234 ( .A(n2407), .Y(n2408) );
  AND2X2 U2235 ( .A(n5072), .B(n1703), .Y(n2409) );
  INVX1 U2236 ( .A(n2409), .Y(n2410) );
  AND2X2 U2237 ( .A(n5078), .B(n1703), .Y(n2411) );
  INVX1 U2238 ( .A(n2411), .Y(n2412) );
  AND2X2 U2239 ( .A(n5084), .B(n1703), .Y(n2413) );
  INVX1 U2240 ( .A(n2413), .Y(n2414) );
  AND2X2 U2241 ( .A(n5089), .B(n1703), .Y(n2415) );
  INVX1 U2242 ( .A(n2415), .Y(n2416) );
  AND2X2 U2243 ( .A(n5095), .B(n1703), .Y(n2417) );
  INVX1 U2244 ( .A(n2417), .Y(n2418) );
  AND2X2 U2245 ( .A(n5099), .B(n1703), .Y(n2419) );
  INVX1 U2246 ( .A(n2419), .Y(n2420) );
  AND2X2 U2247 ( .A(n5103), .B(n1703), .Y(n2421) );
  INVX1 U2248 ( .A(n2421), .Y(n2422) );
  AND2X2 U2249 ( .A(n5108), .B(n1703), .Y(n2423) );
  INVX1 U2250 ( .A(n2423), .Y(n2424) );
  AND2X2 U2251 ( .A(n5072), .B(n1705), .Y(n2425) );
  INVX1 U2252 ( .A(n2425), .Y(n2426) );
  AND2X2 U2253 ( .A(n5078), .B(n1705), .Y(n2427) );
  INVX1 U2254 ( .A(n2427), .Y(n2428) );
  AND2X2 U2255 ( .A(n5084), .B(n1705), .Y(n2429) );
  INVX1 U2256 ( .A(n2429), .Y(n2430) );
  AND2X2 U2257 ( .A(n5089), .B(n1705), .Y(n2431) );
  INVX1 U2258 ( .A(n2431), .Y(n2432) );
  AND2X2 U2259 ( .A(n5095), .B(n1705), .Y(n2433) );
  INVX1 U2260 ( .A(n2433), .Y(n2434) );
  AND2X2 U2261 ( .A(n5099), .B(n1705), .Y(n2435) );
  INVX1 U2262 ( .A(n2435), .Y(n2436) );
  AND2X2 U2263 ( .A(n5103), .B(n1705), .Y(n2437) );
  INVX1 U2264 ( .A(n2437), .Y(n2438) );
  AND2X2 U2265 ( .A(n5107), .B(n1705), .Y(n2439) );
  INVX1 U2266 ( .A(n2439), .Y(n2440) );
  AND2X2 U2267 ( .A(n5072), .B(n1708), .Y(n2441) );
  INVX1 U2268 ( .A(n2441), .Y(n2442) );
  AND2X2 U2269 ( .A(n5078), .B(n1708), .Y(n2443) );
  INVX1 U2270 ( .A(n2443), .Y(n2444) );
  AND2X2 U2271 ( .A(n5084), .B(n1708), .Y(n2445) );
  INVX1 U2272 ( .A(n2445), .Y(n2446) );
  AND2X2 U2273 ( .A(n5089), .B(n1708), .Y(n2447) );
  INVX1 U2274 ( .A(n2447), .Y(n2448) );
  AND2X2 U2275 ( .A(n5095), .B(n1708), .Y(n2449) );
  INVX1 U2276 ( .A(n2449), .Y(n2450) );
  AND2X2 U2277 ( .A(n5099), .B(n1708), .Y(n2451) );
  INVX1 U2278 ( .A(n2451), .Y(n2452) );
  AND2X2 U2279 ( .A(n5103), .B(n1708), .Y(n2453) );
  INVX1 U2280 ( .A(n2453), .Y(n2454) );
  AND2X2 U2281 ( .A(n5108), .B(n1708), .Y(n2455) );
  INVX1 U2282 ( .A(n2455), .Y(n2456) );
  AND2X2 U2283 ( .A(n5072), .B(n1710), .Y(n2457) );
  INVX1 U2284 ( .A(n2457), .Y(n2458) );
  AND2X2 U2285 ( .A(n5077), .B(n1710), .Y(n2459) );
  INVX1 U2286 ( .A(n2459), .Y(n2460) );
  AND2X2 U2287 ( .A(n5082), .B(n1710), .Y(n2461) );
  INVX1 U2288 ( .A(n2461), .Y(n2462) );
  AND2X2 U2289 ( .A(n5089), .B(n1710), .Y(n2463) );
  INVX1 U2290 ( .A(n2463), .Y(n2464) );
  AND2X2 U2291 ( .A(n5094), .B(n1710), .Y(n2465) );
  INVX1 U2292 ( .A(n2465), .Y(n2466) );
  AND2X2 U2293 ( .A(n5098), .B(n1710), .Y(n2467) );
  INVX1 U2294 ( .A(n2467), .Y(n2468) );
  AND2X2 U2295 ( .A(n5102), .B(n1710), .Y(n2469) );
  INVX1 U2296 ( .A(n2469), .Y(n2470) );
  AND2X2 U2297 ( .A(n5108), .B(n1710), .Y(n2471) );
  INVX1 U2298 ( .A(n2471), .Y(n2472) );
  AND2X2 U2299 ( .A(n5072), .B(n1712), .Y(n2473) );
  INVX1 U2300 ( .A(n2473), .Y(n2474) );
  AND2X2 U2301 ( .A(n5077), .B(n1712), .Y(n2475) );
  INVX1 U2302 ( .A(n2475), .Y(n2476) );
  AND2X2 U2303 ( .A(n5082), .B(n1712), .Y(n2477) );
  INVX1 U2304 ( .A(n2477), .Y(n2478) );
  AND2X2 U2305 ( .A(n5089), .B(n1712), .Y(n2479) );
  INVX1 U2306 ( .A(n2479), .Y(n2480) );
  AND2X2 U2307 ( .A(n5094), .B(n1712), .Y(n2481) );
  INVX1 U2308 ( .A(n2481), .Y(n2482) );
  AND2X2 U2309 ( .A(n5098), .B(n1712), .Y(n2483) );
  INVX1 U2310 ( .A(n2483), .Y(n2484) );
  AND2X2 U2311 ( .A(n5102), .B(n1712), .Y(n2485) );
  INVX1 U2312 ( .A(n2485), .Y(n2486) );
  AND2X2 U2313 ( .A(n5108), .B(n1712), .Y(n2487) );
  INVX1 U2314 ( .A(n2487), .Y(n2488) );
  AND2X2 U2315 ( .A(n5072), .B(n1717), .Y(n2489) );
  INVX1 U2316 ( .A(n2489), .Y(n2490) );
  AND2X2 U2317 ( .A(n5077), .B(n1717), .Y(n2491) );
  INVX1 U2318 ( .A(n2491), .Y(n2492) );
  AND2X2 U2319 ( .A(n5082), .B(n1717), .Y(n2493) );
  INVX1 U2320 ( .A(n2493), .Y(n2494) );
  AND2X2 U2321 ( .A(n5089), .B(n1717), .Y(n2495) );
  INVX1 U2322 ( .A(n2495), .Y(n2496) );
  AND2X2 U2323 ( .A(n5094), .B(n1717), .Y(n2497) );
  INVX1 U2324 ( .A(n2497), .Y(n2498) );
  AND2X2 U2325 ( .A(n5098), .B(n1717), .Y(n2499) );
  INVX1 U2326 ( .A(n2499), .Y(n2500) );
  AND2X2 U2327 ( .A(n5102), .B(n1717), .Y(n2501) );
  INVX1 U2328 ( .A(n2501), .Y(n2502) );
  AND2X2 U2329 ( .A(n5108), .B(n1717), .Y(n2503) );
  INVX1 U2330 ( .A(n2503), .Y(n2504) );
  AND2X2 U2331 ( .A(n5072), .B(n1719), .Y(n2505) );
  INVX1 U2332 ( .A(n2505), .Y(n2506) );
  AND2X2 U2333 ( .A(n5077), .B(n1719), .Y(n2507) );
  INVX1 U2334 ( .A(n2507), .Y(n2508) );
  AND2X2 U2335 ( .A(n5082), .B(n1719), .Y(n2509) );
  INVX1 U2336 ( .A(n2509), .Y(n2510) );
  AND2X2 U2337 ( .A(n5089), .B(n1719), .Y(n2511) );
  INVX1 U2338 ( .A(n2511), .Y(n2512) );
  AND2X2 U2339 ( .A(n5094), .B(n1719), .Y(n2513) );
  INVX1 U2340 ( .A(n2513), .Y(n2514) );
  AND2X2 U2341 ( .A(n5098), .B(n1719), .Y(n2515) );
  INVX1 U2342 ( .A(n2515), .Y(n2516) );
  AND2X2 U2343 ( .A(n5102), .B(n1719), .Y(n2517) );
  INVX1 U2344 ( .A(n2517), .Y(n2518) );
  AND2X2 U2345 ( .A(n5108), .B(n1719), .Y(n2519) );
  INVX1 U2346 ( .A(n2519), .Y(n2520) );
  AND2X2 U2347 ( .A(n5072), .B(n1721), .Y(n2521) );
  INVX1 U2348 ( .A(n2521), .Y(n2522) );
  AND2X2 U2349 ( .A(n5077), .B(n1721), .Y(n2523) );
  INVX1 U2350 ( .A(n2523), .Y(n2524) );
  AND2X2 U2351 ( .A(n5082), .B(n1721), .Y(n2525) );
  INVX1 U2352 ( .A(n2525), .Y(n2526) );
  AND2X2 U2353 ( .A(n5089), .B(n1721), .Y(n2527) );
  INVX1 U2354 ( .A(n2527), .Y(n2528) );
  AND2X2 U2355 ( .A(n5094), .B(n1721), .Y(n2529) );
  INVX1 U2356 ( .A(n2529), .Y(n2530) );
  AND2X2 U2357 ( .A(n5098), .B(n1721), .Y(n2531) );
  INVX1 U2358 ( .A(n2531), .Y(n2532) );
  AND2X2 U2359 ( .A(n5102), .B(n1721), .Y(n2533) );
  INVX1 U2360 ( .A(n2533), .Y(n2534) );
  AND2X2 U2361 ( .A(n5108), .B(n1721), .Y(n2535) );
  INVX1 U2362 ( .A(n2535), .Y(n2536) );
  AND2X2 U2363 ( .A(n5072), .B(n1723), .Y(n2537) );
  INVX1 U2364 ( .A(n2537), .Y(n2538) );
  AND2X2 U2365 ( .A(n5077), .B(n1723), .Y(n2539) );
  INVX1 U2366 ( .A(n2539), .Y(n2540) );
  AND2X2 U2367 ( .A(n5082), .B(n1723), .Y(n2541) );
  INVX1 U2368 ( .A(n2541), .Y(n2542) );
  AND2X2 U2369 ( .A(n5089), .B(n1723), .Y(n2543) );
  INVX1 U2370 ( .A(n2543), .Y(n2544) );
  AND2X2 U2371 ( .A(n5094), .B(n1723), .Y(n2545) );
  INVX1 U2372 ( .A(n2545), .Y(n2546) );
  AND2X2 U2373 ( .A(n5098), .B(n1723), .Y(n2547) );
  INVX1 U2374 ( .A(n2547), .Y(n2548) );
  AND2X2 U2375 ( .A(n5102), .B(n1723), .Y(n2549) );
  INVX1 U2376 ( .A(n2549), .Y(n2550) );
  AND2X2 U2377 ( .A(n5108), .B(n1723), .Y(n2551) );
  INVX1 U2378 ( .A(n2551), .Y(n2552) );
  AND2X2 U2379 ( .A(n5072), .B(n1725), .Y(n2553) );
  INVX1 U2380 ( .A(n2553), .Y(n2554) );
  AND2X2 U2381 ( .A(n5077), .B(n1725), .Y(n2555) );
  INVX1 U2382 ( .A(n2555), .Y(n2556) );
  AND2X2 U2383 ( .A(n5082), .B(n1725), .Y(n2557) );
  INVX1 U2384 ( .A(n2557), .Y(n2558) );
  AND2X2 U2385 ( .A(n5089), .B(n1725), .Y(n2559) );
  INVX1 U2386 ( .A(n2559), .Y(n2560) );
  AND2X2 U2387 ( .A(n5094), .B(n1725), .Y(n2561) );
  INVX1 U2388 ( .A(n2561), .Y(n2562) );
  AND2X2 U2389 ( .A(n5098), .B(n1725), .Y(n2563) );
  INVX1 U2390 ( .A(n2563), .Y(n2564) );
  AND2X2 U2391 ( .A(n5102), .B(n1725), .Y(n2565) );
  INVX1 U2392 ( .A(n2565), .Y(n2566) );
  AND2X2 U2393 ( .A(n5108), .B(n1725), .Y(n2567) );
  INVX1 U2394 ( .A(n2567), .Y(n2568) );
  AND2X2 U2395 ( .A(n5072), .B(n1727), .Y(n2569) );
  INVX1 U2396 ( .A(n2569), .Y(n2570) );
  AND2X2 U2397 ( .A(n5077), .B(n1727), .Y(n2571) );
  INVX1 U2398 ( .A(n2571), .Y(n2572) );
  AND2X2 U2399 ( .A(n5082), .B(n1727), .Y(n2573) );
  INVX1 U2400 ( .A(n2573), .Y(n2574) );
  AND2X2 U2401 ( .A(n5089), .B(n1727), .Y(n2575) );
  INVX1 U2402 ( .A(n2575), .Y(n2576) );
  AND2X2 U2403 ( .A(n5094), .B(n1727), .Y(n2577) );
  INVX1 U2404 ( .A(n2577), .Y(n2578) );
  AND2X2 U2405 ( .A(n5098), .B(n1727), .Y(n2579) );
  INVX1 U2406 ( .A(n2579), .Y(n2580) );
  AND2X2 U2407 ( .A(n5102), .B(n1727), .Y(n2581) );
  INVX1 U2408 ( .A(n2581), .Y(n2582) );
  AND2X2 U2409 ( .A(n5108), .B(n1727), .Y(n2583) );
  INVX1 U2410 ( .A(n2583), .Y(n2584) );
  AND2X2 U2411 ( .A(n5072), .B(n1729), .Y(n2585) );
  INVX1 U2412 ( .A(n2585), .Y(n2586) );
  AND2X2 U2413 ( .A(n5077), .B(n1729), .Y(n2587) );
  INVX1 U2414 ( .A(n2587), .Y(n2588) );
  AND2X2 U2415 ( .A(n5082), .B(n1729), .Y(n2589) );
  INVX1 U2416 ( .A(n2589), .Y(n2590) );
  AND2X2 U2417 ( .A(n5089), .B(n1729), .Y(n2591) );
  INVX1 U2418 ( .A(n2591), .Y(n2592) );
  AND2X2 U2419 ( .A(n5094), .B(n1729), .Y(n2593) );
  INVX1 U2420 ( .A(n2593), .Y(n2594) );
  AND2X2 U2421 ( .A(n5098), .B(n1729), .Y(n2595) );
  INVX1 U2422 ( .A(n2595), .Y(n2596) );
  AND2X2 U2423 ( .A(n5102), .B(n1729), .Y(n2597) );
  INVX1 U2424 ( .A(n2597), .Y(n2598) );
  AND2X2 U2425 ( .A(n5108), .B(n1729), .Y(n2599) );
  INVX1 U2426 ( .A(n2599), .Y(n2600) );
  AND2X2 U2427 ( .A(n5072), .B(n1731), .Y(n2601) );
  INVX1 U2428 ( .A(n2601), .Y(n2602) );
  AND2X2 U2429 ( .A(n5077), .B(n1731), .Y(n2603) );
  INVX1 U2430 ( .A(n2603), .Y(n2604) );
  AND2X2 U2431 ( .A(n5082), .B(n1731), .Y(n2605) );
  INVX1 U2432 ( .A(n2605), .Y(n2606) );
  AND2X2 U2433 ( .A(n5089), .B(n1731), .Y(n2607) );
  INVX1 U2434 ( .A(n2607), .Y(n2608) );
  AND2X2 U2435 ( .A(n5094), .B(n1731), .Y(n2609) );
  INVX1 U2436 ( .A(n2609), .Y(n2610) );
  AND2X2 U2437 ( .A(n5098), .B(n1731), .Y(n2611) );
  INVX1 U2438 ( .A(n2611), .Y(n2612) );
  AND2X2 U2439 ( .A(n5102), .B(n1731), .Y(n2613) );
  INVX1 U2440 ( .A(n2613), .Y(n2614) );
  AND2X2 U2441 ( .A(n5108), .B(n1731), .Y(n2615) );
  INVX1 U2442 ( .A(n2615), .Y(n2616) );
  AND2X2 U2443 ( .A(n5073), .B(n1733), .Y(n2617) );
  INVX1 U2444 ( .A(n2617), .Y(n2618) );
  AND2X2 U2445 ( .A(n5078), .B(n1733), .Y(n2619) );
  INVX1 U2446 ( .A(n2619), .Y(n2620) );
  AND2X2 U2447 ( .A(n5082), .B(n1733), .Y(n2621) );
  INVX1 U2448 ( .A(n2621), .Y(n2622) );
  AND2X2 U2449 ( .A(n5087), .B(n1733), .Y(n2623) );
  INVX1 U2450 ( .A(n2623), .Y(n2624) );
  AND2X2 U2451 ( .A(n5095), .B(n1733), .Y(n2625) );
  INVX1 U2452 ( .A(n2625), .Y(n2626) );
  AND2X2 U2453 ( .A(n5099), .B(n1733), .Y(n2627) );
  INVX1 U2454 ( .A(n2627), .Y(n2628) );
  AND2X2 U2455 ( .A(n5103), .B(n1733), .Y(n2629) );
  INVX1 U2456 ( .A(n2629), .Y(n2630) );
  AND2X2 U2457 ( .A(n5107), .B(n1733), .Y(n2631) );
  INVX1 U2458 ( .A(n2631), .Y(n2632) );
  AND2X2 U2459 ( .A(n5073), .B(n1735), .Y(n2633) );
  INVX1 U2460 ( .A(n2633), .Y(n2634) );
  AND2X2 U2461 ( .A(n5078), .B(n1735), .Y(n2635) );
  INVX1 U2462 ( .A(n2635), .Y(n2636) );
  AND2X2 U2463 ( .A(n5082), .B(n1735), .Y(n2637) );
  INVX1 U2464 ( .A(n2637), .Y(n2638) );
  AND2X2 U2465 ( .A(n5087), .B(n1735), .Y(n2639) );
  INVX1 U2466 ( .A(n2639), .Y(n2640) );
  AND2X2 U2467 ( .A(n5095), .B(n1735), .Y(n2641) );
  INVX1 U2468 ( .A(n2641), .Y(n2642) );
  AND2X2 U2469 ( .A(n5099), .B(n1735), .Y(n2643) );
  INVX1 U2470 ( .A(n2643), .Y(n2644) );
  AND2X2 U2471 ( .A(n5103), .B(n1735), .Y(n2645) );
  INVX1 U2472 ( .A(n2645), .Y(n2646) );
  AND2X2 U2473 ( .A(n5107), .B(n1735), .Y(n2647) );
  INVX1 U2474 ( .A(n2647), .Y(n2648) );
  AND2X2 U2475 ( .A(n5073), .B(n1737), .Y(n2649) );
  INVX1 U2476 ( .A(n2649), .Y(n2650) );
  AND2X2 U2477 ( .A(n5078), .B(n1737), .Y(n2651) );
  INVX1 U2478 ( .A(n2651), .Y(n2652) );
  AND2X2 U2479 ( .A(n5082), .B(n1737), .Y(n2653) );
  INVX1 U2480 ( .A(n2653), .Y(n2654) );
  AND2X2 U2481 ( .A(n5087), .B(n1737), .Y(n2655) );
  INVX1 U2482 ( .A(n2655), .Y(n2656) );
  AND2X2 U2483 ( .A(n5095), .B(n1737), .Y(n2657) );
  INVX1 U2484 ( .A(n2657), .Y(n2658) );
  AND2X2 U2485 ( .A(n5099), .B(n1737), .Y(n2659) );
  INVX1 U2486 ( .A(n2659), .Y(n2660) );
  AND2X2 U2487 ( .A(n5103), .B(n1737), .Y(n2661) );
  INVX1 U2488 ( .A(n2661), .Y(n2662) );
  AND2X2 U2489 ( .A(n5107), .B(n1737), .Y(n2663) );
  INVX1 U2490 ( .A(n2663), .Y(n2664) );
  AND2X2 U2491 ( .A(n5073), .B(n1739), .Y(n2665) );
  INVX1 U2492 ( .A(n2665), .Y(n2666) );
  AND2X2 U2493 ( .A(n5078), .B(n1739), .Y(n2667) );
  INVX1 U2494 ( .A(n2667), .Y(n2668) );
  AND2X2 U2495 ( .A(n5082), .B(n1739), .Y(n2669) );
  INVX1 U2496 ( .A(n2669), .Y(n2670) );
  AND2X2 U2497 ( .A(n5087), .B(n1739), .Y(n2671) );
  INVX1 U2498 ( .A(n2671), .Y(n2672) );
  AND2X2 U2499 ( .A(n5095), .B(n1739), .Y(n2673) );
  INVX1 U2500 ( .A(n2673), .Y(n2674) );
  AND2X2 U2501 ( .A(n5099), .B(n1739), .Y(n2675) );
  INVX1 U2502 ( .A(n2675), .Y(n2676) );
  AND2X2 U2503 ( .A(n5103), .B(n1739), .Y(n2677) );
  INVX1 U2504 ( .A(n2677), .Y(n2678) );
  AND2X2 U2505 ( .A(n5107), .B(n1739), .Y(n2679) );
  INVX1 U2506 ( .A(n2679), .Y(n2680) );
  AND2X2 U2507 ( .A(n5073), .B(n1741), .Y(n2681) );
  INVX1 U2508 ( .A(n2681), .Y(n2682) );
  AND2X2 U2509 ( .A(n5078), .B(n1741), .Y(n2683) );
  INVX1 U2510 ( .A(n2683), .Y(n2684) );
  AND2X2 U2511 ( .A(n5082), .B(n1741), .Y(n2685) );
  INVX1 U2512 ( .A(n2685), .Y(n2686) );
  AND2X2 U2513 ( .A(n5087), .B(n1741), .Y(n2687) );
  INVX1 U2514 ( .A(n2687), .Y(n2688) );
  AND2X2 U2515 ( .A(n5095), .B(n1741), .Y(n2689) );
  INVX1 U2516 ( .A(n2689), .Y(n2690) );
  AND2X2 U2517 ( .A(n5099), .B(n1741), .Y(n2691) );
  INVX1 U2518 ( .A(n2691), .Y(n2692) );
  AND2X2 U2519 ( .A(n5103), .B(n1741), .Y(n2693) );
  INVX1 U2520 ( .A(n2693), .Y(n2694) );
  AND2X2 U2521 ( .A(n5107), .B(n1741), .Y(n2695) );
  INVX1 U2522 ( .A(n2695), .Y(n2696) );
  AND2X2 U2523 ( .A(n5073), .B(n1743), .Y(n2697) );
  INVX1 U2524 ( .A(n2697), .Y(n2698) );
  AND2X2 U2525 ( .A(n5078), .B(n1743), .Y(n2699) );
  INVX1 U2526 ( .A(n2699), .Y(n2700) );
  AND2X2 U2527 ( .A(n5082), .B(n1743), .Y(n2701) );
  INVX1 U2528 ( .A(n2701), .Y(n2702) );
  AND2X2 U2529 ( .A(n5087), .B(n1743), .Y(n2703) );
  INVX1 U2530 ( .A(n2703), .Y(n2704) );
  AND2X2 U2531 ( .A(n5095), .B(n1743), .Y(n2705) );
  INVX1 U2532 ( .A(n2705), .Y(n2706) );
  AND2X2 U2533 ( .A(n5099), .B(n1743), .Y(n2707) );
  INVX1 U2534 ( .A(n2707), .Y(n2708) );
  AND2X2 U2535 ( .A(n5103), .B(n1743), .Y(n2709) );
  INVX1 U2536 ( .A(n2709), .Y(n2710) );
  AND2X2 U2537 ( .A(n5107), .B(n1743), .Y(n2711) );
  INVX1 U2538 ( .A(n2711), .Y(n2712) );
  AND2X2 U2539 ( .A(n5073), .B(n1745), .Y(n2713) );
  INVX1 U2540 ( .A(n2713), .Y(n2714) );
  AND2X2 U2541 ( .A(n5078), .B(n1745), .Y(n2715) );
  INVX1 U2542 ( .A(n2715), .Y(n2716) );
  AND2X2 U2543 ( .A(n5082), .B(n1745), .Y(n2717) );
  INVX1 U2544 ( .A(n2717), .Y(n2718) );
  AND2X2 U2545 ( .A(n5087), .B(n1745), .Y(n2719) );
  INVX1 U2546 ( .A(n2719), .Y(n2720) );
  AND2X2 U2547 ( .A(n5095), .B(n1745), .Y(n2721) );
  INVX1 U2548 ( .A(n2721), .Y(n2722) );
  AND2X2 U2549 ( .A(n5099), .B(n1745), .Y(n2723) );
  INVX1 U2550 ( .A(n2723), .Y(n2724) );
  AND2X2 U2551 ( .A(n5103), .B(n1745), .Y(n2725) );
  INVX1 U2552 ( .A(n2725), .Y(n2726) );
  AND2X2 U2553 ( .A(n5107), .B(n1745), .Y(n2727) );
  INVX1 U2554 ( .A(n2727), .Y(n2728) );
  AND2X2 U2555 ( .A(n5073), .B(n1752), .Y(n2729) );
  INVX1 U2556 ( .A(n2729), .Y(n2730) );
  AND2X2 U2557 ( .A(n5078), .B(n1752), .Y(n2731) );
  INVX1 U2558 ( .A(n2731), .Y(n2732) );
  AND2X2 U2559 ( .A(n5082), .B(n1752), .Y(n2733) );
  INVX1 U2560 ( .A(n2733), .Y(n2734) );
  AND2X2 U2561 ( .A(n5087), .B(n1752), .Y(n2735) );
  INVX1 U2562 ( .A(n2735), .Y(n2736) );
  AND2X2 U2563 ( .A(n5095), .B(n1752), .Y(n2737) );
  INVX1 U2564 ( .A(n2737), .Y(n2738) );
  AND2X2 U2565 ( .A(n5099), .B(n1752), .Y(n2739) );
  INVX1 U2566 ( .A(n2739), .Y(n2740) );
  AND2X2 U2567 ( .A(n5103), .B(n1752), .Y(n2741) );
  INVX1 U2568 ( .A(n2741), .Y(n2742) );
  AND2X2 U2569 ( .A(n5107), .B(n1752), .Y(n2743) );
  INVX1 U2570 ( .A(n2743), .Y(n2744) );
  AND2X2 U2571 ( .A(n5072), .B(n1754), .Y(n2745) );
  INVX1 U2572 ( .A(n2745), .Y(n2746) );
  AND2X2 U2573 ( .A(n5078), .B(n1754), .Y(n2747) );
  INVX1 U2574 ( .A(n2747), .Y(n2748) );
  AND2X2 U2575 ( .A(n5083), .B(n1754), .Y(n2749) );
  INVX1 U2576 ( .A(n2749), .Y(n2750) );
  AND2X2 U2577 ( .A(n5088), .B(n1754), .Y(n2751) );
  INVX1 U2578 ( .A(n2751), .Y(n2752) );
  AND2X2 U2579 ( .A(n5095), .B(n1754), .Y(n2753) );
  INVX1 U2580 ( .A(n2753), .Y(n2754) );
  AND2X2 U2581 ( .A(n5099), .B(n1754), .Y(n2755) );
  INVX1 U2582 ( .A(n2755), .Y(n2756) );
  AND2X2 U2583 ( .A(n5103), .B(n1754), .Y(n2757) );
  INVX1 U2584 ( .A(n2757), .Y(n2758) );
  AND2X2 U2585 ( .A(n5108), .B(n1754), .Y(n2759) );
  INVX1 U2586 ( .A(n2759), .Y(n2760) );
  AND2X2 U2587 ( .A(n5072), .B(n1756), .Y(n2761) );
  INVX1 U2588 ( .A(n2761), .Y(n2762) );
  AND2X2 U2589 ( .A(n5078), .B(n1756), .Y(n2763) );
  INVX1 U2590 ( .A(n2763), .Y(n2764) );
  AND2X2 U2591 ( .A(n5083), .B(n1756), .Y(n2765) );
  INVX1 U2592 ( .A(n2765), .Y(n2766) );
  AND2X2 U2593 ( .A(n5088), .B(n1756), .Y(n2767) );
  INVX1 U2594 ( .A(n2767), .Y(n2768) );
  AND2X2 U2595 ( .A(n5095), .B(n1756), .Y(n2769) );
  INVX1 U2596 ( .A(n2769), .Y(n2770) );
  AND2X2 U2597 ( .A(n5099), .B(n1756), .Y(n2771) );
  INVX1 U2598 ( .A(n2771), .Y(n2772) );
  AND2X2 U2599 ( .A(n5103), .B(n1756), .Y(n2773) );
  INVX1 U2600 ( .A(n2773), .Y(n2774) );
  AND2X2 U2601 ( .A(n5108), .B(n1756), .Y(n2775) );
  INVX1 U2602 ( .A(n2775), .Y(n2776) );
  AND2X2 U2603 ( .A(n5074), .B(n1761), .Y(n2777) );
  INVX1 U2604 ( .A(n2777), .Y(n2778) );
  AND2X2 U2605 ( .A(n5078), .B(n1761), .Y(n2779) );
  INVX1 U2606 ( .A(n2779), .Y(n2780) );
  AND2X2 U2607 ( .A(n5083), .B(n1761), .Y(n2781) );
  INVX1 U2608 ( .A(n2781), .Y(n2782) );
  AND2X2 U2609 ( .A(n5088), .B(n1761), .Y(n2783) );
  INVX1 U2610 ( .A(n2783), .Y(n2784) );
  AND2X2 U2611 ( .A(n5095), .B(n1761), .Y(n2785) );
  INVX1 U2612 ( .A(n2785), .Y(n2786) );
  AND2X2 U2613 ( .A(n5099), .B(n1761), .Y(n2787) );
  INVX1 U2614 ( .A(n2787), .Y(n2788) );
  AND2X2 U2615 ( .A(n5103), .B(n1761), .Y(n2789) );
  INVX1 U2616 ( .A(n2789), .Y(n2790) );
  AND2X2 U2617 ( .A(n5108), .B(n1761), .Y(n2791) );
  INVX1 U2618 ( .A(n2791), .Y(n2792) );
  AND2X2 U2619 ( .A(n5074), .B(n1763), .Y(n2793) );
  INVX1 U2620 ( .A(n2793), .Y(n2794) );
  AND2X2 U2621 ( .A(n5078), .B(n1763), .Y(n2795) );
  INVX1 U2622 ( .A(n2795), .Y(n2796) );
  AND2X2 U2623 ( .A(n5083), .B(n1763), .Y(n2797) );
  INVX1 U2624 ( .A(n2797), .Y(n2798) );
  AND2X2 U2625 ( .A(n5088), .B(n1763), .Y(n2799) );
  INVX1 U2626 ( .A(n2799), .Y(n2800) );
  AND2X2 U2627 ( .A(n5095), .B(n1763), .Y(n2801) );
  INVX1 U2628 ( .A(n2801), .Y(n2802) );
  AND2X2 U2629 ( .A(n5099), .B(n1763), .Y(n2803) );
  INVX1 U2630 ( .A(n2803), .Y(n2804) );
  AND2X2 U2631 ( .A(n5103), .B(n1763), .Y(n2805) );
  INVX1 U2632 ( .A(n2805), .Y(n2806) );
  AND2X2 U2633 ( .A(n5108), .B(n1763), .Y(n2807) );
  INVX1 U2634 ( .A(n2807), .Y(n2808) );
  AND2X2 U2635 ( .A(n5072), .B(n1765), .Y(n2809) );
  INVX1 U2636 ( .A(n2809), .Y(n2810) );
  AND2X2 U2637 ( .A(n5078), .B(n1765), .Y(n2811) );
  INVX1 U2638 ( .A(n2811), .Y(n2812) );
  AND2X2 U2639 ( .A(n5083), .B(n1765), .Y(n2813) );
  INVX1 U2640 ( .A(n2813), .Y(n2814) );
  AND2X2 U2641 ( .A(n5088), .B(n1765), .Y(n2815) );
  INVX1 U2642 ( .A(n2815), .Y(n2816) );
  AND2X2 U2643 ( .A(n5095), .B(n1765), .Y(n2817) );
  INVX1 U2644 ( .A(n2817), .Y(n2818) );
  AND2X2 U2645 ( .A(n5099), .B(n1765), .Y(n2819) );
  INVX1 U2646 ( .A(n2819), .Y(n2820) );
  AND2X2 U2647 ( .A(n5103), .B(n1765), .Y(n2821) );
  INVX1 U2648 ( .A(n2821), .Y(n2822) );
  AND2X2 U2649 ( .A(n5108), .B(n1765), .Y(n2823) );
  INVX1 U2650 ( .A(n2823), .Y(n2824) );
  AND2X2 U2651 ( .A(n5072), .B(n1767), .Y(n2825) );
  INVX1 U2652 ( .A(n2825), .Y(n2826) );
  AND2X2 U2653 ( .A(n5078), .B(n1767), .Y(n2827) );
  INVX1 U2654 ( .A(n2827), .Y(n2828) );
  AND2X2 U2655 ( .A(n5083), .B(n1767), .Y(n2829) );
  INVX1 U2656 ( .A(n2829), .Y(n2830) );
  AND2X2 U2657 ( .A(n5088), .B(n1767), .Y(n2831) );
  INVX1 U2658 ( .A(n2831), .Y(n2832) );
  AND2X2 U2659 ( .A(n5095), .B(n1767), .Y(n2833) );
  INVX1 U2660 ( .A(n2833), .Y(n2834) );
  AND2X2 U2661 ( .A(n5099), .B(n1767), .Y(n2835) );
  INVX1 U2662 ( .A(n2835), .Y(n2836) );
  AND2X2 U2663 ( .A(n5103), .B(n1767), .Y(n2837) );
  INVX1 U2664 ( .A(n2837), .Y(n2838) );
  AND2X2 U2665 ( .A(n5108), .B(n1767), .Y(n2839) );
  INVX1 U2666 ( .A(n2839), .Y(n2840) );
  AND2X2 U2667 ( .A(n5072), .B(n1769), .Y(n2841) );
  INVX1 U2668 ( .A(n2841), .Y(n2842) );
  AND2X2 U2669 ( .A(n5078), .B(n1769), .Y(n2843) );
  INVX1 U2670 ( .A(n2843), .Y(n2844) );
  AND2X2 U2671 ( .A(n5083), .B(n1769), .Y(n2845) );
  INVX1 U2672 ( .A(n2845), .Y(n2846) );
  AND2X2 U2673 ( .A(n5088), .B(n1769), .Y(n2847) );
  INVX1 U2674 ( .A(n2847), .Y(n2848) );
  AND2X2 U2675 ( .A(n5095), .B(n1769), .Y(n2849) );
  INVX1 U2676 ( .A(n2849), .Y(n2850) );
  AND2X2 U2677 ( .A(n5099), .B(n1769), .Y(n2851) );
  INVX1 U2678 ( .A(n2851), .Y(n2852) );
  AND2X2 U2679 ( .A(n5103), .B(n1769), .Y(n2853) );
  INVX1 U2680 ( .A(n2853), .Y(n2854) );
  AND2X2 U2681 ( .A(n5108), .B(n1769), .Y(n2855) );
  INVX1 U2682 ( .A(n2855), .Y(n2856) );
  AND2X2 U2683 ( .A(n5074), .B(n1771), .Y(n2857) );
  INVX1 U2684 ( .A(n2857), .Y(n2858) );
  AND2X2 U2685 ( .A(n5078), .B(n1771), .Y(n2859) );
  INVX1 U2686 ( .A(n2859), .Y(n2860) );
  AND2X2 U2687 ( .A(n5083), .B(n1771), .Y(n2861) );
  INVX1 U2688 ( .A(n2861), .Y(n2862) );
  AND2X2 U2689 ( .A(n5088), .B(n1771), .Y(n2863) );
  INVX1 U2690 ( .A(n2863), .Y(n2864) );
  AND2X2 U2691 ( .A(n5095), .B(n1771), .Y(n2865) );
  INVX1 U2692 ( .A(n2865), .Y(n2866) );
  AND2X2 U2693 ( .A(n5099), .B(n1771), .Y(n2867) );
  INVX1 U2694 ( .A(n2867), .Y(n2868) );
  AND2X2 U2695 ( .A(n5103), .B(n1771), .Y(n2869) );
  INVX1 U2696 ( .A(n2869), .Y(n2870) );
  AND2X2 U2697 ( .A(n5108), .B(n1771), .Y(n2871) );
  INVX1 U2698 ( .A(n2871), .Y(n2872) );
  AND2X2 U2699 ( .A(n5074), .B(n1776), .Y(n2873) );
  INVX1 U2700 ( .A(n2873), .Y(n2874) );
  AND2X2 U2701 ( .A(n5078), .B(n1776), .Y(n2875) );
  INVX1 U2702 ( .A(n2875), .Y(n2876) );
  AND2X2 U2703 ( .A(n5084), .B(n1776), .Y(n2877) );
  INVX1 U2704 ( .A(n2877), .Y(n2878) );
  AND2X2 U2705 ( .A(n5089), .B(n1776), .Y(n2879) );
  INVX1 U2706 ( .A(n2879), .Y(n2880) );
  AND2X2 U2707 ( .A(n5095), .B(n1776), .Y(n2881) );
  INVX1 U2708 ( .A(n2881), .Y(n2882) );
  AND2X2 U2709 ( .A(n5099), .B(n1776), .Y(n2883) );
  INVX1 U2710 ( .A(n2883), .Y(n2884) );
  AND2X2 U2711 ( .A(n5103), .B(n1776), .Y(n2885) );
  INVX1 U2712 ( .A(n2885), .Y(n2886) );
  AND2X2 U2713 ( .A(n5108), .B(n1776), .Y(n2887) );
  INVX1 U2714 ( .A(n2887), .Y(n2888) );
  AND2X2 U2715 ( .A(n5074), .B(n1778), .Y(n2889) );
  INVX1 U2716 ( .A(n2889), .Y(n2890) );
  AND2X2 U2717 ( .A(n5078), .B(n1778), .Y(n2891) );
  INVX1 U2718 ( .A(n2891), .Y(n2892) );
  AND2X2 U2719 ( .A(n5084), .B(n1778), .Y(n2893) );
  INVX1 U2720 ( .A(n2893), .Y(n2894) );
  AND2X2 U2721 ( .A(n5089), .B(n1778), .Y(n2895) );
  INVX1 U2722 ( .A(n2895), .Y(n2896) );
  AND2X2 U2723 ( .A(n5095), .B(n1778), .Y(n2897) );
  INVX1 U2724 ( .A(n2897), .Y(n2898) );
  AND2X2 U2725 ( .A(n5099), .B(n1778), .Y(n2899) );
  INVX1 U2726 ( .A(n2899), .Y(n2900) );
  AND2X2 U2727 ( .A(n5103), .B(n1778), .Y(n2901) );
  INVX1 U2728 ( .A(n2901), .Y(n2902) );
  AND2X2 U2729 ( .A(n5108), .B(n1778), .Y(n2903) );
  INVX1 U2730 ( .A(n2903), .Y(n2904) );
  AND2X2 U2731 ( .A(n5074), .B(n1780), .Y(n2905) );
  INVX1 U2732 ( .A(n2905), .Y(n2906) );
  AND2X2 U2733 ( .A(n5078), .B(n1780), .Y(n2907) );
  INVX1 U2734 ( .A(n2907), .Y(n2908) );
  AND2X2 U2735 ( .A(n5084), .B(n1780), .Y(n2909) );
  INVX1 U2736 ( .A(n2909), .Y(n2910) );
  AND2X2 U2737 ( .A(n5089), .B(n1780), .Y(n2911) );
  INVX1 U2738 ( .A(n2911), .Y(n2912) );
  AND2X2 U2739 ( .A(n5095), .B(n1780), .Y(n2913) );
  INVX1 U2740 ( .A(n2913), .Y(n2914) );
  AND2X2 U2741 ( .A(n5099), .B(n1780), .Y(n2915) );
  INVX1 U2742 ( .A(n2915), .Y(n2916) );
  AND2X2 U2743 ( .A(n5103), .B(n1780), .Y(n2917) );
  INVX1 U2744 ( .A(n2917), .Y(n2918) );
  AND2X2 U2745 ( .A(n5108), .B(n1780), .Y(n2919) );
  INVX1 U2746 ( .A(n2919), .Y(n2920) );
  AND2X2 U2747 ( .A(n5074), .B(n1782), .Y(n2921) );
  INVX1 U2748 ( .A(n2921), .Y(n2922) );
  AND2X2 U2749 ( .A(n5078), .B(n1782), .Y(n2923) );
  INVX1 U2750 ( .A(n2923), .Y(n2924) );
  AND2X2 U2751 ( .A(n5084), .B(n1782), .Y(n2925) );
  INVX1 U2752 ( .A(n2925), .Y(n2926) );
  AND2X2 U2753 ( .A(n5089), .B(n1782), .Y(n2927) );
  INVX1 U2754 ( .A(n2927), .Y(n2928) );
  AND2X2 U2755 ( .A(n5095), .B(n1782), .Y(n2929) );
  INVX1 U2756 ( .A(n2929), .Y(n2930) );
  AND2X2 U2757 ( .A(n5099), .B(n1782), .Y(n2931) );
  INVX1 U2758 ( .A(n2931), .Y(n2932) );
  AND2X2 U2759 ( .A(n5103), .B(n1782), .Y(n2933) );
  INVX1 U2760 ( .A(n2933), .Y(n2934) );
  AND2X2 U2761 ( .A(n5108), .B(n1782), .Y(n2935) );
  INVX1 U2762 ( .A(n2935), .Y(n2936) );
  AND2X2 U2763 ( .A(n5074), .B(n1784), .Y(n2937) );
  INVX1 U2764 ( .A(n2937), .Y(n2938) );
  AND2X2 U2765 ( .A(n5078), .B(n1784), .Y(n2939) );
  INVX1 U2766 ( .A(n2939), .Y(n2940) );
  AND2X2 U2767 ( .A(n5084), .B(n1784), .Y(n2941) );
  INVX1 U2768 ( .A(n2941), .Y(n2942) );
  AND2X2 U2769 ( .A(n5089), .B(n1784), .Y(n2943) );
  INVX1 U2770 ( .A(n2943), .Y(n2944) );
  AND2X2 U2771 ( .A(n5095), .B(n1784), .Y(n2945) );
  INVX1 U2772 ( .A(n2945), .Y(n2946) );
  AND2X2 U2773 ( .A(n5099), .B(n1784), .Y(n2947) );
  INVX1 U2774 ( .A(n2947), .Y(n2948) );
  AND2X2 U2775 ( .A(n5103), .B(n1784), .Y(n2949) );
  INVX1 U2776 ( .A(n2949), .Y(n2950) );
  AND2X2 U2777 ( .A(n5108), .B(n1784), .Y(n2951) );
  INVX1 U2778 ( .A(n2951), .Y(n2952) );
  AND2X2 U2779 ( .A(n5074), .B(n1786), .Y(n2953) );
  INVX1 U2780 ( .A(n2953), .Y(n2954) );
  AND2X2 U2781 ( .A(n5078), .B(n1786), .Y(n2955) );
  INVX1 U2782 ( .A(n2955), .Y(n2956) );
  AND2X2 U2783 ( .A(n5084), .B(n1786), .Y(n2957) );
  INVX1 U2784 ( .A(n2957), .Y(n2958) );
  AND2X2 U2785 ( .A(n5089), .B(n1786), .Y(n2959) );
  INVX1 U2786 ( .A(n2959), .Y(n2960) );
  AND2X2 U2787 ( .A(n5095), .B(n1786), .Y(n2961) );
  INVX1 U2788 ( .A(n2961), .Y(n2962) );
  AND2X2 U2789 ( .A(n5099), .B(n1786), .Y(n2963) );
  INVX1 U2790 ( .A(n2963), .Y(n2964) );
  AND2X2 U2791 ( .A(n5103), .B(n1786), .Y(n2965) );
  INVX1 U2792 ( .A(n2965), .Y(n2966) );
  AND2X2 U2793 ( .A(n5108), .B(n1786), .Y(n2967) );
  INVX1 U2794 ( .A(n2967), .Y(n2968) );
  AND2X2 U2795 ( .A(n5074), .B(n1788), .Y(n2969) );
  INVX1 U2796 ( .A(n2969), .Y(n2970) );
  AND2X2 U2797 ( .A(n5078), .B(n1788), .Y(n2971) );
  INVX1 U2798 ( .A(n2971), .Y(n2972) );
  AND2X2 U2799 ( .A(n5084), .B(n1788), .Y(n2973) );
  INVX1 U2800 ( .A(n2973), .Y(n2974) );
  AND2X2 U2801 ( .A(n5089), .B(n1788), .Y(n2975) );
  INVX1 U2802 ( .A(n2975), .Y(n2976) );
  AND2X2 U2803 ( .A(n5095), .B(n1788), .Y(n2977) );
  INVX1 U2804 ( .A(n2977), .Y(n2978) );
  AND2X2 U2805 ( .A(n5099), .B(n1788), .Y(n2979) );
  INVX1 U2806 ( .A(n2979), .Y(n2980) );
  AND2X2 U2807 ( .A(n5103), .B(n1788), .Y(n2981) );
  INVX1 U2808 ( .A(n2981), .Y(n2982) );
  AND2X2 U2809 ( .A(n5108), .B(n1788), .Y(n2983) );
  INVX1 U2810 ( .A(n2983), .Y(n2984) );
  AND2X2 U2811 ( .A(n5074), .B(n1790), .Y(n2985) );
  INVX1 U2812 ( .A(n2985), .Y(n2986) );
  AND2X2 U2813 ( .A(n5078), .B(n1790), .Y(n2987) );
  INVX1 U2814 ( .A(n2987), .Y(n2988) );
  AND2X2 U2815 ( .A(n5084), .B(n1790), .Y(n2989) );
  INVX1 U2816 ( .A(n2989), .Y(n2990) );
  AND2X2 U2817 ( .A(n5089), .B(n1790), .Y(n2991) );
  INVX1 U2818 ( .A(n2991), .Y(n2992) );
  AND2X2 U2819 ( .A(n5095), .B(n1790), .Y(n2993) );
  INVX1 U2820 ( .A(n2993), .Y(n2994) );
  AND2X2 U2821 ( .A(n5099), .B(n1790), .Y(n2995) );
  INVX1 U2822 ( .A(n2995), .Y(n2996) );
  AND2X2 U2823 ( .A(n5103), .B(n1790), .Y(n2997) );
  INVX1 U2824 ( .A(n2997), .Y(n2998) );
  AND2X2 U2825 ( .A(n5074), .B(n1792), .Y(n2999) );
  INVX1 U2826 ( .A(n2999), .Y(n3000) );
  AND2X2 U2827 ( .A(n5078), .B(n1792), .Y(n3001) );
  INVX1 U2828 ( .A(n3001), .Y(n3002) );
  AND2X2 U2829 ( .A(n5084), .B(n1792), .Y(n3003) );
  INVX1 U2830 ( .A(n3003), .Y(n3004) );
  AND2X2 U2831 ( .A(n5089), .B(n1792), .Y(n3005) );
  INVX1 U2832 ( .A(n3005), .Y(n3006) );
  AND2X2 U2833 ( .A(n5095), .B(n1792), .Y(n3007) );
  INVX1 U2834 ( .A(n3007), .Y(n3008) );
  AND2X2 U2835 ( .A(n5099), .B(n1792), .Y(n3009) );
  INVX1 U2836 ( .A(n3009), .Y(n3010) );
  AND2X2 U2837 ( .A(n5103), .B(n1792), .Y(n3011) );
  INVX1 U2838 ( .A(n3011), .Y(n3012) );
  AND2X2 U2839 ( .A(n5108), .B(n1792), .Y(n3013) );
  INVX1 U2840 ( .A(n3013), .Y(n3014) );
  AND2X2 U2841 ( .A(n5074), .B(n1794), .Y(n3015) );
  INVX1 U2842 ( .A(n3015), .Y(n3016) );
  AND2X2 U2843 ( .A(n5078), .B(n1794), .Y(n3017) );
  INVX1 U2844 ( .A(n3017), .Y(n3018) );
  AND2X2 U2845 ( .A(n5084), .B(n1794), .Y(n3019) );
  INVX1 U2846 ( .A(n3019), .Y(n3020) );
  AND2X2 U2847 ( .A(n5089), .B(n1794), .Y(n3021) );
  INVX1 U2848 ( .A(n3021), .Y(n3022) );
  AND2X2 U2849 ( .A(n5095), .B(n1794), .Y(n3023) );
  INVX1 U2850 ( .A(n3023), .Y(n3024) );
  AND2X2 U2851 ( .A(n5099), .B(n1794), .Y(n3025) );
  INVX1 U2852 ( .A(n3025), .Y(n3026) );
  AND2X2 U2853 ( .A(n5103), .B(n1794), .Y(n3027) );
  INVX1 U2854 ( .A(n3027), .Y(n3028) );
  AND2X2 U2855 ( .A(n5108), .B(n1794), .Y(n3029) );
  INVX1 U2856 ( .A(n3029), .Y(n3030) );
  AND2X2 U2857 ( .A(n5074), .B(n1796), .Y(n3031) );
  INVX1 U2858 ( .A(n3031), .Y(n3032) );
  AND2X2 U2859 ( .A(n5078), .B(n1796), .Y(n3033) );
  INVX1 U2860 ( .A(n3033), .Y(n3034) );
  AND2X2 U2861 ( .A(n5084), .B(n1796), .Y(n3035) );
  INVX1 U2862 ( .A(n3035), .Y(n3036) );
  AND2X2 U2863 ( .A(n5089), .B(n1796), .Y(n3037) );
  INVX1 U2864 ( .A(n3037), .Y(n3038) );
  AND2X2 U2865 ( .A(n5095), .B(n1796), .Y(n3039) );
  INVX1 U2866 ( .A(n3039), .Y(n3040) );
  AND2X2 U2867 ( .A(n5099), .B(n1796), .Y(n3041) );
  INVX1 U2868 ( .A(n3041), .Y(n3042) );
  AND2X2 U2869 ( .A(n5103), .B(n1796), .Y(n3043) );
  INVX1 U2870 ( .A(n3043), .Y(n3044) );
  AND2X2 U2871 ( .A(n5108), .B(n1796), .Y(n3045) );
  INVX1 U2872 ( .A(n3045), .Y(n3046) );
  AND2X2 U2873 ( .A(n5074), .B(n1798), .Y(n3047) );
  INVX1 U2874 ( .A(n3047), .Y(n3048) );
  AND2X2 U2875 ( .A(n5078), .B(n1798), .Y(n3049) );
  INVX1 U2876 ( .A(n3049), .Y(n3050) );
  AND2X2 U2877 ( .A(n5084), .B(n1798), .Y(n3051) );
  INVX1 U2878 ( .A(n3051), .Y(n3052) );
  AND2X2 U2879 ( .A(n5089), .B(n1798), .Y(n3053) );
  INVX1 U2880 ( .A(n3053), .Y(n3054) );
  AND2X2 U2881 ( .A(n5095), .B(n1798), .Y(n3055) );
  INVX1 U2882 ( .A(n3055), .Y(n3056) );
  AND2X2 U2883 ( .A(n5099), .B(n1798), .Y(n3057) );
  INVX1 U2884 ( .A(n3057), .Y(n3058) );
  AND2X2 U2885 ( .A(n5103), .B(n1798), .Y(n3059) );
  INVX1 U2886 ( .A(n3059), .Y(n3060) );
  AND2X2 U2887 ( .A(n5108), .B(n1798), .Y(n3061) );
  INVX1 U2888 ( .A(n3061), .Y(n3062) );
  AND2X2 U2889 ( .A(n5075), .B(n1800), .Y(n3063) );
  INVX1 U2890 ( .A(n3063), .Y(n3064) );
  AND2X2 U2891 ( .A(n5079), .B(n1800), .Y(n3065) );
  INVX1 U2892 ( .A(n3065), .Y(n3066) );
  AND2X2 U2893 ( .A(n5085), .B(n1800), .Y(n3067) );
  INVX1 U2894 ( .A(n3067), .Y(n3068) );
  AND2X2 U2895 ( .A(n5090), .B(n1800), .Y(n3069) );
  INVX1 U2896 ( .A(n3069), .Y(n3070) );
  AND2X2 U2897 ( .A(n5096), .B(n1800), .Y(n3071) );
  INVX1 U2898 ( .A(n3071), .Y(n3072) );
  AND2X2 U2899 ( .A(n5100), .B(n1800), .Y(n3073) );
  INVX1 U2900 ( .A(n3073), .Y(n3074) );
  AND2X2 U2901 ( .A(n5104), .B(n1800), .Y(n3075) );
  INVX1 U2902 ( .A(n3075), .Y(n3076) );
  AND2X2 U2903 ( .A(n5109), .B(n1800), .Y(n3077) );
  INVX1 U2904 ( .A(n3077), .Y(n3078) );
  AND2X2 U2905 ( .A(n5075), .B(n1802), .Y(n3079) );
  INVX1 U2906 ( .A(n3079), .Y(n3080) );
  AND2X2 U2907 ( .A(n5079), .B(n1802), .Y(n3081) );
  INVX1 U2908 ( .A(n3081), .Y(n3082) );
  AND2X2 U2909 ( .A(n5085), .B(n1802), .Y(n3083) );
  INVX1 U2910 ( .A(n3083), .Y(n3084) );
  AND2X2 U2911 ( .A(n5090), .B(n1802), .Y(n3085) );
  INVX1 U2912 ( .A(n3085), .Y(n3086) );
  AND2X2 U2913 ( .A(n5096), .B(n1802), .Y(n3087) );
  INVX1 U2914 ( .A(n3087), .Y(n3088) );
  AND2X2 U2915 ( .A(n5100), .B(n1802), .Y(n3089) );
  INVX1 U2916 ( .A(n3089), .Y(n3090) );
  AND2X2 U2917 ( .A(n5104), .B(n1802), .Y(n3091) );
  INVX1 U2918 ( .A(n3091), .Y(n3092) );
  AND2X2 U2919 ( .A(n5109), .B(n1802), .Y(n3093) );
  INVX1 U2920 ( .A(n3093), .Y(n3094) );
  BUFX2 U2921 ( .A(n5184), .Y(n3095) );
  BUFX2 U2922 ( .A(n5288), .Y(n3096) );
  AND2X2 U2923 ( .A(\mem<22><1> ), .B(n4957), .Y(n3097) );
  INVX1 U2924 ( .A(n3097), .Y(n3098) );
  AND2X2 U2925 ( .A(\mem<63><2> ), .B(n4692), .Y(n3099) );
  INVX1 U2926 ( .A(n3099), .Y(n3100) );
  AND2X2 U2927 ( .A(\mem<63><5> ), .B(n4693), .Y(n3101) );
  INVX1 U2928 ( .A(n3101), .Y(n3102) );
  AND2X2 U2929 ( .A(n5039), .B(n1690), .Y(n3103) );
  INVX1 U2930 ( .A(n3103), .Y(n3104) );
  AND2X2 U2931 ( .A(n5044), .B(n1690), .Y(n3105) );
  INVX1 U2932 ( .A(n3105), .Y(n3106) );
  AND2X2 U2933 ( .A(\data_in<2> ), .B(n1690), .Y(n3107) );
  INVX1 U2934 ( .A(n3107), .Y(n3108) );
  AND2X2 U2935 ( .A(n5052), .B(n1690), .Y(n3109) );
  INVX1 U2936 ( .A(n3109), .Y(n3110) );
  AND2X2 U2937 ( .A(n5057), .B(n1690), .Y(n3111) );
  INVX1 U2938 ( .A(n3111), .Y(n3112) );
  AND2X2 U2939 ( .A(n5061), .B(n1690), .Y(n3113) );
  INVX1 U2940 ( .A(n3113), .Y(n3114) );
  AND2X2 U2941 ( .A(n5066), .B(n1690), .Y(n3115) );
  INVX1 U2942 ( .A(n3115), .Y(n3116) );
  AND2X2 U2943 ( .A(n5070), .B(n1690), .Y(n3117) );
  INVX1 U2944 ( .A(n3117), .Y(n3118) );
  AND2X2 U2945 ( .A(n5039), .B(n1696), .Y(n3119) );
  INVX1 U2946 ( .A(n3119), .Y(n3120) );
  AND2X2 U2947 ( .A(n5045), .B(n1696), .Y(n3121) );
  INVX1 U2948 ( .A(n3121), .Y(n3122) );
  AND2X2 U2949 ( .A(n5048), .B(n1696), .Y(n3123) );
  INVX1 U2950 ( .A(n3123), .Y(n3124) );
  AND2X2 U2951 ( .A(n5052), .B(n1696), .Y(n3125) );
  INVX1 U2952 ( .A(n3125), .Y(n3126) );
  AND2X2 U2953 ( .A(n5057), .B(n1696), .Y(n3127) );
  INVX1 U2954 ( .A(n3127), .Y(n3128) );
  AND2X2 U2955 ( .A(n5061), .B(n1696), .Y(n3129) );
  INVX1 U2956 ( .A(n3129), .Y(n3130) );
  AND2X2 U2957 ( .A(n5066), .B(n1696), .Y(n3131) );
  INVX1 U2958 ( .A(n3131), .Y(n3132) );
  AND2X2 U2959 ( .A(n5070), .B(n1696), .Y(n3133) );
  INVX1 U2960 ( .A(n3133), .Y(n3134) );
  AND2X2 U2961 ( .A(\mem<57><0> ), .B(n3580), .Y(n3135) );
  INVX1 U2962 ( .A(n3135), .Y(n3136) );
  AND2X2 U2963 ( .A(\mem<57><1> ), .B(n3580), .Y(n3137) );
  INVX1 U2964 ( .A(n3137), .Y(n3138) );
  AND2X2 U2965 ( .A(\mem<57><2> ), .B(n3580), .Y(n3139) );
  INVX1 U2966 ( .A(n3139), .Y(n3140) );
  AND2X2 U2967 ( .A(\mem<57><3> ), .B(n3580), .Y(n3141) );
  INVX1 U2968 ( .A(n3141), .Y(n3142) );
  AND2X2 U2969 ( .A(\mem<57><4> ), .B(n3580), .Y(n3143) );
  INVX1 U2970 ( .A(n3143), .Y(n3144) );
  AND2X2 U2971 ( .A(\mem<57><5> ), .B(n3580), .Y(n3145) );
  INVX1 U2972 ( .A(n3145), .Y(n3146) );
  AND2X2 U2973 ( .A(\mem<57><6> ), .B(n3580), .Y(n3147) );
  INVX1 U2974 ( .A(n3147), .Y(n3148) );
  AND2X2 U2975 ( .A(n5039), .B(n1704), .Y(n3149) );
  INVX1 U2976 ( .A(n3149), .Y(n3150) );
  AND2X2 U2977 ( .A(n5045), .B(n1704), .Y(n3151) );
  INVX1 U2978 ( .A(n3151), .Y(n3152) );
  AND2X2 U2979 ( .A(n5047), .B(n1704), .Y(n3153) );
  INVX1 U2980 ( .A(n3153), .Y(n3154) );
  AND2X2 U2981 ( .A(n5051), .B(n1704), .Y(n3155) );
  INVX1 U2982 ( .A(n3155), .Y(n3156) );
  AND2X2 U2983 ( .A(n5057), .B(n1704), .Y(n3157) );
  INVX1 U2984 ( .A(n3157), .Y(n3158) );
  AND2X2 U2985 ( .A(n5061), .B(n1704), .Y(n3159) );
  INVX1 U2986 ( .A(n3159), .Y(n3160) );
  AND2X2 U2987 ( .A(n5066), .B(n1704), .Y(n3161) );
  INVX1 U2988 ( .A(n3161), .Y(n3162) );
  AND2X2 U2989 ( .A(n5070), .B(n1704), .Y(n3163) );
  INVX1 U2990 ( .A(n3163), .Y(n3164) );
  AND2X2 U2991 ( .A(n5039), .B(n1711), .Y(n3165) );
  INVX1 U2992 ( .A(n3165), .Y(n3166) );
  AND2X2 U2993 ( .A(n5045), .B(n1711), .Y(n3167) );
  INVX1 U2994 ( .A(n3167), .Y(n3168) );
  AND2X2 U2995 ( .A(n5049), .B(n1711), .Y(n3169) );
  INVX1 U2996 ( .A(n3169), .Y(n3170) );
  AND2X2 U2997 ( .A(n5052), .B(n1711), .Y(n3171) );
  INVX1 U2998 ( .A(n3171), .Y(n3172) );
  AND2X2 U2999 ( .A(n5057), .B(n1711), .Y(n3173) );
  INVX1 U3000 ( .A(n3173), .Y(n3174) );
  AND2X2 U3001 ( .A(n5061), .B(n1711), .Y(n3175) );
  INVX1 U3002 ( .A(n3175), .Y(n3176) );
  AND2X2 U3003 ( .A(n5066), .B(n1711), .Y(n3177) );
  INVX1 U3004 ( .A(n3177), .Y(n3178) );
  AND2X2 U3005 ( .A(n5070), .B(n1711), .Y(n3179) );
  INVX1 U3006 ( .A(n3179), .Y(n3180) );
  AND2X2 U3007 ( .A(n5039), .B(n1718), .Y(n3181) );
  INVX1 U3008 ( .A(n3181), .Y(n3182) );
  AND2X2 U3009 ( .A(n5044), .B(n1718), .Y(n3183) );
  INVX1 U3010 ( .A(n3183), .Y(n3184) );
  AND2X2 U3011 ( .A(\data_in<2> ), .B(n1718), .Y(n3185) );
  INVX1 U3012 ( .A(n3185), .Y(n3186) );
  AND2X2 U3013 ( .A(n5052), .B(n1718), .Y(n3187) );
  INVX1 U3014 ( .A(n3187), .Y(n3188) );
  AND2X2 U3015 ( .A(n5057), .B(n1718), .Y(n3189) );
  INVX1 U3016 ( .A(n3189), .Y(n3190) );
  AND2X2 U3017 ( .A(n5061), .B(n1718), .Y(n3191) );
  INVX1 U3018 ( .A(n3191), .Y(n3192) );
  AND2X2 U3019 ( .A(n5066), .B(n1718), .Y(n3193) );
  INVX1 U3020 ( .A(n3193), .Y(n3194) );
  AND2X2 U3021 ( .A(n5070), .B(n1718), .Y(n3195) );
  INVX1 U3022 ( .A(n3195), .Y(n3196) );
  AND2X2 U3023 ( .A(n5039), .B(n1720), .Y(n3197) );
  INVX1 U3024 ( .A(n3197), .Y(n3198) );
  AND2X2 U3025 ( .A(n5044), .B(n1720), .Y(n3199) );
  INVX1 U3026 ( .A(n3199), .Y(n3200) );
  AND2X2 U3027 ( .A(\data_in<2> ), .B(n1720), .Y(n3201) );
  INVX1 U3028 ( .A(n3201), .Y(n3202) );
  AND2X2 U3029 ( .A(n5052), .B(n1720), .Y(n3203) );
  INVX1 U3030 ( .A(n3203), .Y(n3204) );
  AND2X2 U3031 ( .A(n5057), .B(n1720), .Y(n3205) );
  INVX1 U3032 ( .A(n3205), .Y(n3206) );
  AND2X2 U3033 ( .A(n5061), .B(n1720), .Y(n3207) );
  INVX1 U3034 ( .A(n3207), .Y(n3208) );
  AND2X2 U3035 ( .A(n5066), .B(n1720), .Y(n3209) );
  INVX1 U3036 ( .A(n3209), .Y(n3210) );
  AND2X2 U3037 ( .A(n5070), .B(n1720), .Y(n3211) );
  INVX1 U3038 ( .A(n3211), .Y(n3212) );
  AND2X2 U3039 ( .A(n5039), .B(n1722), .Y(n3213) );
  INVX1 U3040 ( .A(n3213), .Y(n3214) );
  AND2X2 U3041 ( .A(n5044), .B(n1722), .Y(n3215) );
  INVX1 U3042 ( .A(n3215), .Y(n3216) );
  AND2X2 U3043 ( .A(\data_in<2> ), .B(n1722), .Y(n3217) );
  INVX1 U3044 ( .A(n3217), .Y(n3218) );
  AND2X2 U3045 ( .A(n5052), .B(n1722), .Y(n3219) );
  INVX1 U3046 ( .A(n3219), .Y(n3220) );
  AND2X2 U3047 ( .A(n5057), .B(n1722), .Y(n3221) );
  INVX1 U3048 ( .A(n3221), .Y(n3222) );
  AND2X2 U3049 ( .A(n5061), .B(n1722), .Y(n3223) );
  INVX1 U3050 ( .A(n3223), .Y(n3224) );
  AND2X2 U3051 ( .A(n5066), .B(n1722), .Y(n3225) );
  INVX1 U3052 ( .A(n3225), .Y(n3226) );
  AND2X2 U3053 ( .A(n5070), .B(n1722), .Y(n3227) );
  INVX1 U3054 ( .A(n3227), .Y(n3228) );
  AND2X2 U3055 ( .A(n5039), .B(n1724), .Y(n3229) );
  INVX1 U3056 ( .A(n3229), .Y(n3230) );
  AND2X2 U3057 ( .A(n5044), .B(n1724), .Y(n3231) );
  INVX1 U3058 ( .A(n3231), .Y(n3232) );
  AND2X2 U3059 ( .A(\data_in<2> ), .B(n1724), .Y(n3233) );
  INVX1 U3060 ( .A(n3233), .Y(n3234) );
  AND2X2 U3061 ( .A(n5052), .B(n1724), .Y(n3235) );
  INVX1 U3062 ( .A(n3235), .Y(n3236) );
  AND2X2 U3063 ( .A(n5057), .B(n1724), .Y(n3237) );
  INVX1 U3064 ( .A(n3237), .Y(n3238) );
  AND2X2 U3065 ( .A(n5061), .B(n1724), .Y(n3239) );
  INVX1 U3066 ( .A(n3239), .Y(n3240) );
  AND2X2 U3067 ( .A(n5066), .B(n1724), .Y(n3241) );
  INVX1 U3068 ( .A(n3241), .Y(n3242) );
  AND2X2 U3069 ( .A(n5070), .B(n1724), .Y(n3243) );
  INVX1 U3070 ( .A(n3243), .Y(n3244) );
  AND2X2 U3071 ( .A(n5039), .B(n1726), .Y(n3245) );
  INVX1 U3072 ( .A(n3245), .Y(n3246) );
  AND2X2 U3073 ( .A(n5044), .B(n1726), .Y(n3247) );
  INVX1 U3074 ( .A(n3247), .Y(n3248) );
  AND2X2 U3075 ( .A(\data_in<2> ), .B(n1726), .Y(n3249) );
  INVX1 U3076 ( .A(n3249), .Y(n3250) );
  AND2X2 U3077 ( .A(n5052), .B(n1726), .Y(n3251) );
  INVX1 U3078 ( .A(n3251), .Y(n3252) );
  AND2X2 U3079 ( .A(n5057), .B(n1726), .Y(n3253) );
  INVX1 U3080 ( .A(n3253), .Y(n3254) );
  AND2X2 U3081 ( .A(n5061), .B(n1726), .Y(n3255) );
  INVX1 U3082 ( .A(n3255), .Y(n3256) );
  AND2X2 U3083 ( .A(n5066), .B(n1726), .Y(n3257) );
  INVX1 U3084 ( .A(n3257), .Y(n3258) );
  AND2X2 U3085 ( .A(n5070), .B(n1726), .Y(n3259) );
  INVX1 U3086 ( .A(n3259), .Y(n3260) );
  AND2X2 U3087 ( .A(n5039), .B(n1732), .Y(n3261) );
  INVX1 U3088 ( .A(n3261), .Y(n3262) );
  AND2X2 U3089 ( .A(n5044), .B(n1732), .Y(n3263) );
  INVX1 U3090 ( .A(n3263), .Y(n3264) );
  AND2X2 U3091 ( .A(\data_in<2> ), .B(n1732), .Y(n3265) );
  INVX1 U3092 ( .A(n3265), .Y(n3266) );
  AND2X2 U3093 ( .A(n5052), .B(n1732), .Y(n3267) );
  INVX1 U3094 ( .A(n3267), .Y(n3268) );
  AND2X2 U3095 ( .A(n5057), .B(n1732), .Y(n3269) );
  INVX1 U3096 ( .A(n3269), .Y(n3270) );
  AND2X2 U3097 ( .A(n5061), .B(n1732), .Y(n3271) );
  INVX1 U3098 ( .A(n3271), .Y(n3272) );
  AND2X2 U3099 ( .A(n5066), .B(n1732), .Y(n3273) );
  INVX1 U3100 ( .A(n3273), .Y(n3274) );
  AND2X2 U3101 ( .A(n5070), .B(n1732), .Y(n3275) );
  INVX1 U3102 ( .A(n3275), .Y(n3276) );
  AND2X2 U3103 ( .A(n5039), .B(n1734), .Y(n3277) );
  INVX1 U3104 ( .A(n3277), .Y(n3278) );
  AND2X2 U3105 ( .A(n5044), .B(n1734), .Y(n3279) );
  INVX1 U3106 ( .A(n3279), .Y(n3280) );
  AND2X2 U3107 ( .A(\data_in<2> ), .B(n1734), .Y(n3281) );
  INVX1 U3108 ( .A(n3281), .Y(n3282) );
  AND2X2 U3109 ( .A(n5052), .B(n1734), .Y(n3283) );
  INVX1 U3110 ( .A(n3283), .Y(n3284) );
  AND2X2 U3111 ( .A(n5057), .B(n1734), .Y(n3285) );
  INVX1 U3112 ( .A(n3285), .Y(n3286) );
  AND2X2 U3113 ( .A(n5061), .B(n1734), .Y(n3287) );
  INVX1 U3114 ( .A(n3287), .Y(n3288) );
  AND2X2 U3115 ( .A(n5066), .B(n1734), .Y(n3289) );
  INVX1 U3116 ( .A(n3289), .Y(n3290) );
  AND2X2 U3117 ( .A(n5070), .B(n1734), .Y(n3291) );
  INVX1 U3118 ( .A(n3291), .Y(n3292) );
  AND2X2 U3119 ( .A(n5039), .B(n1736), .Y(n3293) );
  INVX1 U3120 ( .A(n3293), .Y(n3294) );
  AND2X2 U3121 ( .A(n5044), .B(n1736), .Y(n3295) );
  INVX1 U3122 ( .A(n3295), .Y(n3296) );
  AND2X2 U3123 ( .A(\data_in<2> ), .B(n1736), .Y(n3297) );
  INVX1 U3124 ( .A(n3297), .Y(n3298) );
  AND2X2 U3125 ( .A(n5052), .B(n1736), .Y(n3299) );
  INVX1 U3126 ( .A(n3299), .Y(n3300) );
  AND2X2 U3127 ( .A(n5057), .B(n1736), .Y(n3301) );
  INVX1 U3128 ( .A(n3301), .Y(n3302) );
  AND2X2 U3129 ( .A(n5061), .B(n1736), .Y(n3303) );
  INVX1 U3130 ( .A(n3303), .Y(n3304) );
  AND2X2 U3131 ( .A(n5066), .B(n1736), .Y(n3305) );
  INVX1 U3132 ( .A(n3305), .Y(n3306) );
  AND2X2 U3133 ( .A(n5070), .B(n1736), .Y(n3307) );
  INVX1 U3134 ( .A(n3307), .Y(n3308) );
  AND2X2 U3135 ( .A(n5038), .B(n1742), .Y(n3309) );
  INVX1 U3136 ( .A(n3309), .Y(n3310) );
  AND2X2 U3137 ( .A(n5043), .B(n1742), .Y(n3311) );
  INVX1 U3138 ( .A(n3311), .Y(n3312) );
  AND2X2 U3139 ( .A(n5049), .B(n1742), .Y(n3313) );
  INVX1 U3140 ( .A(n3313), .Y(n3314) );
  AND2X2 U3141 ( .A(n5053), .B(n1742), .Y(n3315) );
  INVX1 U3142 ( .A(n3315), .Y(n3316) );
  AND2X2 U3143 ( .A(n5055), .B(n1742), .Y(n3317) );
  INVX1 U3144 ( .A(n3317), .Y(n3318) );
  AND2X2 U3145 ( .A(n5060), .B(n1742), .Y(n3319) );
  INVX1 U3146 ( .A(n3319), .Y(n3320) );
  AND2X2 U3147 ( .A(n5064), .B(n1742), .Y(n3321) );
  INVX1 U3148 ( .A(n3321), .Y(n3322) );
  AND2X2 U3149 ( .A(n5069), .B(n1742), .Y(n3323) );
  INVX1 U3150 ( .A(n3323), .Y(n3324) );
  AND2X2 U3151 ( .A(n5073), .B(n3715), .Y(n3325) );
  INVX1 U3152 ( .A(n3325), .Y(n3326) );
  AND2X2 U3153 ( .A(n5078), .B(n3715), .Y(n3327) );
  INVX1 U3154 ( .A(n3327), .Y(n3328) );
  AND2X2 U3155 ( .A(n5082), .B(n3715), .Y(n3329) );
  INVX1 U3156 ( .A(n3329), .Y(n3330) );
  AND2X2 U3157 ( .A(n5087), .B(n3715), .Y(n3331) );
  INVX1 U3158 ( .A(n3331), .Y(n3332) );
  AND2X2 U3159 ( .A(n5095), .B(n3715), .Y(n3333) );
  INVX1 U3160 ( .A(n3333), .Y(n3334) );
  AND2X2 U3161 ( .A(n5099), .B(n3715), .Y(n3335) );
  INVX1 U3162 ( .A(n3335), .Y(n3336) );
  AND2X2 U3163 ( .A(n5103), .B(n3715), .Y(n3337) );
  INVX1 U3164 ( .A(n3337), .Y(n3338) );
  AND2X2 U3165 ( .A(n5107), .B(n3715), .Y(n3339) );
  INVX1 U3166 ( .A(n3339), .Y(n3340) );
  AND2X2 U3167 ( .A(n5038), .B(n1751), .Y(n3341) );
  INVX1 U3168 ( .A(n3341), .Y(n3342) );
  AND2X2 U3169 ( .A(n5043), .B(n1751), .Y(n3343) );
  INVX1 U3170 ( .A(n3343), .Y(n3344) );
  AND2X2 U3171 ( .A(n5049), .B(n1751), .Y(n3345) );
  INVX1 U3172 ( .A(n3345), .Y(n3346) );
  AND2X2 U3173 ( .A(n5053), .B(n1751), .Y(n3347) );
  INVX1 U3174 ( .A(n3347), .Y(n3348) );
  AND2X2 U3175 ( .A(n5056), .B(n1751), .Y(n3349) );
  INVX1 U3176 ( .A(n3349), .Y(n3350) );
  AND2X2 U3177 ( .A(n5060), .B(n1751), .Y(n3351) );
  INVX1 U3178 ( .A(n3351), .Y(n3352) );
  AND2X2 U3179 ( .A(n5065), .B(n1751), .Y(n3353) );
  INVX1 U3180 ( .A(n3353), .Y(n3354) );
  AND2X2 U3181 ( .A(n5069), .B(n1751), .Y(n3355) );
  INVX1 U3182 ( .A(n3355), .Y(n3356) );
  AND2X2 U3183 ( .A(n5038), .B(n50), .Y(n3357) );
  INVX1 U3184 ( .A(n3357), .Y(n3358) );
  AND2X2 U3185 ( .A(n5043), .B(n50), .Y(n3359) );
  INVX1 U3186 ( .A(n3359), .Y(n3360) );
  AND2X2 U3187 ( .A(n5049), .B(n50), .Y(n3361) );
  INVX1 U3188 ( .A(n3361), .Y(n3362) );
  AND2X2 U3189 ( .A(n5053), .B(n1753), .Y(n3363) );
  INVX1 U3190 ( .A(n3363), .Y(n3364) );
  AND2X2 U3191 ( .A(n5056), .B(n1753), .Y(n3365) );
  INVX1 U3192 ( .A(n3365), .Y(n3366) );
  AND2X2 U3193 ( .A(n5060), .B(n50), .Y(n3367) );
  INVX1 U3194 ( .A(n3367), .Y(n3368) );
  AND2X2 U3195 ( .A(n5064), .B(n1753), .Y(n3369) );
  INVX1 U3196 ( .A(n3369), .Y(n3370) );
  AND2X2 U3197 ( .A(n5069), .B(n50), .Y(n3371) );
  INVX1 U3198 ( .A(n3371), .Y(n3372) );
  AND2X2 U3199 ( .A(n5038), .B(n1762), .Y(n3373) );
  INVX1 U3200 ( .A(n3373), .Y(n3374) );
  AND2X2 U3201 ( .A(n5042), .B(n1762), .Y(n3375) );
  INVX1 U3202 ( .A(n3375), .Y(n3376) );
  AND2X2 U3203 ( .A(n5048), .B(n1762), .Y(n3377) );
  INVX1 U3204 ( .A(n3377), .Y(n3378) );
  AND2X2 U3205 ( .A(n5052), .B(n1762), .Y(n3379) );
  INVX1 U3206 ( .A(n3379), .Y(n3380) );
  AND2X2 U3207 ( .A(n5056), .B(n1762), .Y(n3381) );
  INVX1 U3208 ( .A(n3381), .Y(n3382) );
  AND2X2 U3209 ( .A(n5060), .B(n1762), .Y(n3383) );
  INVX1 U3210 ( .A(n3383), .Y(n3384) );
  AND2X2 U3211 ( .A(n5065), .B(n1762), .Y(n3385) );
  INVX1 U3212 ( .A(n3385), .Y(n3386) );
  AND2X2 U3213 ( .A(n5069), .B(n1762), .Y(n3387) );
  INVX1 U3214 ( .A(n3387), .Y(n3388) );
  AND2X2 U3215 ( .A(n5038), .B(n1764), .Y(n3389) );
  INVX1 U3216 ( .A(n3389), .Y(n3390) );
  AND2X2 U3217 ( .A(n5042), .B(n1764), .Y(n3391) );
  INVX1 U3218 ( .A(n3391), .Y(n3392) );
  AND2X2 U3219 ( .A(n5048), .B(n1764), .Y(n3393) );
  INVX1 U3220 ( .A(n3393), .Y(n3394) );
  AND2X2 U3221 ( .A(n5052), .B(n1764), .Y(n3395) );
  INVX1 U3222 ( .A(n3395), .Y(n3396) );
  AND2X2 U3223 ( .A(n5056), .B(n1764), .Y(n3397) );
  INVX1 U3224 ( .A(n3397), .Y(n3398) );
  AND2X2 U3225 ( .A(n5060), .B(n1764), .Y(n3399) );
  INVX1 U3226 ( .A(n3399), .Y(n3400) );
  AND2X2 U3227 ( .A(n5065), .B(n1764), .Y(n3401) );
  INVX1 U3228 ( .A(n3401), .Y(n3402) );
  AND2X2 U3229 ( .A(n5069), .B(n1764), .Y(n3403) );
  INVX1 U3230 ( .A(n3403), .Y(n3404) );
  AND2X2 U3231 ( .A(n5038), .B(n1770), .Y(n3405) );
  INVX1 U3232 ( .A(n3405), .Y(n3406) );
  AND2X2 U3233 ( .A(n5042), .B(n1770), .Y(n3407) );
  INVX1 U3234 ( .A(n3407), .Y(n3408) );
  AND2X2 U3235 ( .A(n5048), .B(n1770), .Y(n3409) );
  INVX1 U3236 ( .A(n3409), .Y(n3410) );
  AND2X2 U3237 ( .A(n5052), .B(n1770), .Y(n3411) );
  INVX1 U3238 ( .A(n3411), .Y(n3412) );
  AND2X2 U3239 ( .A(n5056), .B(n1770), .Y(n3413) );
  INVX1 U3240 ( .A(n3413), .Y(n3414) );
  AND2X2 U3241 ( .A(n5060), .B(n1770), .Y(n3415) );
  INVX1 U3242 ( .A(n3415), .Y(n3416) );
  AND2X2 U3243 ( .A(n5065), .B(n1770), .Y(n3417) );
  INVX1 U3244 ( .A(n3417), .Y(n3418) );
  AND2X2 U3245 ( .A(n5069), .B(n1770), .Y(n3419) );
  INVX1 U3246 ( .A(n3419), .Y(n3420) );
  AND2X2 U3247 ( .A(n5038), .B(n1774), .Y(n3421) );
  INVX1 U3248 ( .A(n3421), .Y(n3422) );
  AND2X2 U3249 ( .A(n5042), .B(n1774), .Y(n3423) );
  INVX1 U3250 ( .A(n3423), .Y(n3424) );
  AND2X2 U3251 ( .A(n5048), .B(n1774), .Y(n3425) );
  INVX1 U3252 ( .A(n3425), .Y(n3426) );
  AND2X2 U3253 ( .A(n5038), .B(n1777), .Y(n3427) );
  INVX1 U3254 ( .A(n3427), .Y(n3428) );
  AND2X2 U3255 ( .A(n5042), .B(n1777), .Y(n3429) );
  INVX1 U3256 ( .A(n3429), .Y(n3430) );
  AND2X2 U3257 ( .A(n5048), .B(n1777), .Y(n3431) );
  INVX1 U3258 ( .A(n3431), .Y(n3432) );
  AND2X2 U3259 ( .A(n5052), .B(n1777), .Y(n3433) );
  INVX1 U3260 ( .A(n3433), .Y(n3434) );
  AND2X2 U3261 ( .A(n5056), .B(n1777), .Y(n3435) );
  INVX1 U3262 ( .A(n3435), .Y(n3436) );
  AND2X2 U3263 ( .A(n5060), .B(n1777), .Y(n3437) );
  INVX1 U3264 ( .A(n3437), .Y(n3438) );
  AND2X2 U3265 ( .A(n5065), .B(n1777), .Y(n3439) );
  INVX1 U3266 ( .A(n3439), .Y(n3440) );
  AND2X2 U3267 ( .A(n5069), .B(n1777), .Y(n3441) );
  INVX1 U3268 ( .A(n3441), .Y(n3442) );
  AND2X2 U3269 ( .A(n5038), .B(n1779), .Y(n3443) );
  INVX1 U3270 ( .A(n3443), .Y(n3444) );
  AND2X2 U3271 ( .A(n5042), .B(n1779), .Y(n3445) );
  INVX1 U3272 ( .A(n3445), .Y(n3446) );
  AND2X2 U3273 ( .A(n5048), .B(n1779), .Y(n3447) );
  INVX1 U3274 ( .A(n3447), .Y(n3448) );
  AND2X2 U3275 ( .A(n5052), .B(n1779), .Y(n3449) );
  INVX1 U3276 ( .A(n3449), .Y(n3450) );
  AND2X2 U3277 ( .A(n5056), .B(n1779), .Y(n3451) );
  INVX1 U3278 ( .A(n3451), .Y(n3452) );
  AND2X2 U3279 ( .A(n5060), .B(n1779), .Y(n3453) );
  INVX1 U3280 ( .A(n3453), .Y(n3454) );
  AND2X2 U3281 ( .A(n5065), .B(n1779), .Y(n3455) );
  INVX1 U3282 ( .A(n3455), .Y(n3456) );
  AND2X2 U3283 ( .A(n5069), .B(n1779), .Y(n3457) );
  INVX1 U3284 ( .A(n3457), .Y(n3458) );
  AND2X2 U3285 ( .A(n5038), .B(n1785), .Y(n3459) );
  INVX1 U3286 ( .A(n3459), .Y(n3460) );
  AND2X2 U3287 ( .A(n5041), .B(n1785), .Y(n3461) );
  INVX1 U3288 ( .A(n3461), .Y(n3462) );
  AND2X2 U3289 ( .A(n5047), .B(n1785), .Y(n3463) );
  INVX1 U3290 ( .A(n3463), .Y(n3464) );
  AND2X2 U3291 ( .A(n5051), .B(n1785), .Y(n3465) );
  INVX1 U3292 ( .A(n3465), .Y(n3466) );
  AND2X2 U3293 ( .A(n5055), .B(n1785), .Y(n3467) );
  INVX1 U3294 ( .A(n3467), .Y(n3468) );
  AND2X2 U3295 ( .A(n5060), .B(n1785), .Y(n3469) );
  INVX1 U3296 ( .A(n3469), .Y(n3470) );
  AND2X2 U3297 ( .A(n5064), .B(n1785), .Y(n3471) );
  INVX1 U3298 ( .A(n3471), .Y(n3472) );
  AND2X2 U3299 ( .A(n5069), .B(n1785), .Y(n3473) );
  INVX1 U3300 ( .A(n3473), .Y(n3474) );
  AND2X2 U3301 ( .A(n5038), .B(n1787), .Y(n3475) );
  INVX1 U3302 ( .A(n3475), .Y(n3476) );
  AND2X2 U3303 ( .A(n5041), .B(n1787), .Y(n3477) );
  INVX1 U3304 ( .A(n3477), .Y(n3478) );
  AND2X2 U3305 ( .A(n5047), .B(n1787), .Y(n3479) );
  INVX1 U3306 ( .A(n3479), .Y(n3480) );
  AND2X2 U3307 ( .A(n5051), .B(n1787), .Y(n3481) );
  INVX1 U3308 ( .A(n3481), .Y(n3482) );
  AND2X2 U3309 ( .A(n5055), .B(n1787), .Y(n3483) );
  INVX1 U3310 ( .A(n3483), .Y(n3484) );
  AND2X2 U3311 ( .A(n5060), .B(n1787), .Y(n3485) );
  INVX1 U3312 ( .A(n3485), .Y(n3486) );
  AND2X2 U3313 ( .A(n5064), .B(n1787), .Y(n3487) );
  INVX1 U3314 ( .A(n3487), .Y(n3488) );
  AND2X2 U3315 ( .A(n5069), .B(n1787), .Y(n3489) );
  INVX1 U3316 ( .A(n3489), .Y(n3490) );
  AND2X2 U3317 ( .A(n5069), .B(n1789), .Y(n3491) );
  INVX1 U3318 ( .A(n3491), .Y(n3492) );
  AND2X2 U3319 ( .A(n5038), .B(n1791), .Y(n3493) );
  INVX1 U3320 ( .A(n3493), .Y(n3494) );
  AND2X2 U3321 ( .A(n5041), .B(n1791), .Y(n3495) );
  INVX1 U3322 ( .A(n3495), .Y(n3496) );
  AND2X2 U3323 ( .A(n5047), .B(n1791), .Y(n3497) );
  INVX1 U3324 ( .A(n3497), .Y(n3498) );
  AND2X2 U3325 ( .A(n5051), .B(n1791), .Y(n3499) );
  INVX1 U3326 ( .A(n3499), .Y(n3500) );
  AND2X2 U3327 ( .A(n5055), .B(n1791), .Y(n3501) );
  INVX1 U3328 ( .A(n3501), .Y(n3502) );
  AND2X2 U3329 ( .A(n5060), .B(n1791), .Y(n3503) );
  INVX1 U3330 ( .A(n3503), .Y(n3504) );
  AND2X2 U3331 ( .A(n5064), .B(n1791), .Y(n3505) );
  INVX1 U3332 ( .A(n3505), .Y(n3506) );
  AND2X2 U3333 ( .A(n5069), .B(n1791), .Y(n3507) );
  INVX1 U3334 ( .A(n3507), .Y(n3508) );
  AND2X2 U3335 ( .A(n5038), .B(n1793), .Y(n3509) );
  INVX1 U3336 ( .A(n3509), .Y(n3510) );
  AND2X2 U3337 ( .A(n5041), .B(n1793), .Y(n3511) );
  INVX1 U3338 ( .A(n3511), .Y(n3512) );
  AND2X2 U3339 ( .A(n5047), .B(n1793), .Y(n3513) );
  INVX1 U3340 ( .A(n3513), .Y(n3514) );
  AND2X2 U3341 ( .A(n5051), .B(n1793), .Y(n3515) );
  INVX1 U3342 ( .A(n3515), .Y(n3516) );
  AND2X2 U3343 ( .A(n5055), .B(n1793), .Y(n3517) );
  INVX1 U3344 ( .A(n3517), .Y(n3518) );
  AND2X2 U3345 ( .A(n5060), .B(n1793), .Y(n3519) );
  INVX1 U3346 ( .A(n3519), .Y(n3520) );
  AND2X2 U3347 ( .A(n5064), .B(n1793), .Y(n3521) );
  INVX1 U3348 ( .A(n3521), .Y(n3522) );
  AND2X2 U3349 ( .A(n5069), .B(n1793), .Y(n3523) );
  INVX1 U3350 ( .A(n3523), .Y(n3524) );
  AND2X2 U3351 ( .A(n5038), .B(n1795), .Y(n3525) );
  INVX1 U3352 ( .A(n3525), .Y(n3526) );
  AND2X2 U3353 ( .A(n5041), .B(n1795), .Y(n3527) );
  INVX1 U3354 ( .A(n3527), .Y(n3528) );
  AND2X2 U3355 ( .A(n5047), .B(n1795), .Y(n3529) );
  INVX1 U3356 ( .A(n3529), .Y(n3530) );
  AND2X2 U3357 ( .A(n5051), .B(n1795), .Y(n3531) );
  INVX1 U3358 ( .A(n3531), .Y(n3532) );
  AND2X2 U3359 ( .A(n5055), .B(n1795), .Y(n3533) );
  INVX1 U3360 ( .A(n3533), .Y(n3534) );
  AND2X2 U3361 ( .A(n5060), .B(n1795), .Y(n3535) );
  INVX1 U3362 ( .A(n3535), .Y(n3536) );
  AND2X2 U3363 ( .A(n5064), .B(n1795), .Y(n3537) );
  INVX1 U3364 ( .A(n3537), .Y(n3538) );
  AND2X2 U3365 ( .A(n5069), .B(n1795), .Y(n3539) );
  INVX1 U3366 ( .A(n3539), .Y(n3540) );
  AND2X2 U3367 ( .A(n5038), .B(n1801), .Y(n3541) );
  INVX1 U3368 ( .A(n3541), .Y(n3542) );
  AND2X2 U3369 ( .A(n5041), .B(n1801), .Y(n3543) );
  INVX1 U3370 ( .A(n3543), .Y(n3544) );
  AND2X2 U3371 ( .A(n5047), .B(n1801), .Y(n3545) );
  INVX1 U3372 ( .A(n3545), .Y(n3546) );
  AND2X2 U3373 ( .A(n5051), .B(n1801), .Y(n3547) );
  INVX1 U3374 ( .A(n3547), .Y(n3548) );
  AND2X2 U3375 ( .A(n5055), .B(n1801), .Y(n3549) );
  INVX1 U3376 ( .A(n3549), .Y(n3550) );
  AND2X2 U3377 ( .A(n5060), .B(n1801), .Y(n3551) );
  INVX1 U3378 ( .A(n3551), .Y(n3552) );
  AND2X2 U3379 ( .A(n5064), .B(n1801), .Y(n3553) );
  INVX1 U3380 ( .A(n3553), .Y(n3554) );
  AND2X2 U3381 ( .A(n5069), .B(n1801), .Y(n3555) );
  INVX1 U3382 ( .A(n3555), .Y(n3556) );
  INVX1 U3383 ( .A(n5724), .Y(n3557) );
  INVX1 U3384 ( .A(n5725), .Y(n3558) );
  AND2X2 U3385 ( .A(n4957), .B(n3661), .Y(n3559) );
  INVX1 U3386 ( .A(n3559), .Y(n3560) );
  AND2X2 U3387 ( .A(n4969), .B(n3661), .Y(n3561) );
  INVX1 U3388 ( .A(n3561), .Y(n3562) );
  OR2X2 U3389 ( .A(n103), .B(n6352), .Y(n3563) );
  INVX1 U3390 ( .A(n3563), .Y(n3564) );
  AND2X2 U3391 ( .A(n4884), .B(n4767), .Y(n3565) );
  INVX1 U3392 ( .A(n3565), .Y(n3566) );
  OR2X2 U3393 ( .A(n4754), .B(n133), .Y(n3567) );
  INVX1 U3394 ( .A(n3567), .Y(n3568) );
  BUFX2 U3395 ( .A(n5180), .Y(n3569) );
  BUFX2 U3396 ( .A(n5284), .Y(n3570) );
  BUFX2 U3397 ( .A(n5347), .Y(n3571) );
  OR2X2 U3398 ( .A(n81), .B(n103), .Y(n3572) );
  AND2X2 U3399 ( .A(n4949), .B(n4967), .Y(n3573) );
  INVX1 U3400 ( .A(n3573), .Y(n3574) );
  OR2X2 U3401 ( .A(n6352), .B(n103), .Y(n3575) );
  INVX1 U3402 ( .A(n3575), .Y(n3576) );
  AND2X2 U3403 ( .A(n562), .B(n80), .Y(n3577) );
  AND2X2 U3404 ( .A(n1064), .B(n4973), .Y(n3579) );
  AND2X2 U3405 ( .A(n1066), .B(n4973), .Y(n3581) );
  INVX1 U3406 ( .A(n3581), .Y(n3582) );
  AND2X2 U3407 ( .A(n1068), .B(n4973), .Y(n3583) );
  AND2X2 U3408 ( .A(n6311), .B(n4973), .Y(n3585) );
  AND2X2 U3409 ( .A(n1070), .B(n4973), .Y(n3587) );
  INVX1 U3410 ( .A(n3587), .Y(n3588) );
  AND2X2 U3411 ( .A(n1072), .B(n4973), .Y(n3589) );
  INVX1 U3412 ( .A(n3589), .Y(n3590) );
  AND2X2 U3413 ( .A(n1074), .B(n4973), .Y(n3591) );
  AND2X2 U3414 ( .A(n1076), .B(n4973), .Y(n3593) );
  AND2X2 U3415 ( .A(n1078), .B(n4973), .Y(n3595) );
  AND2X2 U3416 ( .A(n1080), .B(n4973), .Y(n3597) );
  AND2X2 U3417 ( .A(n1082), .B(n4973), .Y(n3599) );
  INVX1 U3418 ( .A(n3599), .Y(n3600) );
  AND2X2 U3419 ( .A(n1084), .B(n4973), .Y(n3601) );
  INVX1 U3420 ( .A(n3601), .Y(n3602) );
  AND2X2 U3421 ( .A(n1086), .B(n4974), .Y(n3603) );
  INVX1 U3422 ( .A(n3603), .Y(n3604) );
  AND2X2 U3423 ( .A(n1088), .B(n4974), .Y(n3605) );
  INVX1 U3424 ( .A(n3605), .Y(n3606) );
  AND2X2 U3425 ( .A(n1090), .B(n4974), .Y(n3607) );
  INVX1 U3426 ( .A(n3607), .Y(n3608) );
  AND2X2 U3427 ( .A(n1092), .B(n4974), .Y(n3609) );
  AND2X2 U3428 ( .A(n1094), .B(n4974), .Y(n3611) );
  INVX1 U3429 ( .A(n3611), .Y(n3612) );
  AND2X2 U3430 ( .A(n1096), .B(n4974), .Y(n3613) );
  AND2X2 U3431 ( .A(n4974), .B(n1098), .Y(n3615) );
  AND2X2 U3432 ( .A(n1100), .B(n4974), .Y(n3617) );
  AND2X2 U3433 ( .A(n4974), .B(n1102), .Y(n3619) );
  AND2X2 U3434 ( .A(n1104), .B(n4974), .Y(n3621) );
  AND2X2 U3435 ( .A(n4974), .B(n1106), .Y(n3623) );
  AND2X2 U3436 ( .A(n1108), .B(n4975), .Y(n3625) );
  AND2X2 U3437 ( .A(n1110), .B(n4975), .Y(n3627) );
  AND2X2 U3438 ( .A(n1112), .B(n4975), .Y(n3629) );
  INVX1 U3439 ( .A(n3629), .Y(n3630) );
  AND2X2 U3440 ( .A(n1114), .B(n4975), .Y(n3631) );
  AND2X2 U3441 ( .A(n4975), .B(n1116), .Y(n3633) );
  INVX1 U3442 ( .A(n3633), .Y(n3634) );
  AND2X2 U3443 ( .A(n4975), .B(n1118), .Y(n3635) );
  INVX1 U3444 ( .A(n3635), .Y(n3636) );
  AND2X2 U3445 ( .A(n1120), .B(n4975), .Y(n3637) );
  AND2X2 U3446 ( .A(n1122), .B(n4976), .Y(n3639) );
  INVX1 U3447 ( .A(n3639), .Y(n3640) );
  AND2X2 U3448 ( .A(n1124), .B(n4976), .Y(n3641) );
  INVX1 U3449 ( .A(n3641), .Y(n3642) );
  AND2X2 U3450 ( .A(n1126), .B(n4975), .Y(n3643) );
  INVX1 U3451 ( .A(n3643), .Y(n3644) );
  AND2X2 U3452 ( .A(n1128), .B(n4976), .Y(n3645) );
  INVX1 U3453 ( .A(n3645), .Y(n3646) );
  AND2X2 U3454 ( .A(n1130), .B(n4975), .Y(n3647) );
  INVX1 U3455 ( .A(n3647), .Y(n3648) );
  OR2X2 U3456 ( .A(n4764), .B(n3870), .Y(n3649) );
  INVX1 U3457 ( .A(n3649), .Y(n3650) );
  INVX1 U3458 ( .A(n3649), .Y(n3651) );
  OR2X2 U3459 ( .A(n560), .B(n4735), .Y(n3652) );
  OR2X2 U3460 ( .A(n4673), .B(n750), .Y(n3653) );
  OR2X2 U3461 ( .A(n4724), .B(n4725), .Y(n3655) );
  INVX1 U3462 ( .A(n3655), .Y(n3656) );
  INVX1 U3463 ( .A(n3655), .Y(n3657) );
  OR2X2 U3464 ( .A(n4815), .B(n3874), .Y(n3658) );
  INVX1 U3465 ( .A(n3658), .Y(n3659) );
  OR2X2 U3466 ( .A(n4980), .B(n4628), .Y(n3660) );
  OR2X2 U3467 ( .A(n115), .B(n748), .Y(n3662) );
  OR2X2 U3468 ( .A(n6288), .B(n750), .Y(n3664) );
  AND2X2 U3469 ( .A(n1055), .B(n4975), .Y(n3666) );
  INVX1 U3470 ( .A(n3666), .Y(n3667) );
  AND2X2 U3471 ( .A(n122), .B(n4873), .Y(n3668) );
  OR2X2 U3472 ( .A(n4623), .B(n4955), .Y(n3670) );
  INVX1 U3473 ( .A(n3670), .Y(n3671) );
  INVX1 U3474 ( .A(n3670), .Y(n3672) );
  OR2X2 U3475 ( .A(n4867), .B(n749), .Y(n3673) );
  AND2X2 U3476 ( .A(n45), .B(n5167), .Y(n3674) );
  INVX1 U3477 ( .A(n3674), .Y(n3675) );
  INVX1 U3478 ( .A(n3674), .Y(n3676) );
  INVX1 U3479 ( .A(n6333), .Y(n3677) );
  BUFX2 U3480 ( .A(n3567), .Y(n4917) );
  AND2X2 U3481 ( .A(n54), .B(n5726), .Y(n3678) );
  INVX1 U3482 ( .A(n3678), .Y(n3679) );
  AND2X2 U3483 ( .A(\mem<16><0> ), .B(n4816), .Y(n3680) );
  INVX1 U3484 ( .A(n3680), .Y(n3681) );
  AND2X2 U3485 ( .A(\mem<16><1> ), .B(n4816), .Y(n3682) );
  INVX1 U3486 ( .A(n3682), .Y(n3683) );
  AND2X2 U3487 ( .A(\mem<43><7> ), .B(n151), .Y(n3684) );
  INVX1 U3488 ( .A(n3684), .Y(n3685) );
  INVX1 U3489 ( .A(n5437), .Y(n3686) );
  INVX1 U3490 ( .A(n3686), .Y(n3687) );
  AND2X2 U3491 ( .A(n5038), .B(n1746), .Y(n3688) );
  INVX1 U3492 ( .A(n3688), .Y(n3689) );
  AND2X2 U3493 ( .A(n5043), .B(n1746), .Y(n3690) );
  INVX1 U3494 ( .A(n3690), .Y(n3691) );
  AND2X2 U3495 ( .A(n5053), .B(n1746), .Y(n3692) );
  INVX1 U3496 ( .A(n3692), .Y(n3693) );
  AND2X2 U3497 ( .A(n5069), .B(n1746), .Y(n3694) );
  INVX1 U3498 ( .A(n3694), .Y(n3695) );
  AND2X2 U3499 ( .A(n5075), .B(n3719), .Y(n3696) );
  INVX1 U3500 ( .A(n3696), .Y(n3697) );
  AND2X2 U3501 ( .A(n5079), .B(n3719), .Y(n3698) );
  INVX1 U3502 ( .A(n3698), .Y(n3699) );
  AND2X2 U3503 ( .A(n5085), .B(n3719), .Y(n3700) );
  INVX1 U3504 ( .A(n3700), .Y(n3701) );
  AND2X2 U3505 ( .A(n5090), .B(n3719), .Y(n3702) );
  INVX1 U3506 ( .A(n3702), .Y(n3703) );
  AND2X2 U3507 ( .A(n5096), .B(n3719), .Y(n3704) );
  INVX1 U3508 ( .A(n3704), .Y(n3705) );
  AND2X2 U3509 ( .A(n5100), .B(n3719), .Y(n3706) );
  INVX1 U3510 ( .A(n3706), .Y(n3707) );
  AND2X2 U3511 ( .A(n5104), .B(n3719), .Y(n3708) );
  INVX1 U3512 ( .A(n3708), .Y(n3709) );
  AND2X2 U3513 ( .A(n5109), .B(n3719), .Y(n3710) );
  INVX1 U3514 ( .A(n3710), .Y(n3711) );
  AND2X2 U3515 ( .A(n3861), .B(n5033), .Y(n3712) );
  AND2X2 U3516 ( .A(n4949), .B(n3), .Y(n3713) );
  AND2X2 U3517 ( .A(n4850), .B(n3591), .Y(n3714) );
  AND2X2 U3518 ( .A(n6347), .B(n6346), .Y(n3715) );
  AND2X2 U3519 ( .A(n4751), .B(n3621), .Y(n3716) );
  AND2X2 U3520 ( .A(n4957), .B(n4967), .Y(n3717) );
  AND2X2 U3521 ( .A(n4961), .B(n4967), .Y(n3718) );
  AND2X2 U3522 ( .A(n3572), .B(n6418), .Y(n3719) );
  AND2X2 U3523 ( .A(\mem<22><3> ), .B(n4957), .Y(n3720) );
  INVX1 U3524 ( .A(n3720), .Y(n3721) );
  AND2X2 U3525 ( .A(\mem<22><4> ), .B(n4957), .Y(n3722) );
  INVX1 U3526 ( .A(n3722), .Y(n3723) );
  AND2X2 U3527 ( .A(\mem<22><5> ), .B(n4959), .Y(n3724) );
  INVX1 U3528 ( .A(n3724), .Y(n3725) );
  AND2X2 U3529 ( .A(\mem<22><6> ), .B(n4957), .Y(n3726) );
  INVX1 U3530 ( .A(n3726), .Y(n3727) );
  AND2X2 U3531 ( .A(n5107), .B(n1699), .Y(n3728) );
  INVX1 U3532 ( .A(n3728), .Y(n3729) );
  AND2X2 U3533 ( .A(n5072), .B(n3855), .Y(n3730) );
  INVX1 U3534 ( .A(n3730), .Y(n3731) );
  AND2X2 U3535 ( .A(n5078), .B(n3855), .Y(n3732) );
  INVX1 U3536 ( .A(n3732), .Y(n3733) );
  AND2X2 U3537 ( .A(n5084), .B(n3855), .Y(n3734) );
  INVX1 U3538 ( .A(n3734), .Y(n3735) );
  AND2X2 U3539 ( .A(n5089), .B(n3855), .Y(n3736) );
  INVX1 U3540 ( .A(n3736), .Y(n3737) );
  AND2X2 U3541 ( .A(n5095), .B(n3855), .Y(n3738) );
  INVX1 U3542 ( .A(n3738), .Y(n3739) );
  AND2X2 U3543 ( .A(n5099), .B(n3855), .Y(n3740) );
  INVX1 U3544 ( .A(n3740), .Y(n3741) );
  AND2X2 U3545 ( .A(n5103), .B(n3855), .Y(n3742) );
  INVX1 U3546 ( .A(n3742), .Y(n3743) );
  AND2X2 U3547 ( .A(n5108), .B(n3855), .Y(n3744) );
  INVX1 U3548 ( .A(n3744), .Y(n3745) );
  AND2X2 U3549 ( .A(n5073), .B(n1748), .Y(n3746) );
  INVX1 U3550 ( .A(n3746), .Y(n3747) );
  AND2X2 U3551 ( .A(n5078), .B(n1748), .Y(n3748) );
  INVX1 U3552 ( .A(n3748), .Y(n3749) );
  AND2X2 U3553 ( .A(n5082), .B(n1748), .Y(n3750) );
  INVX1 U3554 ( .A(n3750), .Y(n3751) );
  AND2X2 U3555 ( .A(n5087), .B(n1748), .Y(n3752) );
  INVX1 U3556 ( .A(n3752), .Y(n3753) );
  AND2X2 U3557 ( .A(n5095), .B(n1748), .Y(n3754) );
  INVX1 U3558 ( .A(n3754), .Y(n3755) );
  AND2X2 U3559 ( .A(n5099), .B(n1748), .Y(n3756) );
  INVX1 U3560 ( .A(n3756), .Y(n3757) );
  AND2X2 U3561 ( .A(n5103), .B(n1748), .Y(n3758) );
  INVX1 U3562 ( .A(n3758), .Y(n3759) );
  AND2X2 U3563 ( .A(n5107), .B(n1748), .Y(n3760) );
  INVX1 U3564 ( .A(n3760), .Y(n3761) );
  AND2X2 U3565 ( .A(n5073), .B(n1750), .Y(n3762) );
  INVX1 U3566 ( .A(n3762), .Y(n3763) );
  AND2X2 U3567 ( .A(n5078), .B(n1750), .Y(n3764) );
  INVX1 U3568 ( .A(n3764), .Y(n3765) );
  AND2X2 U3569 ( .A(n5082), .B(n1750), .Y(n3766) );
  INVX1 U3570 ( .A(n3766), .Y(n3767) );
  AND2X2 U3571 ( .A(n5087), .B(n1750), .Y(n3768) );
  INVX1 U3572 ( .A(n3768), .Y(n3769) );
  AND2X2 U3573 ( .A(n5095), .B(n1750), .Y(n3770) );
  INVX1 U3574 ( .A(n3770), .Y(n3771) );
  AND2X2 U3575 ( .A(n5099), .B(n1750), .Y(n3772) );
  INVX1 U3576 ( .A(n3772), .Y(n3773) );
  AND2X2 U3577 ( .A(n5103), .B(n1750), .Y(n3774) );
  INVX1 U3578 ( .A(n3774), .Y(n3775) );
  AND2X2 U3579 ( .A(n5107), .B(n1750), .Y(n3776) );
  INVX1 U3580 ( .A(n3776), .Y(n3777) );
  INVX1 U3581 ( .A(n1017), .Y(n3778) );
  INVX1 U3582 ( .A(n1018), .Y(n3779) );
  OR2X2 U3583 ( .A(n5458), .B(n5457), .Y(n3780) );
  AND2X2 U3584 ( .A(n5039), .B(n1689), .Y(n3781) );
  INVX1 U3585 ( .A(n3781), .Y(n3782) );
  AND2X2 U3586 ( .A(n5044), .B(n1689), .Y(n3783) );
  INVX1 U3587 ( .A(n3783), .Y(n3784) );
  AND2X2 U3588 ( .A(\data_in<2> ), .B(n1689), .Y(n3785) );
  INVX1 U3589 ( .A(n3785), .Y(n3786) );
  AND2X2 U3590 ( .A(n5052), .B(n1689), .Y(n3787) );
  INVX1 U3591 ( .A(n3787), .Y(n3788) );
  AND2X2 U3592 ( .A(n5057), .B(n1689), .Y(n3789) );
  INVX1 U3593 ( .A(n3789), .Y(n3790) );
  AND2X2 U3594 ( .A(n5061), .B(n1689), .Y(n3791) );
  INVX1 U3595 ( .A(n3791), .Y(n3792) );
  AND2X2 U3596 ( .A(n5066), .B(n1689), .Y(n3793) );
  INVX1 U3597 ( .A(n3793), .Y(n3794) );
  AND2X2 U3598 ( .A(n5070), .B(n1689), .Y(n3795) );
  INVX1 U3599 ( .A(n3795), .Y(n3796) );
  AND2X2 U3600 ( .A(n5039), .B(n1706), .Y(n3797) );
  INVX1 U3601 ( .A(n3797), .Y(n3798) );
  AND2X2 U3602 ( .A(n5045), .B(n1706), .Y(n3799) );
  INVX1 U3603 ( .A(n3799), .Y(n3800) );
  AND2X2 U3604 ( .A(n5053), .B(n1706), .Y(n3801) );
  INVX1 U3605 ( .A(n3801), .Y(n3802) );
  AND2X2 U3606 ( .A(n5070), .B(n1706), .Y(n3803) );
  INVX1 U3607 ( .A(n3803), .Y(n3804) );
  AND2X2 U3608 ( .A(\mem<25><0> ), .B(n3620), .Y(n3805) );
  INVX1 U3609 ( .A(n3805), .Y(n3806) );
  AND2X2 U3610 ( .A(\mem<25><1> ), .B(n3620), .Y(n3807) );
  INVX1 U3611 ( .A(n3807), .Y(n3808) );
  AND2X2 U3612 ( .A(\mem<25><2> ), .B(n3620), .Y(n3809) );
  INVX1 U3613 ( .A(n3809), .Y(n3810) );
  AND2X2 U3614 ( .A(\mem<25><3> ), .B(n3620), .Y(n3811) );
  INVX1 U3615 ( .A(n3811), .Y(n3812) );
  AND2X2 U3616 ( .A(\mem<25><5> ), .B(n3620), .Y(n3813) );
  INVX1 U3617 ( .A(n3813), .Y(n3814) );
  AND2X2 U3618 ( .A(\mem<25><6> ), .B(n3620), .Y(n3815) );
  INVX1 U3619 ( .A(n3815), .Y(n3816) );
  AND2X2 U3620 ( .A(\mem<25><7> ), .B(n3620), .Y(n3817) );
  INVX1 U3621 ( .A(n3817), .Y(n3818) );
  AND2X2 U3622 ( .A(\mem<24><0> ), .B(n3622), .Y(n3819) );
  INVX1 U3623 ( .A(n3819), .Y(n3820) );
  AND2X2 U3624 ( .A(\mem<24><1> ), .B(n3622), .Y(n3821) );
  INVX1 U3625 ( .A(n3821), .Y(n3822) );
  AND2X2 U3626 ( .A(\mem<24><2> ), .B(n3622), .Y(n3823) );
  INVX1 U3627 ( .A(n3823), .Y(n3824) );
  AND2X2 U3628 ( .A(\mem<24><3> ), .B(n3622), .Y(n3825) );
  INVX1 U3629 ( .A(n3825), .Y(n3826) );
  AND2X2 U3630 ( .A(\mem<24><5> ), .B(n3622), .Y(n3827) );
  INVX1 U3631 ( .A(n3827), .Y(n3828) );
  AND2X2 U3632 ( .A(\mem<24><6> ), .B(n3622), .Y(n3829) );
  INVX1 U3633 ( .A(n3829), .Y(n3830) );
  AND2X2 U3634 ( .A(\mem<24><7> ), .B(n3622), .Y(n3831) );
  INVX1 U3635 ( .A(n3831), .Y(n3832) );
  AND2X2 U3636 ( .A(n5038), .B(n1772), .Y(n3833) );
  INVX1 U3637 ( .A(n3833), .Y(n3834) );
  AND2X2 U3638 ( .A(n5042), .B(n1772), .Y(n3835) );
  INVX1 U3639 ( .A(n3835), .Y(n3836) );
  AND2X2 U3640 ( .A(n5048), .B(n1772), .Y(n3837) );
  INVX1 U3641 ( .A(n3837), .Y(n3838) );
  AND2X2 U3642 ( .A(n5052), .B(n1772), .Y(n3839) );
  INVX1 U3643 ( .A(n3839), .Y(n3840) );
  INVX1 U3644 ( .A(n1008), .Y(n3841) );
  AND2X2 U3645 ( .A(n5069), .B(n1772), .Y(n3842) );
  INVX1 U3646 ( .A(n3842), .Y(n3843) );
  INVX1 U3647 ( .A(n4858), .Y(n6352) );
  INVX2 U3648 ( .A(n4968), .Y(n4967) );
  INVX1 U3649 ( .A(n119), .Y(n6332) );
  INVX1 U3650 ( .A(n5203), .Y(n3844) );
  INVX1 U3651 ( .A(n4952), .Y(n3845) );
  INVX1 U3652 ( .A(n953), .Y(n3860) );
  INVX1 U3653 ( .A(n3717), .Y(n3846) );
  INVX2 U3654 ( .A(n1687), .Y(n3847) );
  INVX1 U3655 ( .A(n3651), .Y(n3848) );
  INVX1 U3656 ( .A(n3656), .Y(n3850) );
  INVX1 U3657 ( .A(n3657), .Y(n6367) );
  INVX1 U3658 ( .A(n3659), .Y(n5649) );
  AND2X2 U3659 ( .A(n65), .B(n747), .Y(n4868) );
  INVX1 U3660 ( .A(n6404), .Y(n6405) );
  INVX2 U3661 ( .A(n1684), .Y(n6331) );
  BUFX2 U3662 ( .A(n3850), .Y(n4918) );
  INVX1 U3663 ( .A(n3655), .Y(n6366) );
  NAND3X1 U3664 ( .A(n148), .B(n5203), .C(n4881), .Y(n3852) );
  INVX1 U3665 ( .A(n5013), .Y(n5012) );
  INVX1 U3666 ( .A(\addr<15> ), .Y(n3853) );
  INVX1 U3667 ( .A(n3853), .Y(n3854) );
  BUFX2 U3668 ( .A(n6310), .Y(n4925) );
  AND2X2 U3669 ( .A(n6309), .B(n4652), .Y(n3855) );
  INVX1 U3670 ( .A(n6369), .Y(n3856) );
  INVX1 U3671 ( .A(n6369), .Y(n6368) );
  NAND2X1 U3672 ( .A(\mem<49><2> ), .B(n4835), .Y(n3857) );
  NAND2X1 U3673 ( .A(\mem<9><2> ), .B(n97), .Y(n3858) );
  AND2X2 U3674 ( .A(n3857), .B(n3858), .Y(n5361) );
  AOI21X1 U3675 ( .A(n4655), .B(n6326), .C(n4978), .Y(n3859) );
  INVX1 U3676 ( .A(n6326), .Y(n6328) );
  INVX1 U3677 ( .A(n6401), .Y(n3862) );
  INVX1 U3678 ( .A(n4821), .Y(n3863) );
  INVX1 U3679 ( .A(n797), .Y(n6401) );
  INVX1 U3680 ( .A(n6302), .Y(n3864) );
  INVX1 U3681 ( .A(n4912), .Y(n3865) );
  INVX1 U3682 ( .A(n3865), .Y(n3866) );
  INVX1 U3683 ( .A(n3865), .Y(n3867) );
  INVX1 U3684 ( .A(n3865), .Y(n3868) );
  AND2X2 U3685 ( .A(n1053), .B(n4975), .Y(n3869) );
  INVX4 U3686 ( .A(n3882), .Y(n4966) );
  INVX1 U3687 ( .A(n4813), .Y(n3871) );
  INVX1 U3688 ( .A(n4910), .Y(n6314) );
  NAND2X1 U3689 ( .A(\mem<1><7> ), .B(n4810), .Y(n3872) );
  AND2X2 U3690 ( .A(n3872), .B(n3679), .Y(n5727) );
  INVX1 U3691 ( .A(n4867), .Y(n3874) );
  INVX1 U3692 ( .A(n43), .Y(n3875) );
  INVX1 U3693 ( .A(n3661), .Y(n3876) );
  INVX1 U3694 ( .A(n5192), .Y(n4915) );
  INVX2 U3695 ( .A(n4963), .Y(n4962) );
  AND2X2 U3696 ( .A(n3673), .B(n3650), .Y(n3877) );
  AND2X2 U3697 ( .A(n3673), .B(n3650), .Y(n3878) );
  INVX1 U3698 ( .A(n4855), .Y(n3879) );
  INVX1 U3699 ( .A(n4843), .Y(n3880) );
  INVX1 U3700 ( .A(n6333), .Y(n3881) );
  INVX1 U3701 ( .A(n6410), .Y(n3882) );
  INVX1 U3702 ( .A(n4877), .Y(n6313) );
  AND2X2 U3703 ( .A(n5039), .B(n1713), .Y(n3883) );
  INVX1 U3704 ( .A(n3883), .Y(n3884) );
  AND2X2 U3705 ( .A(n5072), .B(n3714), .Y(n3885) );
  INVX1 U3706 ( .A(n3885), .Y(n3886) );
  OR2X2 U3707 ( .A(n5123), .B(n5122), .Y(n3887) );
  OR2X2 U3708 ( .A(n5238), .B(n5237), .Y(n3888) );
  OR2X2 U3709 ( .A(n5296), .B(n5297), .Y(n3889) );
  INVX1 U3710 ( .A(n3563), .Y(n4916) );
  INVX1 U3711 ( .A(n782), .Y(n6353) );
  NAND2X1 U3712 ( .A(n1216), .B(n751), .Y(n6827) );
  NAND2X1 U3713 ( .A(n1220), .B(n752), .Y(n6826) );
  NAND2X1 U3714 ( .A(n1224), .B(n753), .Y(n6825) );
  NAND2X1 U3715 ( .A(n1228), .B(n754), .Y(n6824) );
  NAND2X1 U3716 ( .A(n1232), .B(n755), .Y(n6823) );
  NAND2X1 U3717 ( .A(n1236), .B(n756), .Y(n6822) );
  NAND2X1 U3718 ( .A(n1240), .B(n757), .Y(n6821) );
  AND2X2 U3719 ( .A(n4904), .B(n5131), .Y(n3890) );
  INVX1 U3720 ( .A(n3890), .Y(n3891) );
  AND2X2 U3721 ( .A(\mem<51><0> ), .B(n4873), .Y(n3892) );
  INVX1 U3722 ( .A(n3892), .Y(n3893) );
  AND2X2 U3723 ( .A(n3851), .B(n5144), .Y(n3894) );
  INVX1 U3724 ( .A(n3894), .Y(n3895) );
  INVX1 U3725 ( .A(n3896), .Y(n3897) );
  AND2X2 U3726 ( .A(\mem<55><0> ), .B(n4873), .Y(n3898) );
  INVX1 U3727 ( .A(n3898), .Y(n3899) );
  INVX1 U3728 ( .A(n3900), .Y(n3901) );
  AND2X2 U3729 ( .A(\mem<10><0> ), .B(n6399), .Y(n3902) );
  INVX1 U3730 ( .A(n3902), .Y(n3903) );
  AND2X2 U3731 ( .A(\mem<10><1> ), .B(n6399), .Y(n3904) );
  INVX1 U3732 ( .A(n3904), .Y(n3905) );
  AND2X2 U3733 ( .A(\mem<51><1> ), .B(n4873), .Y(n3906) );
  INVX1 U3734 ( .A(n3906), .Y(n3907) );
  AND2X2 U3735 ( .A(n3851), .B(n5250), .Y(n3908) );
  INVX1 U3736 ( .A(n3908), .Y(n3909) );
  AND2X2 U3737 ( .A(\mem<55><1> ), .B(n4873), .Y(n3910) );
  INVX1 U3738 ( .A(n3910), .Y(n3911) );
  AND2X2 U3739 ( .A(\mem<53><1> ), .B(n4873), .Y(n3912) );
  INVX1 U3740 ( .A(n3912), .Y(n3913) );
  AND2X2 U3741 ( .A(\mem<54><1> ), .B(n4873), .Y(n3914) );
  INVX1 U3742 ( .A(n3914), .Y(n3915) );
  AND2X2 U3743 ( .A(\mem<51><2> ), .B(n4873), .Y(n3916) );
  INVX1 U3744 ( .A(n3916), .Y(n3917) );
  AND2X2 U3745 ( .A(n5310), .B(n3851), .Y(n3918) );
  INVX1 U3746 ( .A(n3918), .Y(n3919) );
  AND2X2 U3747 ( .A(\mem<53><2> ), .B(n4873), .Y(n3920) );
  INVX1 U3748 ( .A(n3920), .Y(n3921) );
  AND2X2 U3749 ( .A(n114), .B(n5398), .Y(n3922) );
  INVX1 U3750 ( .A(n3922), .Y(n3923) );
  AND2X2 U3751 ( .A(n3671), .B(\mem<40><3> ), .Y(n3924) );
  INVX1 U3752 ( .A(n3924), .Y(n3925) );
  AND2X2 U3753 ( .A(\mem<51><4> ), .B(n4873), .Y(n3926) );
  INVX1 U3754 ( .A(n3926), .Y(n3927) );
  AND2X2 U3755 ( .A(n3851), .B(n5482), .Y(n3928) );
  INVX1 U3756 ( .A(n3928), .Y(n3929) );
  AND2X2 U3757 ( .A(\mem<53><4> ), .B(n4873), .Y(n3930) );
  INVX1 U3758 ( .A(n3930), .Y(n3931) );
  AND2X2 U3759 ( .A(\mem<40><4> ), .B(n3672), .Y(n3932) );
  INVX1 U3760 ( .A(n3932), .Y(n3933) );
  AND2X2 U3761 ( .A(\mem<51><5> ), .B(n4873), .Y(n3934) );
  INVX1 U3762 ( .A(n3934), .Y(n3935) );
  AND2X2 U3763 ( .A(n3851), .B(n5565), .Y(n3936) );
  INVX1 U3764 ( .A(n3936), .Y(n3937) );
  AND2X2 U3765 ( .A(\mem<53><5> ), .B(n4873), .Y(n3938) );
  INVX1 U3766 ( .A(n3938), .Y(n3939) );
  AND2X2 U3767 ( .A(n3851), .B(n5647), .Y(n3940) );
  INVX1 U3768 ( .A(n3940), .Y(n3941) );
  INVX1 U3769 ( .A(n3942), .Y(n3943) );
  INVX1 U3770 ( .A(n3944), .Y(n3945) );
  AND2X2 U3771 ( .A(\mem<40><7> ), .B(n3672), .Y(n3946) );
  INVX1 U3772 ( .A(n3946), .Y(n3947) );
  AND2X2 U3773 ( .A(n6157), .B(n99), .Y(n3948) );
  INVX1 U3774 ( .A(n3948), .Y(n3949) );
  AND2X2 U3775 ( .A(\mem<6><7> ), .B(n80), .Y(n3950) );
  INVX1 U3776 ( .A(n3950), .Y(n3951) );
  INVX1 U3777 ( .A(\addr<9> ), .Y(n3952) );
  INVX1 U3778 ( .A(\addr<10> ), .Y(n3953) );
  AND2X2 U3779 ( .A(n57), .B(\addr<7> ), .Y(n3954) );
  INVX1 U3780 ( .A(n3954), .Y(n3955) );
  AND2X2 U3781 ( .A(n4964), .B(n720), .Y(n3956) );
  INVX1 U3782 ( .A(n3956), .Y(n3957) );
  AND2X2 U3783 ( .A(\mem<14><7> ), .B(n3847), .Y(n3958) );
  INVX1 U3784 ( .A(n3958), .Y(n3959) );
  AND2X2 U3785 ( .A(\mem<62><0> ), .B(n4919), .Y(n3960) );
  INVX1 U3786 ( .A(n3960), .Y(n3961) );
  AND2X2 U3787 ( .A(\mem<62><1> ), .B(n4919), .Y(n3962) );
  INVX1 U3788 ( .A(n3962), .Y(n3963) );
  AND2X2 U3789 ( .A(\mem<62><2> ), .B(n4919), .Y(n3964) );
  INVX1 U3790 ( .A(n3964), .Y(n3965) );
  AND2X2 U3791 ( .A(\mem<62><3> ), .B(n4919), .Y(n3966) );
  INVX1 U3792 ( .A(n3966), .Y(n3967) );
  AND2X2 U3793 ( .A(\mem<62><4> ), .B(n4919), .Y(n3968) );
  INVX1 U3794 ( .A(n3968), .Y(n3969) );
  AND2X2 U3795 ( .A(\mem<62><5> ), .B(n4919), .Y(n3970) );
  INVX1 U3796 ( .A(n3970), .Y(n3971) );
  AND2X2 U3797 ( .A(\mem<62><6> ), .B(n4919), .Y(n3972) );
  INVX1 U3798 ( .A(n3972), .Y(n3973) );
  AND2X2 U3799 ( .A(\mem<62><7> ), .B(n4919), .Y(n3974) );
  INVX1 U3800 ( .A(n3974), .Y(n3975) );
  AND2X2 U3801 ( .A(\mem<61><0> ), .B(n4920), .Y(n3976) );
  INVX1 U3802 ( .A(n3976), .Y(n3977) );
  AND2X2 U3803 ( .A(\mem<61><1> ), .B(n4920), .Y(n3978) );
  INVX1 U3804 ( .A(n3978), .Y(n3979) );
  AND2X2 U3805 ( .A(\mem<61><2> ), .B(n4920), .Y(n3980) );
  INVX1 U3806 ( .A(n3980), .Y(n3981) );
  AND2X2 U3807 ( .A(\mem<61><3> ), .B(n4920), .Y(n3982) );
  INVX1 U3808 ( .A(n3982), .Y(n3983) );
  AND2X2 U3809 ( .A(\mem<61><4> ), .B(n4920), .Y(n3984) );
  INVX1 U3810 ( .A(n3984), .Y(n3985) );
  AND2X2 U3811 ( .A(\mem<61><5> ), .B(n4920), .Y(n3986) );
  INVX1 U3812 ( .A(n3986), .Y(n3987) );
  AND2X2 U3813 ( .A(\mem<61><6> ), .B(n4920), .Y(n3988) );
  INVX1 U3814 ( .A(n3988), .Y(n3989) );
  AND2X2 U3815 ( .A(\mem<61><7> ), .B(n4920), .Y(n3990) );
  INVX1 U3816 ( .A(n3990), .Y(n3991) );
  AND2X2 U3817 ( .A(n5039), .B(n1692), .Y(n3992) );
  INVX1 U3818 ( .A(n3992), .Y(n3993) );
  AND2X2 U3819 ( .A(n1692), .B(n5045), .Y(n3994) );
  INVX1 U3820 ( .A(n3994), .Y(n3995) );
  AND2X2 U3821 ( .A(n1692), .B(n5053), .Y(n3996) );
  INVX1 U3822 ( .A(n3996), .Y(n3997) );
  AND2X2 U3823 ( .A(n1692), .B(n5057), .Y(n3998) );
  INVX1 U3824 ( .A(n3998), .Y(n3999) );
  AND2X2 U3825 ( .A(n1692), .B(n5066), .Y(n4000) );
  INVX1 U3826 ( .A(n4000), .Y(n4001) );
  AND2X2 U3827 ( .A(n1692), .B(n5070), .Y(n4002) );
  INVX1 U3828 ( .A(n4002), .Y(n4003) );
  INVX1 U3829 ( .A(n876), .Y(n4004) );
  INVX1 U3830 ( .A(n909), .Y(n4005) );
  AND2X2 U3831 ( .A(\mem<28><0> ), .B(n4933), .Y(n4006) );
  INVX1 U3832 ( .A(n4006), .Y(n4007) );
  AND2X2 U3833 ( .A(\mem<28><1> ), .B(n4933), .Y(n4008) );
  INVX1 U3834 ( .A(n4008), .Y(n4009) );
  AND2X2 U3835 ( .A(\mem<28><2> ), .B(n4933), .Y(n4010) );
  INVX1 U3836 ( .A(n4010), .Y(n4011) );
  AND2X2 U3837 ( .A(\mem<28><3> ), .B(n4933), .Y(n4012) );
  INVX1 U3838 ( .A(n4012), .Y(n4013) );
  AND2X2 U3839 ( .A(\mem<28><4> ), .B(n4933), .Y(n4014) );
  INVX1 U3840 ( .A(n4014), .Y(n4015) );
  AND2X2 U3841 ( .A(\mem<28><5> ), .B(n4933), .Y(n4016) );
  INVX1 U3842 ( .A(n4016), .Y(n4017) );
  AND2X2 U3843 ( .A(\mem<28><6> ), .B(n4933), .Y(n4018) );
  INVX1 U3844 ( .A(n4018), .Y(n4019) );
  AND2X2 U3845 ( .A(\mem<28><7> ), .B(n4933), .Y(n4020) );
  INVX1 U3846 ( .A(n4020), .Y(n4021) );
  BUFX2 U3847 ( .A(n6362), .Y(n4933) );
  AND2X2 U3848 ( .A(n5038), .B(n20), .Y(n4022) );
  INVX1 U3849 ( .A(n4022), .Y(n4023) );
  AND2X2 U3850 ( .A(n5043), .B(n1757), .Y(n4024) );
  INVX1 U3851 ( .A(n4024), .Y(n4025) );
  INVX1 U3852 ( .A(n4027), .Y(n4026) );
  AND2X2 U3853 ( .A(n5049), .B(n1757), .Y(n4027) );
  AND2X2 U3854 ( .A(n5053), .B(n20), .Y(n4028) );
  INVX1 U3855 ( .A(n4028), .Y(n4029) );
  AND2X2 U3856 ( .A(n5055), .B(n20), .Y(n4030) );
  INVX1 U3857 ( .A(n4030), .Y(n4031) );
  AND2X2 U3858 ( .A(n5060), .B(n1757), .Y(n4032) );
  INVX1 U3859 ( .A(n4032), .Y(n4033) );
  AND2X2 U3860 ( .A(n5065), .B(n1757), .Y(n4034) );
  INVX1 U3861 ( .A(n4034), .Y(n4035) );
  AND2X2 U3862 ( .A(n5069), .B(n20), .Y(n4036) );
  INVX1 U3863 ( .A(n4036), .Y(n4037) );
  AND2X2 U3864 ( .A(n5038), .B(n1759), .Y(n4038) );
  INVX1 U3865 ( .A(n4038), .Y(n4039) );
  AND2X2 U3866 ( .A(n5042), .B(n1759), .Y(n4040) );
  INVX1 U3867 ( .A(n4040), .Y(n4041) );
  AND2X2 U3868 ( .A(n5048), .B(n1759), .Y(n4042) );
  INVX1 U3869 ( .A(n4042), .Y(n4043) );
  AND2X2 U3870 ( .A(n5052), .B(n1759), .Y(n4044) );
  INVX1 U3871 ( .A(n4044), .Y(n4045) );
  AND2X2 U3872 ( .A(n5056), .B(n1759), .Y(n4046) );
  INVX1 U3873 ( .A(n4046), .Y(n4047) );
  AND2X2 U3874 ( .A(n5060), .B(n1759), .Y(n4048) );
  INVX1 U3875 ( .A(n4048), .Y(n4049) );
  INVX1 U3876 ( .A(n4051), .Y(n4050) );
  AND2X2 U3877 ( .A(n5065), .B(n1759), .Y(n4051) );
  AND2X2 U3878 ( .A(n5069), .B(n1759), .Y(n4052) );
  INVX1 U3879 ( .A(n4052), .Y(n4053) );
  INVX1 U3880 ( .A(n6293), .Y(n6290) );
  OR2X2 U3881 ( .A(n1247), .B(n5175), .Y(n4054) );
  INVX1 U3882 ( .A(n4054), .Y(n4055) );
  OR2X2 U3883 ( .A(n1248), .B(n5279), .Y(n4056) );
  INVX1 U3884 ( .A(n4056), .Y(n4057) );
  OR2X2 U3885 ( .A(n1249), .B(n5341), .Y(n4058) );
  INVX1 U3886 ( .A(n4058), .Y(n4059) );
  INVX1 U3887 ( .A(n5352), .Y(n4060) );
  INVX1 U3888 ( .A(n4060), .Y(n4061) );
  AND2X2 U3889 ( .A(n4897), .B(n5172), .Y(n4062) );
  INVX1 U3890 ( .A(n4062), .Y(n4063) );
  AND2X2 U3891 ( .A(n4891), .B(n5338), .Y(n4064) );
  INVX1 U3892 ( .A(n4064), .Y(n4065) );
  OR2X2 U3893 ( .A(n5526), .B(n5525), .Y(n4066) );
  OR2X2 U3894 ( .A(n5693), .B(n5694), .Y(n4067) );
  AND2X2 U3895 ( .A(n4966), .B(n1060), .Y(n4068) );
  INVX1 U3896 ( .A(n4068), .Y(n4069) );
  AND2X2 U3897 ( .A(\mem<46><7> ), .B(n146), .Y(n4070) );
  INVX1 U3898 ( .A(n4070), .Y(n4071) );
  AND2X2 U3899 ( .A(n5072), .B(n1693), .Y(n4072) );
  INVX1 U3900 ( .A(n4072), .Y(n4073) );
  AND2X2 U3901 ( .A(n5078), .B(n5), .Y(n4074) );
  INVX1 U3902 ( .A(n4074), .Y(n4075) );
  AND2X2 U3903 ( .A(n5084), .B(n5), .Y(n4076) );
  INVX1 U3904 ( .A(n4076), .Y(n4077) );
  AND2X2 U3905 ( .A(n5089), .B(n5), .Y(n4078) );
  INVX1 U3906 ( .A(n4078), .Y(n4079) );
  AND2X2 U3907 ( .A(n5095), .B(n5), .Y(n4080) );
  INVX1 U3908 ( .A(n4080), .Y(n4081) );
  AND2X2 U3909 ( .A(n5099), .B(n1693), .Y(n4082) );
  INVX1 U3910 ( .A(n4082), .Y(n4083) );
  AND2X2 U3911 ( .A(n5103), .B(n1693), .Y(n4084) );
  INVX1 U3912 ( .A(n4084), .Y(n4085) );
  AND2X2 U3913 ( .A(n5107), .B(n1693), .Y(n4086) );
  INVX1 U3914 ( .A(n4086), .Y(n4087) );
  INVX1 U3915 ( .A(n4089), .Y(n4088) );
  AND2X2 U3916 ( .A(n5074), .B(n1701), .Y(n4089) );
  INVX1 U3917 ( .A(n4091), .Y(n4090) );
  AND2X2 U3918 ( .A(n5078), .B(n1701), .Y(n4091) );
  AND2X2 U3919 ( .A(n5084), .B(n1701), .Y(n4092) );
  INVX1 U3920 ( .A(n4092), .Y(n4093) );
  AND2X2 U3921 ( .A(n5089), .B(n1701), .Y(n4094) );
  INVX1 U3922 ( .A(n4094), .Y(n4095) );
  AND2X2 U3923 ( .A(n5095), .B(n1701), .Y(n4096) );
  INVX1 U3924 ( .A(n4096), .Y(n4097) );
  AND2X2 U3925 ( .A(n5099), .B(n1701), .Y(n4098) );
  INVX1 U3926 ( .A(n4098), .Y(n4099) );
  AND2X2 U3927 ( .A(n5103), .B(n1701), .Y(n4100) );
  INVX1 U3928 ( .A(n4100), .Y(n4101) );
  AND2X2 U3929 ( .A(n5108), .B(n1701), .Y(n4102) );
  INVX1 U3930 ( .A(n4102), .Y(n4103) );
  AND2X2 U3931 ( .A(n5074), .B(n1758), .Y(n4104) );
  INVX1 U3932 ( .A(n4104), .Y(n4105) );
  AND2X2 U3933 ( .A(n1758), .B(n5078), .Y(n4106) );
  INVX1 U3934 ( .A(n4106), .Y(n4107) );
  AND2X2 U3935 ( .A(n1758), .B(n5083), .Y(n4108) );
  INVX1 U3936 ( .A(n4108), .Y(n4109) );
  AND2X2 U3937 ( .A(n1758), .B(n5088), .Y(n4110) );
  INVX1 U3938 ( .A(n4110), .Y(n4111) );
  AND2X2 U3939 ( .A(n1758), .B(n5096), .Y(n4112) );
  INVX1 U3940 ( .A(n4112), .Y(n4113) );
  AND2X2 U3941 ( .A(n1758), .B(n5099), .Y(n4114) );
  INVX1 U3942 ( .A(n4114), .Y(n4115) );
  AND2X2 U3943 ( .A(n1758), .B(n5103), .Y(n4116) );
  INVX1 U3944 ( .A(n4116), .Y(n4117) );
  AND2X2 U3945 ( .A(n5108), .B(n1758), .Y(n4118) );
  INVX1 U3946 ( .A(n4118), .Y(n4119) );
  OR2X2 U3947 ( .A(n5386), .B(n5385), .Y(n4120) );
  INVX1 U3948 ( .A(n4120), .Y(n4121) );
  OR2X2 U3949 ( .A(n5447), .B(n5446), .Y(n4122) );
  AND2X2 U3950 ( .A(\mem<6><4> ), .B(n80), .Y(n4123) );
  AND2X2 U3951 ( .A(\mem<6><5> ), .B(n80), .Y(n4124) );
  AND2X2 U3952 ( .A(\mem<6><6> ), .B(n4838), .Y(n4125) );
  AND2X2 U3953 ( .A(\mem<58><0> ), .B(n4923), .Y(n4126) );
  INVX1 U3954 ( .A(n4126), .Y(n4127) );
  AND2X2 U3955 ( .A(\mem<58><1> ), .B(n4923), .Y(n4128) );
  INVX1 U3956 ( .A(n4128), .Y(n4129) );
  AND2X2 U3957 ( .A(\mem<58><2> ), .B(n4923), .Y(n4130) );
  INVX1 U3958 ( .A(n4130), .Y(n4131) );
  AND2X2 U3959 ( .A(\mem<58><3> ), .B(n4923), .Y(n4132) );
  INVX1 U3960 ( .A(n4132), .Y(n4133) );
  AND2X2 U3961 ( .A(\mem<58><4> ), .B(n4923), .Y(n4134) );
  INVX1 U3962 ( .A(n4134), .Y(n4135) );
  AND2X2 U3963 ( .A(\mem<58><5> ), .B(n4923), .Y(n4136) );
  INVX1 U3964 ( .A(n4136), .Y(n4137) );
  AND2X2 U3965 ( .A(\mem<58><6> ), .B(n4923), .Y(n4138) );
  INVX1 U3966 ( .A(n4138), .Y(n4139) );
  AND2X2 U3967 ( .A(\mem<58><7> ), .B(n4923), .Y(n4140) );
  INVX1 U3968 ( .A(n4140), .Y(n4141) );
  AND2X2 U3969 ( .A(\mem<54><0> ), .B(n4924), .Y(n4142) );
  INVX1 U3970 ( .A(n4142), .Y(n4143) );
  AND2X2 U3971 ( .A(\mem<54><1> ), .B(n4924), .Y(n4144) );
  INVX1 U3972 ( .A(n4144), .Y(n4145) );
  AND2X2 U3973 ( .A(\mem<54><2> ), .B(n4924), .Y(n4146) );
  INVX1 U3974 ( .A(n4146), .Y(n4147) );
  AND2X2 U3975 ( .A(\mem<54><3> ), .B(n4924), .Y(n4148) );
  INVX1 U3976 ( .A(n4148), .Y(n4149) );
  AND2X2 U3977 ( .A(\mem<54><4> ), .B(n4924), .Y(n4150) );
  INVX1 U3978 ( .A(n4150), .Y(n4151) );
  AND2X2 U3979 ( .A(\mem<54><5> ), .B(n4924), .Y(n4152) );
  INVX1 U3980 ( .A(n4152), .Y(n4153) );
  AND2X2 U3981 ( .A(\mem<54><6> ), .B(n4924), .Y(n4154) );
  INVX1 U3982 ( .A(n4154), .Y(n4155) );
  AND2X2 U3983 ( .A(\mem<54><7> ), .B(n4924), .Y(n4156) );
  INVX1 U3984 ( .A(n4156), .Y(n4157) );
  AND2X2 U3985 ( .A(\mem<53><0> ), .B(n4925), .Y(n4158) );
  INVX1 U3986 ( .A(n4158), .Y(n4159) );
  AND2X2 U3987 ( .A(\mem<53><1> ), .B(n4925), .Y(n4160) );
  INVX1 U3988 ( .A(n4160), .Y(n4161) );
  AND2X2 U3989 ( .A(\mem<53><2> ), .B(n4925), .Y(n4162) );
  INVX1 U3990 ( .A(n4162), .Y(n4163) );
  AND2X2 U3991 ( .A(\mem<53><3> ), .B(n4925), .Y(n4164) );
  INVX1 U3992 ( .A(n4164), .Y(n4165) );
  AND2X2 U3993 ( .A(\mem<53><4> ), .B(n4925), .Y(n4166) );
  INVX1 U3994 ( .A(n4166), .Y(n4167) );
  AND2X2 U3995 ( .A(\mem<53><5> ), .B(n4925), .Y(n4168) );
  INVX1 U3996 ( .A(n4168), .Y(n4169) );
  AND2X2 U3997 ( .A(\mem<53><6> ), .B(n4925), .Y(n4170) );
  INVX1 U3998 ( .A(n4170), .Y(n4171) );
  AND2X2 U3999 ( .A(\mem<53><7> ), .B(n4925), .Y(n4172) );
  INVX1 U4000 ( .A(n4172), .Y(n4173) );
  AND2X2 U4001 ( .A(\mem<50><0> ), .B(n3590), .Y(n4174) );
  INVX1 U4002 ( .A(n4174), .Y(n4175) );
  AND2X2 U4003 ( .A(\mem<50><1> ), .B(n3590), .Y(n4176) );
  INVX1 U4004 ( .A(n4176), .Y(n4177) );
  AND2X2 U4005 ( .A(\mem<50><2> ), .B(n3590), .Y(n4178) );
  INVX1 U4006 ( .A(n4178), .Y(n4179) );
  AND2X2 U4007 ( .A(\mem<50><3> ), .B(n3590), .Y(n4180) );
  INVX1 U4008 ( .A(n4180), .Y(n4181) );
  AND2X2 U4009 ( .A(\mem<50><4> ), .B(n3590), .Y(n4182) );
  INVX1 U4010 ( .A(n4182), .Y(n4183) );
  AND2X2 U4011 ( .A(\mem<50><5> ), .B(n3590), .Y(n4184) );
  INVX1 U4012 ( .A(n4184), .Y(n4185) );
  AND2X2 U4013 ( .A(\mem<50><6> ), .B(n3590), .Y(n4186) );
  INVX1 U4014 ( .A(n4186), .Y(n4187) );
  AND2X2 U4015 ( .A(\mem<50><7> ), .B(n3590), .Y(n4188) );
  INVX1 U4016 ( .A(n4188), .Y(n4189) );
  AND2X2 U4017 ( .A(\mem<46><0> ), .B(n4926), .Y(n4190) );
  INVX1 U4018 ( .A(n4190), .Y(n4191) );
  AND2X2 U4019 ( .A(\mem<46><1> ), .B(n4926), .Y(n4192) );
  INVX1 U4020 ( .A(n4192), .Y(n4193) );
  AND2X2 U4021 ( .A(\mem<46><2> ), .B(n4926), .Y(n4194) );
  INVX1 U4022 ( .A(n4194), .Y(n4195) );
  AND2X2 U4023 ( .A(\mem<46><3> ), .B(n4926), .Y(n4196) );
  INVX1 U4024 ( .A(n4196), .Y(n4197) );
  AND2X2 U4025 ( .A(\mem<46><4> ), .B(n4926), .Y(n4198) );
  INVX1 U4026 ( .A(n4198), .Y(n4199) );
  AND2X2 U4027 ( .A(\mem<46><5> ), .B(n4926), .Y(n4200) );
  INVX1 U4028 ( .A(n4200), .Y(n4201) );
  AND2X2 U4029 ( .A(\mem<46><6> ), .B(n4926), .Y(n4202) );
  INVX1 U4030 ( .A(n4202), .Y(n4203) );
  AND2X2 U4031 ( .A(\mem<46><7> ), .B(n4926), .Y(n4204) );
  INVX1 U4032 ( .A(n4204), .Y(n4205) );
  AND2X2 U4033 ( .A(n6329), .B(\mem<45><0> ), .Y(n4206) );
  INVX1 U4034 ( .A(n4206), .Y(n4207) );
  AND2X2 U4035 ( .A(n6329), .B(\mem<45><1> ), .Y(n4208) );
  INVX1 U4036 ( .A(n4208), .Y(n4209) );
  AND2X2 U4037 ( .A(n6329), .B(\mem<45><2> ), .Y(n4210) );
  INVX1 U4038 ( .A(n4210), .Y(n4211) );
  AND2X2 U4039 ( .A(n6329), .B(\mem<45><3> ), .Y(n4212) );
  INVX1 U4040 ( .A(n4212), .Y(n4213) );
  AND2X2 U4041 ( .A(\mem<45><4> ), .B(n27), .Y(n4214) );
  INVX1 U4042 ( .A(n4214), .Y(n4215) );
  AND2X2 U4043 ( .A(\mem<45><5> ), .B(n27), .Y(n4216) );
  INVX1 U4044 ( .A(n4216), .Y(n4217) );
  AND2X2 U4045 ( .A(\mem<45><6> ), .B(n27), .Y(n4218) );
  INVX1 U4046 ( .A(n4218), .Y(n4219) );
  AND2X2 U4047 ( .A(n6329), .B(\mem<45><7> ), .Y(n4220) );
  INVX1 U4048 ( .A(n4220), .Y(n4221) );
  AND2X2 U4049 ( .A(\mem<44><0> ), .B(n3598), .Y(n4222) );
  INVX1 U4050 ( .A(n4222), .Y(n4223) );
  AND2X2 U4051 ( .A(\mem<44><1> ), .B(n3598), .Y(n4224) );
  INVX1 U4052 ( .A(n4224), .Y(n4225) );
  AND2X2 U4053 ( .A(\mem<44><2> ), .B(n3598), .Y(n4226) );
  INVX1 U4054 ( .A(n4226), .Y(n4227) );
  AND2X2 U4055 ( .A(\mem<44><3> ), .B(n3598), .Y(n4228) );
  INVX1 U4056 ( .A(n4228), .Y(n4229) );
  AND2X2 U4057 ( .A(\mem<44><4> ), .B(n3598), .Y(n4230) );
  INVX1 U4058 ( .A(n4230), .Y(n4231) );
  AND2X2 U4059 ( .A(\mem<44><5> ), .B(n3598), .Y(n4232) );
  INVX1 U4060 ( .A(n4232), .Y(n4233) );
  AND2X2 U4061 ( .A(\mem<44><6> ), .B(n3598), .Y(n4234) );
  INVX1 U4062 ( .A(n4234), .Y(n4235) );
  AND2X2 U4063 ( .A(\mem<44><7> ), .B(n3598), .Y(n4236) );
  INVX1 U4064 ( .A(n4236), .Y(n4237) );
  AND2X2 U4065 ( .A(\mem<43><0> ), .B(n3600), .Y(n4238) );
  INVX1 U4066 ( .A(n4238), .Y(n4239) );
  AND2X2 U4067 ( .A(\mem<43><1> ), .B(n3600), .Y(n4240) );
  INVX1 U4068 ( .A(n4240), .Y(n4241) );
  AND2X2 U4069 ( .A(\mem<43><2> ), .B(n3600), .Y(n4242) );
  INVX1 U4070 ( .A(n4242), .Y(n4243) );
  AND2X2 U4071 ( .A(\mem<43><3> ), .B(n3600), .Y(n4244) );
  INVX1 U4072 ( .A(n4244), .Y(n4245) );
  AND2X2 U4073 ( .A(\mem<43><4> ), .B(n3600), .Y(n4246) );
  INVX1 U4074 ( .A(n4246), .Y(n4247) );
  AND2X2 U4075 ( .A(\mem<43><5> ), .B(n3600), .Y(n4248) );
  INVX1 U4076 ( .A(n4248), .Y(n4249) );
  AND2X2 U4077 ( .A(\mem<43><6> ), .B(n3600), .Y(n4250) );
  INVX1 U4078 ( .A(n4250), .Y(n4251) );
  AND2X2 U4079 ( .A(\mem<43><7> ), .B(n3600), .Y(n4252) );
  INVX1 U4080 ( .A(n4252), .Y(n4253) );
  AND2X2 U4081 ( .A(\mem<42><0> ), .B(n3602), .Y(n4254) );
  INVX1 U4082 ( .A(n4254), .Y(n4255) );
  AND2X2 U4083 ( .A(\mem<42><1> ), .B(n3602), .Y(n4256) );
  INVX1 U4084 ( .A(n4256), .Y(n4257) );
  AND2X2 U4085 ( .A(\mem<42><2> ), .B(n3602), .Y(n4258) );
  INVX1 U4086 ( .A(n4258), .Y(n4259) );
  AND2X2 U4087 ( .A(\mem<42><3> ), .B(n3602), .Y(n4260) );
  INVX1 U4088 ( .A(n4260), .Y(n4261) );
  AND2X2 U4089 ( .A(\mem<42><4> ), .B(n3602), .Y(n4262) );
  INVX1 U4090 ( .A(n4262), .Y(n4263) );
  AND2X2 U4091 ( .A(\mem<42><5> ), .B(n3602), .Y(n4264) );
  INVX1 U4092 ( .A(n4264), .Y(n4265) );
  AND2X2 U4093 ( .A(\mem<42><6> ), .B(n3602), .Y(n4266) );
  INVX1 U4094 ( .A(n4266), .Y(n4267) );
  AND2X2 U4095 ( .A(\mem<42><7> ), .B(n3602), .Y(n4268) );
  INVX1 U4096 ( .A(n4268), .Y(n4269) );
  AND2X2 U4097 ( .A(\mem<40><0> ), .B(n3606), .Y(n4270) );
  INVX1 U4098 ( .A(n4270), .Y(n4271) );
  AND2X2 U4099 ( .A(\mem<40><1> ), .B(n3606), .Y(n4272) );
  INVX1 U4100 ( .A(n4272), .Y(n4273) );
  AND2X2 U4101 ( .A(\mem<40><2> ), .B(n3606), .Y(n4274) );
  INVX1 U4102 ( .A(n4274), .Y(n4275) );
  AND2X2 U4103 ( .A(\mem<40><3> ), .B(n3606), .Y(n4276) );
  INVX1 U4104 ( .A(n4276), .Y(n4277) );
  AND2X2 U4105 ( .A(\mem<40><4> ), .B(n3606), .Y(n4278) );
  INVX1 U4106 ( .A(n4278), .Y(n4279) );
  AND2X2 U4107 ( .A(\mem<40><5> ), .B(n3606), .Y(n4280) );
  INVX1 U4108 ( .A(n4280), .Y(n4281) );
  AND2X2 U4109 ( .A(\mem<40><6> ), .B(n3606), .Y(n4282) );
  INVX1 U4110 ( .A(n4282), .Y(n4283) );
  AND2X2 U4111 ( .A(\mem<40><7> ), .B(n3606), .Y(n4284) );
  INVX1 U4112 ( .A(n4284), .Y(n4285) );
  AND2X2 U4113 ( .A(\mem<39><0> ), .B(n3608), .Y(n4286) );
  INVX1 U4114 ( .A(n4286), .Y(n4287) );
  AND2X2 U4115 ( .A(\mem<39><1> ), .B(n3608), .Y(n4288) );
  INVX1 U4116 ( .A(n4288), .Y(n4289) );
  AND2X2 U4117 ( .A(\mem<39><2> ), .B(n3608), .Y(n4290) );
  INVX1 U4118 ( .A(n4290), .Y(n4291) );
  AND2X2 U4119 ( .A(\mem<39><3> ), .B(n3608), .Y(n4292) );
  INVX1 U4120 ( .A(n4292), .Y(n4293) );
  AND2X2 U4121 ( .A(\mem<39><4> ), .B(n3608), .Y(n4294) );
  INVX1 U4122 ( .A(n4294), .Y(n4295) );
  AND2X2 U4123 ( .A(\mem<39><5> ), .B(n3608), .Y(n4296) );
  INVX1 U4124 ( .A(n4296), .Y(n4297) );
  AND2X2 U4125 ( .A(\mem<39><6> ), .B(n3608), .Y(n4298) );
  INVX1 U4126 ( .A(n4298), .Y(n4299) );
  AND2X2 U4127 ( .A(\mem<39><7> ), .B(n3608), .Y(n4300) );
  INVX1 U4128 ( .A(n4300), .Y(n4301) );
  AND2X2 U4129 ( .A(\mem<38><0> ), .B(n4927), .Y(n4302) );
  INVX1 U4130 ( .A(n4302), .Y(n4303) );
  AND2X2 U4131 ( .A(\mem<38><1> ), .B(n4927), .Y(n4304) );
  INVX1 U4132 ( .A(n4304), .Y(n4305) );
  AND2X2 U4133 ( .A(\mem<38><2> ), .B(n4927), .Y(n4306) );
  INVX1 U4134 ( .A(n4306), .Y(n4307) );
  AND2X2 U4135 ( .A(\mem<38><3> ), .B(n4927), .Y(n4308) );
  INVX1 U4136 ( .A(n4308), .Y(n4309) );
  AND2X2 U4137 ( .A(\mem<38><4> ), .B(n4927), .Y(n4310) );
  INVX1 U4138 ( .A(n4310), .Y(n4311) );
  AND2X2 U4139 ( .A(\mem<38><5> ), .B(n4927), .Y(n4312) );
  INVX1 U4140 ( .A(n4312), .Y(n4313) );
  AND2X2 U4141 ( .A(\mem<38><6> ), .B(n4927), .Y(n4314) );
  INVX1 U4142 ( .A(n4314), .Y(n4315) );
  AND2X2 U4143 ( .A(\mem<38><7> ), .B(n4927), .Y(n4316) );
  INVX1 U4144 ( .A(n4316), .Y(n4317) );
  AND2X2 U4145 ( .A(\mem<37><0> ), .B(n4928), .Y(n4318) );
  INVX1 U4146 ( .A(n4318), .Y(n4319) );
  AND2X2 U4147 ( .A(\mem<37><1> ), .B(n4928), .Y(n4320) );
  INVX1 U4148 ( .A(n4320), .Y(n4321) );
  AND2X2 U4149 ( .A(\mem<37><2> ), .B(n4928), .Y(n4322) );
  INVX1 U4150 ( .A(n4322), .Y(n4323) );
  AND2X2 U4151 ( .A(\mem<37><3> ), .B(n4928), .Y(n4324) );
  INVX1 U4152 ( .A(n4324), .Y(n4325) );
  AND2X2 U4153 ( .A(\mem<37><4> ), .B(n4928), .Y(n4326) );
  INVX1 U4154 ( .A(n4326), .Y(n4327) );
  AND2X2 U4155 ( .A(\mem<37><5> ), .B(n4928), .Y(n4328) );
  INVX1 U4156 ( .A(n4328), .Y(n4329) );
  AND2X2 U4157 ( .A(\mem<37><6> ), .B(n4928), .Y(n4330) );
  INVX1 U4158 ( .A(n4330), .Y(n4331) );
  AND2X2 U4159 ( .A(\mem<37><7> ), .B(n4928), .Y(n4332) );
  INVX1 U4160 ( .A(n4332), .Y(n4333) );
  AND2X2 U4161 ( .A(\mem<34><0> ), .B(n3614), .Y(n4334) );
  INVX1 U4162 ( .A(n4334), .Y(n4335) );
  AND2X2 U4163 ( .A(\mem<34><1> ), .B(n3614), .Y(n4336) );
  INVX1 U4164 ( .A(n4336), .Y(n4337) );
  AND2X2 U4165 ( .A(\mem<34><2> ), .B(n3614), .Y(n4338) );
  INVX1 U4166 ( .A(n4338), .Y(n4339) );
  AND2X2 U4167 ( .A(\mem<34><3> ), .B(n3614), .Y(n4340) );
  INVX1 U4168 ( .A(n4340), .Y(n4341) );
  AND2X2 U4169 ( .A(\mem<34><4> ), .B(n3614), .Y(n4342) );
  INVX1 U4170 ( .A(n4342), .Y(n4343) );
  AND2X2 U4171 ( .A(\mem<34><5> ), .B(n3614), .Y(n4344) );
  INVX1 U4172 ( .A(n4344), .Y(n4345) );
  AND2X2 U4173 ( .A(\mem<34><6> ), .B(n3614), .Y(n4346) );
  INVX1 U4174 ( .A(n4346), .Y(n4347) );
  AND2X2 U4175 ( .A(\mem<34><7> ), .B(n3614), .Y(n4348) );
  INVX1 U4176 ( .A(n4348), .Y(n4349) );
  AND2X2 U4177 ( .A(\mem<32><0> ), .B(n4929), .Y(n4350) );
  INVX1 U4178 ( .A(n4350), .Y(n4351) );
  AND2X2 U4179 ( .A(\mem<32><1> ), .B(n4929), .Y(n4352) );
  INVX1 U4180 ( .A(n4352), .Y(n4353) );
  AND2X2 U4181 ( .A(\mem<32><2> ), .B(n4929), .Y(n4354) );
  INVX1 U4182 ( .A(n4354), .Y(n4355) );
  AND2X2 U4183 ( .A(\mem<32><3> ), .B(n4929), .Y(n4356) );
  INVX1 U4184 ( .A(n4356), .Y(n4357) );
  AND2X2 U4185 ( .A(\mem<32><4> ), .B(n4929), .Y(n4358) );
  INVX1 U4186 ( .A(n4358), .Y(n4359) );
  AND2X2 U4187 ( .A(\mem<32><5> ), .B(n4929), .Y(n4360) );
  INVX1 U4188 ( .A(n4360), .Y(n4361) );
  AND2X2 U4189 ( .A(\mem<32><6> ), .B(n4929), .Y(n4362) );
  INVX1 U4190 ( .A(n4362), .Y(n4363) );
  AND2X2 U4191 ( .A(\mem<32><7> ), .B(n4929), .Y(n4364) );
  INVX1 U4192 ( .A(n4364), .Y(n4365) );
  AND2X2 U4193 ( .A(n5038), .B(n4685), .Y(n4366) );
  INVX1 U4194 ( .A(n4366), .Y(n4367) );
  AND2X2 U4195 ( .A(n5043), .B(n94), .Y(n4368) );
  INVX1 U4196 ( .A(n4368), .Y(n4369) );
  AND2X2 U4197 ( .A(n94), .B(n5049), .Y(n4370) );
  INVX1 U4198 ( .A(n4370), .Y(n4371) );
  INVX1 U4199 ( .A(n4373), .Y(n4372) );
  AND2X2 U4200 ( .A(n5053), .B(n94), .Y(n4373) );
  AND2X2 U4201 ( .A(n5056), .B(n4686), .Y(n4374) );
  INVX1 U4202 ( .A(n4374), .Y(n4375) );
  AND2X2 U4203 ( .A(n5060), .B(n4686), .Y(n4376) );
  INVX1 U4204 ( .A(n4376), .Y(n4377) );
  AND2X2 U4205 ( .A(n5065), .B(n4685), .Y(n4378) );
  INVX1 U4206 ( .A(n4378), .Y(n4379) );
  INVX1 U4207 ( .A(n4381), .Y(n4380) );
  AND2X2 U4208 ( .A(n5069), .B(n4685), .Y(n4381) );
  AND2X2 U4209 ( .A(\mem<27><0> ), .B(n24), .Y(n4382) );
  INVX1 U4210 ( .A(n4382), .Y(n4383) );
  AND2X2 U4211 ( .A(\mem<27><1> ), .B(n49), .Y(n4384) );
  INVX1 U4212 ( .A(n4384), .Y(n4385) );
  AND2X2 U4213 ( .A(\mem<27><2> ), .B(n49), .Y(n4386) );
  INVX1 U4214 ( .A(n4386), .Y(n4387) );
  AND2X2 U4215 ( .A(\mem<27><3> ), .B(n49), .Y(n4388) );
  INVX1 U4216 ( .A(n4388), .Y(n4389) );
  AND2X2 U4217 ( .A(n23), .B(\mem<27><4> ), .Y(n4390) );
  INVX1 U4218 ( .A(n4390), .Y(n4391) );
  AND2X2 U4219 ( .A(\mem<27><5> ), .B(n22), .Y(n4392) );
  INVX1 U4220 ( .A(n4392), .Y(n4393) );
  AND2X2 U4221 ( .A(\mem<27><6> ), .B(n23), .Y(n4394) );
  INVX1 U4222 ( .A(n4394), .Y(n4395) );
  AND2X2 U4223 ( .A(\mem<27><7> ), .B(n22), .Y(n4396) );
  INVX1 U4224 ( .A(n4396), .Y(n4397) );
  AND2X2 U4225 ( .A(\mem<22><1> ), .B(n4934), .Y(n4398) );
  INVX1 U4226 ( .A(n4398), .Y(n4399) );
  AND2X2 U4227 ( .A(\mem<22><2> ), .B(n4934), .Y(n4400) );
  INVX1 U4228 ( .A(n4400), .Y(n4401) );
  AND2X2 U4229 ( .A(\mem<22><3> ), .B(n4934), .Y(n4402) );
  INVX1 U4230 ( .A(n4402), .Y(n4403) );
  AND2X2 U4231 ( .A(\mem<22><4> ), .B(n4934), .Y(n4404) );
  INVX1 U4232 ( .A(n4404), .Y(n4405) );
  AND2X2 U4233 ( .A(\mem<22><5> ), .B(n4934), .Y(n4406) );
  INVX1 U4234 ( .A(n4406), .Y(n4407) );
  AND2X2 U4235 ( .A(\mem<22><6> ), .B(n4934), .Y(n4408) );
  INVX1 U4236 ( .A(n4408), .Y(n4409) );
  AND2X2 U4237 ( .A(\mem<22><7> ), .B(n4934), .Y(n4410) );
  INVX1 U4238 ( .A(n4410), .Y(n4411) );
  AND2X2 U4239 ( .A(\mem<21><0> ), .B(n4935), .Y(n4412) );
  INVX1 U4240 ( .A(n4412), .Y(n4413) );
  AND2X2 U4241 ( .A(\mem<21><1> ), .B(n4935), .Y(n4414) );
  INVX1 U4242 ( .A(n4414), .Y(n4415) );
  AND2X2 U4243 ( .A(\mem<21><2> ), .B(n4935), .Y(n4416) );
  INVX1 U4244 ( .A(n4416), .Y(n4417) );
  AND2X2 U4245 ( .A(\mem<21><3> ), .B(n4935), .Y(n4418) );
  INVX1 U4246 ( .A(n4418), .Y(n4419) );
  AND2X2 U4247 ( .A(\mem<21><4> ), .B(n4935), .Y(n4420) );
  INVX1 U4248 ( .A(n4420), .Y(n4421) );
  AND2X2 U4249 ( .A(\mem<21><5> ), .B(n4935), .Y(n4422) );
  INVX1 U4250 ( .A(n4422), .Y(n4423) );
  AND2X2 U4251 ( .A(\mem<21><6> ), .B(n4935), .Y(n4424) );
  INVX1 U4252 ( .A(n4424), .Y(n4425) );
  AND2X2 U4253 ( .A(\mem<21><7> ), .B(n4935), .Y(n4426) );
  INVX1 U4254 ( .A(n4426), .Y(n4427) );
  AND2X2 U4255 ( .A(\mem<18><0> ), .B(n3630), .Y(n4428) );
  INVX1 U4256 ( .A(n4428), .Y(n4429) );
  AND2X2 U4257 ( .A(\mem<18><1> ), .B(n3630), .Y(n4430) );
  INVX1 U4258 ( .A(n4430), .Y(n4431) );
  AND2X2 U4259 ( .A(\mem<18><2> ), .B(n3630), .Y(n4432) );
  INVX1 U4260 ( .A(n4432), .Y(n4433) );
  AND2X2 U4261 ( .A(\mem<18><3> ), .B(n3630), .Y(n4434) );
  INVX1 U4262 ( .A(n4434), .Y(n4435) );
  AND2X2 U4263 ( .A(\mem<18><4> ), .B(n3630), .Y(n4436) );
  INVX1 U4264 ( .A(n4436), .Y(n4437) );
  AND2X2 U4265 ( .A(\mem<18><5> ), .B(n3630), .Y(n4438) );
  INVX1 U4266 ( .A(n4438), .Y(n4439) );
  AND2X2 U4267 ( .A(\mem<18><6> ), .B(n3630), .Y(n4440) );
  INVX1 U4268 ( .A(n4440), .Y(n4441) );
  AND2X2 U4269 ( .A(\mem<18><7> ), .B(n3630), .Y(n4442) );
  INVX1 U4270 ( .A(n4442), .Y(n4443) );
  AND2X2 U4271 ( .A(\mem<17><0> ), .B(n85), .Y(n4444) );
  INVX1 U4272 ( .A(n4444), .Y(n4445) );
  AND2X2 U4273 ( .A(\mem<17><1> ), .B(n11), .Y(n4446) );
  INVX1 U4274 ( .A(n4446), .Y(n4447) );
  AND2X2 U4275 ( .A(\mem<17><2> ), .B(n3632), .Y(n4448) );
  INVX1 U4276 ( .A(n4448), .Y(n4449) );
  AND2X2 U4277 ( .A(\mem<17><3> ), .B(n85), .Y(n4450) );
  INVX1 U4278 ( .A(n4450), .Y(n4451) );
  AND2X2 U4279 ( .A(\mem<17><4> ), .B(n11), .Y(n4452) );
  INVX1 U4280 ( .A(n4452), .Y(n4453) );
  AND2X2 U4281 ( .A(\mem<17><5> ), .B(n3632), .Y(n4454) );
  INVX1 U4282 ( .A(n4454), .Y(n4455) );
  AND2X2 U4283 ( .A(\mem<17><6> ), .B(n85), .Y(n4456) );
  INVX1 U4284 ( .A(n4456), .Y(n4457) );
  AND2X2 U4285 ( .A(\mem<17><7> ), .B(n3632), .Y(n4458) );
  INVX1 U4286 ( .A(n4458), .Y(n4459) );
  AND2X2 U4287 ( .A(\mem<16><0> ), .B(n3848), .Y(n4460) );
  INVX1 U4288 ( .A(n4460), .Y(n4461) );
  AND2X2 U4289 ( .A(\mem<16><1> ), .B(n3848), .Y(n4462) );
  INVX1 U4290 ( .A(n4462), .Y(n4463) );
  AND2X2 U4291 ( .A(\mem<16><2> ), .B(n3848), .Y(n4464) );
  INVX1 U4292 ( .A(n4464), .Y(n4465) );
  AND2X2 U4293 ( .A(\mem<16><3> ), .B(n6389), .Y(n4466) );
  INVX1 U4294 ( .A(n4466), .Y(n4467) );
  AND2X2 U4295 ( .A(\mem<16><4> ), .B(n6389), .Y(n4468) );
  INVX1 U4296 ( .A(n4468), .Y(n4469) );
  AND2X2 U4297 ( .A(\mem<16><5> ), .B(n6389), .Y(n4470) );
  INVX1 U4298 ( .A(n4470), .Y(n4471) );
  AND2X2 U4299 ( .A(\mem<16><6> ), .B(n6389), .Y(n4472) );
  INVX1 U4300 ( .A(n4472), .Y(n4473) );
  AND2X2 U4301 ( .A(\mem<16><7> ), .B(n6389), .Y(n4474) );
  INVX1 U4302 ( .A(n4474), .Y(n4475) );
  AND2X2 U4303 ( .A(\mem<14><0> ), .B(n4936), .Y(n4476) );
  INVX1 U4304 ( .A(n4476), .Y(n4477) );
  AND2X2 U4305 ( .A(\mem<14><1> ), .B(n4936), .Y(n4478) );
  INVX1 U4306 ( .A(n4478), .Y(n4479) );
  AND2X2 U4307 ( .A(\mem<14><2> ), .B(n4936), .Y(n4480) );
  INVX1 U4308 ( .A(n4480), .Y(n4481) );
  AND2X2 U4309 ( .A(\mem<14><3> ), .B(n4936), .Y(n4482) );
  INVX1 U4310 ( .A(n4482), .Y(n4483) );
  AND2X2 U4311 ( .A(\mem<14><4> ), .B(n4936), .Y(n4484) );
  INVX1 U4312 ( .A(n4484), .Y(n4485) );
  AND2X2 U4313 ( .A(\mem<14><5> ), .B(n4936), .Y(n4486) );
  INVX1 U4314 ( .A(n4486), .Y(n4487) );
  AND2X2 U4315 ( .A(\mem<14><6> ), .B(n4936), .Y(n4488) );
  INVX1 U4316 ( .A(n4488), .Y(n4489) );
  AND2X2 U4317 ( .A(\mem<14><7> ), .B(n4936), .Y(n4490) );
  INVX1 U4318 ( .A(n4490), .Y(n4491) );
  AND2X2 U4319 ( .A(\mem<13><0> ), .B(n4937), .Y(n4492) );
  INVX1 U4320 ( .A(n4492), .Y(n4493) );
  AND2X2 U4321 ( .A(\mem<13><1> ), .B(n4937), .Y(n4494) );
  INVX1 U4322 ( .A(n4494), .Y(n4495) );
  AND2X2 U4323 ( .A(\mem<13><2> ), .B(n4937), .Y(n4496) );
  INVX1 U4324 ( .A(n4496), .Y(n4497) );
  AND2X2 U4325 ( .A(\mem<13><3> ), .B(n4937), .Y(n4498) );
  INVX1 U4326 ( .A(n4498), .Y(n4499) );
  AND2X2 U4327 ( .A(\mem<13><4> ), .B(n4937), .Y(n4500) );
  INVX1 U4328 ( .A(n4500), .Y(n4501) );
  AND2X2 U4329 ( .A(\mem<13><5> ), .B(n4937), .Y(n4502) );
  INVX1 U4330 ( .A(n4502), .Y(n4503) );
  AND2X2 U4331 ( .A(\mem<13><6> ), .B(n4937), .Y(n4504) );
  INVX1 U4332 ( .A(n4504), .Y(n4505) );
  AND2X2 U4333 ( .A(\mem<13><7> ), .B(n4937), .Y(n4506) );
  INVX1 U4334 ( .A(n4506), .Y(n4507) );
  AND2X2 U4335 ( .A(\mem<10><0> ), .B(n3636), .Y(n4508) );
  INVX1 U4336 ( .A(n4508), .Y(n4509) );
  AND2X2 U4337 ( .A(\mem<10><1> ), .B(n3636), .Y(n4510) );
  INVX1 U4338 ( .A(n4510), .Y(n4511) );
  AND2X2 U4339 ( .A(\mem<10><2> ), .B(n3636), .Y(n4512) );
  INVX1 U4340 ( .A(n4512), .Y(n4513) );
  AND2X2 U4341 ( .A(\mem<10><3> ), .B(n3636), .Y(n4514) );
  INVX1 U4342 ( .A(n4514), .Y(n4515) );
  AND2X2 U4343 ( .A(\mem<10><4> ), .B(n3636), .Y(n4516) );
  INVX1 U4344 ( .A(n4516), .Y(n4517) );
  AND2X2 U4345 ( .A(\mem<10><5> ), .B(n3636), .Y(n4518) );
  INVX1 U4346 ( .A(n4518), .Y(n4519) );
  AND2X2 U4347 ( .A(\mem<10><6> ), .B(n3636), .Y(n4520) );
  INVX1 U4348 ( .A(n4520), .Y(n4521) );
  AND2X2 U4349 ( .A(\mem<10><7> ), .B(n3636), .Y(n4522) );
  INVX1 U4350 ( .A(n4522), .Y(n4523) );
  AND2X2 U4351 ( .A(\mem<9><0> ), .B(n3638), .Y(n4524) );
  INVX1 U4352 ( .A(n4524), .Y(n4525) );
  AND2X2 U4353 ( .A(\mem<9><1> ), .B(n3638), .Y(n4526) );
  INVX1 U4354 ( .A(n4526), .Y(n4527) );
  AND2X2 U4355 ( .A(\mem<9><2> ), .B(n3638), .Y(n4528) );
  INVX1 U4356 ( .A(n4528), .Y(n4529) );
  AND2X2 U4357 ( .A(\mem<9><3> ), .B(n3638), .Y(n4530) );
  INVX1 U4358 ( .A(n4530), .Y(n4531) );
  AND2X2 U4359 ( .A(\mem<9><4> ), .B(n3638), .Y(n4532) );
  INVX1 U4360 ( .A(n4532), .Y(n4533) );
  AND2X2 U4361 ( .A(\mem<9><5> ), .B(n3638), .Y(n4534) );
  INVX1 U4362 ( .A(n4534), .Y(n4535) );
  AND2X2 U4363 ( .A(\mem<9><6> ), .B(n3638), .Y(n4536) );
  INVX1 U4364 ( .A(n4536), .Y(n4537) );
  AND2X2 U4365 ( .A(\mem<9><7> ), .B(n3638), .Y(n4538) );
  INVX1 U4366 ( .A(n4538), .Y(n4539) );
  AND2X2 U4367 ( .A(\mem<8><0> ), .B(n3640), .Y(n4540) );
  INVX1 U4368 ( .A(n4540), .Y(n4541) );
  AND2X2 U4369 ( .A(\mem<8><1> ), .B(n3640), .Y(n4542) );
  INVX1 U4370 ( .A(n4542), .Y(n4543) );
  AND2X2 U4371 ( .A(\mem<8><2> ), .B(n3640), .Y(n4544) );
  INVX1 U4372 ( .A(n4544), .Y(n4545) );
  AND2X2 U4373 ( .A(\mem<8><3> ), .B(n3640), .Y(n4546) );
  INVX1 U4374 ( .A(n4546), .Y(n4547) );
  AND2X2 U4375 ( .A(\mem<8><4> ), .B(n3640), .Y(n4548) );
  INVX1 U4376 ( .A(n4548), .Y(n4549) );
  AND2X2 U4377 ( .A(\mem<8><5> ), .B(n3640), .Y(n4550) );
  INVX1 U4378 ( .A(n4550), .Y(n4551) );
  AND2X2 U4379 ( .A(\mem<8><6> ), .B(n3640), .Y(n4552) );
  INVX1 U4380 ( .A(n4552), .Y(n4553) );
  AND2X2 U4381 ( .A(\mem<8><7> ), .B(n3640), .Y(n4554) );
  INVX1 U4382 ( .A(n4554), .Y(n4555) );
  AND2X2 U4383 ( .A(\mem<7><0> ), .B(n3642), .Y(n4556) );
  INVX1 U4384 ( .A(n4556), .Y(n4557) );
  AND2X2 U4385 ( .A(\mem<7><1> ), .B(n3642), .Y(n4558) );
  INVX1 U4386 ( .A(n4558), .Y(n4559) );
  AND2X2 U4387 ( .A(\mem<7><2> ), .B(n3642), .Y(n4560) );
  INVX1 U4388 ( .A(n4560), .Y(n4561) );
  AND2X2 U4389 ( .A(\mem<7><3> ), .B(n3642), .Y(n4562) );
  INVX1 U4390 ( .A(n4562), .Y(n4563) );
  AND2X2 U4391 ( .A(\mem<7><4> ), .B(n3642), .Y(n4564) );
  INVX1 U4392 ( .A(n4564), .Y(n4565) );
  AND2X2 U4393 ( .A(\mem<7><5> ), .B(n3642), .Y(n4566) );
  INVX1 U4394 ( .A(n4566), .Y(n4567) );
  AND2X2 U4395 ( .A(\mem<7><6> ), .B(n3642), .Y(n4568) );
  INVX1 U4396 ( .A(n4568), .Y(n4569) );
  AND2X2 U4397 ( .A(\mem<7><7> ), .B(n3642), .Y(n4570) );
  INVX1 U4398 ( .A(n4570), .Y(n4571) );
  AND2X2 U4399 ( .A(\mem<6><0> ), .B(n4938), .Y(n4572) );
  INVX1 U4400 ( .A(n4572), .Y(n4573) );
  AND2X2 U4401 ( .A(\mem<6><1> ), .B(n4938), .Y(n4574) );
  INVX1 U4402 ( .A(n4574), .Y(n4575) );
  AND2X2 U4403 ( .A(\mem<6><2> ), .B(n4938), .Y(n4576) );
  INVX1 U4404 ( .A(n4576), .Y(n4577) );
  AND2X2 U4405 ( .A(\mem<6><3> ), .B(n4938), .Y(n4578) );
  INVX1 U4406 ( .A(n4578), .Y(n4579) );
  AND2X2 U4407 ( .A(\mem<6><4> ), .B(n4938), .Y(n4580) );
  INVX1 U4408 ( .A(n4580), .Y(n4581) );
  AND2X2 U4409 ( .A(\mem<6><5> ), .B(n4938), .Y(n4582) );
  INVX1 U4410 ( .A(n4582), .Y(n4583) );
  AND2X2 U4411 ( .A(\mem<6><6> ), .B(n4938), .Y(n4584) );
  INVX1 U4412 ( .A(n4584), .Y(n4585) );
  AND2X2 U4413 ( .A(\mem<6><7> ), .B(n4938), .Y(n4586) );
  INVX1 U4414 ( .A(n4586), .Y(n4587) );
  AND2X2 U4415 ( .A(\mem<5><0> ), .B(n4939), .Y(n4588) );
  INVX1 U4416 ( .A(n4588), .Y(n4589) );
  AND2X2 U4417 ( .A(\mem<5><1> ), .B(n4939), .Y(n4590) );
  INVX1 U4418 ( .A(n4590), .Y(n4591) );
  AND2X2 U4419 ( .A(\mem<5><2> ), .B(n4939), .Y(n4592) );
  INVX1 U4420 ( .A(n4592), .Y(n4593) );
  AND2X2 U4421 ( .A(\mem<5><3> ), .B(n4939), .Y(n4594) );
  INVX1 U4422 ( .A(n4594), .Y(n4595) );
  AND2X2 U4423 ( .A(\mem<5><4> ), .B(n4939), .Y(n4596) );
  INVX1 U4424 ( .A(n4596), .Y(n4597) );
  AND2X2 U4425 ( .A(\mem<5><5> ), .B(n4939), .Y(n4598) );
  INVX1 U4426 ( .A(n4598), .Y(n4599) );
  AND2X2 U4427 ( .A(\mem<5><6> ), .B(n4939), .Y(n4600) );
  INVX1 U4428 ( .A(n4600), .Y(n4601) );
  AND2X2 U4429 ( .A(\mem<5><7> ), .B(n4939), .Y(n4602) );
  INVX1 U4430 ( .A(n4602), .Y(n4603) );
  AND2X2 U4431 ( .A(\mem<2><0> ), .B(n3648), .Y(n4604) );
  INVX1 U4432 ( .A(n4604), .Y(n4605) );
  AND2X2 U4433 ( .A(\mem<2><1> ), .B(n3648), .Y(n4606) );
  INVX1 U4434 ( .A(n4606), .Y(n4607) );
  AND2X2 U4435 ( .A(\mem<2><2> ), .B(n3648), .Y(n4608) );
  INVX1 U4436 ( .A(n4608), .Y(n4609) );
  AND2X2 U4437 ( .A(\mem<2><3> ), .B(n3648), .Y(n4610) );
  INVX1 U4438 ( .A(n4610), .Y(n4611) );
  AND2X2 U4439 ( .A(\mem<2><4> ), .B(n3648), .Y(n4612) );
  INVX1 U4440 ( .A(n4612), .Y(n4613) );
  AND2X2 U4441 ( .A(\mem<2><5> ), .B(n3648), .Y(n4614) );
  INVX1 U4442 ( .A(n4614), .Y(n4615) );
  AND2X2 U4443 ( .A(\mem<2><6> ), .B(n3648), .Y(n4616) );
  INVX1 U4444 ( .A(n4616), .Y(n4617) );
  AND2X2 U4445 ( .A(\mem<2><7> ), .B(n3648), .Y(n4618) );
  INVX1 U4446 ( .A(n4618), .Y(n4619) );
  AND2X2 U4447 ( .A(n1051), .B(n5018), .Y(n4620) );
  INVX1 U4448 ( .A(n4620), .Y(n4621) );
  INVX1 U4449 ( .A(n5756), .Y(n4731) );
  INVX1 U4450 ( .A(n3718), .Y(n4622) );
  INVX1 U4451 ( .A(n4809), .Y(n4623) );
  INVX1 U4452 ( .A(n775), .Y(n4624) );
  AND2X2 U4453 ( .A(\mem<46><5> ), .B(n152), .Y(n4625) );
  AND2X2 U4454 ( .A(n4992), .B(n5002), .Y(n4626) );
  INVX1 U4455 ( .A(n4626), .Y(n4627) );
  INVX1 U4456 ( .A(n4626), .Y(n4628) );
  AND2X2 U4457 ( .A(n6415), .B(n4949), .Y(n4629) );
  INVX1 U4458 ( .A(n4629), .Y(n4630) );
  INVX1 U4459 ( .A(n4629), .Y(n4631) );
  AND2X2 U4460 ( .A(n6415), .B(n150), .Y(n4632) );
  INVX1 U4461 ( .A(n4632), .Y(n4633) );
  INVX1 U4462 ( .A(n4632), .Y(n4634) );
  AND2X2 U4463 ( .A(n6415), .B(n4818), .Y(n4635) );
  INVX1 U4464 ( .A(n4635), .Y(n4636) );
  INVX1 U4465 ( .A(n4635), .Y(n4637) );
  AND2X2 U4466 ( .A(n6415), .B(n4957), .Y(n4638) );
  INVX1 U4467 ( .A(n4638), .Y(n4639) );
  INVX1 U4468 ( .A(n4638), .Y(n4640) );
  INVX1 U4469 ( .A(n4638), .Y(n4641) );
  AND2X2 U4470 ( .A(n6415), .B(n4961), .Y(n4642) );
  INVX1 U4471 ( .A(n4642), .Y(n4643) );
  INVX1 U4472 ( .A(n4642), .Y(n4644) );
  INVX1 U4473 ( .A(n4642), .Y(n4645) );
  AND2X2 U4474 ( .A(n6415), .B(n4969), .Y(n4646) );
  INVX1 U4475 ( .A(n4646), .Y(n4647) );
  INVX1 U4476 ( .A(n4646), .Y(n4648) );
  BUFX2 U4477 ( .A(n6334), .Y(n4649) );
  AND2X2 U4478 ( .A(n4966), .B(n4858), .Y(n4650) );
  INVX1 U4479 ( .A(n28), .Y(n4651) );
  INVX1 U4480 ( .A(n3573), .Y(n4652) );
  INVX1 U4481 ( .A(n3713), .Y(n4653) );
  INVX1 U4482 ( .A(n952), .Y(n4654) );
  INVX1 U4483 ( .A(n953), .Y(n4655) );
  INVX1 U4484 ( .A(n954), .Y(n4656) );
  INVX1 U4485 ( .A(n955), .Y(n4657) );
  INVX1 U4486 ( .A(n3717), .Y(n4658) );
  AND2X2 U4487 ( .A(n4961), .B(n3661), .Y(n4659) );
  INVX1 U4488 ( .A(n4659), .Y(n4660) );
  INVX1 U4489 ( .A(n4659), .Y(n4661) );
  INVX1 U4490 ( .A(n3718), .Y(n4662) );
  INVX1 U4491 ( .A(n1031), .Y(n4663) );
  INVX1 U4492 ( .A(n82), .Y(n4969) );
  INVX1 U4493 ( .A(n4666), .Y(n4664) );
  INVX1 U4494 ( .A(n4666), .Y(n4665) );
  AND2X2 U4495 ( .A(n6415), .B(n4858), .Y(n4666) );
  INVX1 U4496 ( .A(n771), .Y(n4667) );
  INVX1 U4497 ( .A(n771), .Y(n4668) );
  INVX1 U4498 ( .A(n4671), .Y(n4669) );
  INVX1 U4499 ( .A(n4671), .Y(n4670) );
  AND2X2 U4500 ( .A(n5018), .B(n5008), .Y(n4671) );
  INVX1 U4501 ( .A(n4880), .Y(n4672) );
  INVX1 U4502 ( .A(n4672), .Y(n4673) );
  INVX1 U4503 ( .A(n4674), .Y(n4675) );
  INVX1 U4504 ( .A(n797), .Y(n4676) );
  INVX1 U4505 ( .A(n4679), .Y(n4677) );
  INVX1 U4506 ( .A(n4679), .Y(n4678) );
  AND2X2 U4507 ( .A(n573), .B(n3847), .Y(n4679) );
  INVX1 U4508 ( .A(n798), .Y(n4680) );
  INVX1 U4509 ( .A(n806), .Y(n4682) );
  INVX1 U4510 ( .A(wr), .Y(n4683) );
  INVX1 U4511 ( .A(enable), .Y(n4684) );
  INVX1 U4512 ( .A(n792), .Y(n4685) );
  INVX1 U4513 ( .A(n792), .Y(n4686) );
  INVX1 U4514 ( .A(n4691), .Y(n4687) );
  INVX1 U4515 ( .A(n4691), .Y(n4688) );
  INVX1 U4516 ( .A(n4691), .Y(n4689) );
  INVX1 U4517 ( .A(n4691), .Y(n4690) );
  AND2X2 U4518 ( .A(n810), .B(n5143), .Y(n4691) );
  INVX1 U4519 ( .A(n831), .Y(n4692) );
  INVX1 U4520 ( .A(n831), .Y(n4693) );
  INVX1 U4521 ( .A(n4698), .Y(n4694) );
  INVX1 U4522 ( .A(n4698), .Y(n4695) );
  INVX1 U4523 ( .A(n4698), .Y(n4696) );
  INVX1 U4524 ( .A(n4698), .Y(n4697) );
  AND2X2 U4525 ( .A(enable), .B(n4683), .Y(n4698) );
  OAI21X1 U4526 ( .A(n5456), .B(n6367), .C(n5455), .Y(n5457) );
  INVX1 U4527 ( .A(\mem<26><3> ), .Y(n5456) );
  AND2X2 U4528 ( .A(n4831), .B(n5203), .Y(n5187) );
  OAI21X1 U4529 ( .A(n4699), .B(n3673), .C(n4700), .Y(n4701) );
  INVX1 U4530 ( .A(\mem<16><4> ), .Y(n4699) );
  INVX1 U4531 ( .A(n5532), .Y(n4700) );
  INVX1 U4532 ( .A(n4701), .Y(n5539) );
  OAI21X1 U4533 ( .A(n4702), .B(n3849), .C(n4703), .Y(n4704) );
  INVX1 U4534 ( .A(\mem<26><0> ), .Y(n4702) );
  INVX1 U4535 ( .A(n5201), .Y(n4703) );
  INVX1 U4536 ( .A(n4704), .Y(n5208) );
  OAI21X1 U4537 ( .A(n4705), .B(n4719), .C(n70), .Y(n4706) );
  INVX1 U4538 ( .A(\mem<56><4> ), .Y(n4705) );
  INVX1 U4539 ( .A(n4706), .Y(n5470) );
  AOI21X1 U4540 ( .A(n4707), .B(n701), .C(n6404), .Y(n4708) );
  INVX1 U4541 ( .A(n5678), .Y(n4707) );
  INVX1 U4542 ( .A(n4708), .Y(n5679) );
  INVX1 U4543 ( .A(n5610), .Y(n4709) );
  INVX1 U4544 ( .A(n5611), .Y(n4710) );
  INVX1 U4545 ( .A(n583), .Y(n4781) );
  AOI22X1 U4546 ( .A(\mem<9><1> ), .B(n4676), .C(n6402), .D(\mem<8><1> ), .Y(
        n5221) );
  INVX2 U4547 ( .A(n3578), .Y(n6402) );
  OAI21X1 U4548 ( .A(n5608), .B(n93), .C(n5607), .Y(n5611) );
  INVX1 U4549 ( .A(\mem<48><5> ), .Y(n5608) );
  INVX1 U4550 ( .A(n6035), .Y(n4711) );
  INVX1 U4551 ( .A(n3564), .Y(n6369) );
  AND2X2 U4552 ( .A(n4712), .B(n4713), .Y(n5625) );
  INVX1 U4553 ( .A(n5623), .Y(n4712) );
  INVX1 U4554 ( .A(n5622), .Y(n4713) );
  NAND3X1 U4555 ( .A(n772), .B(n5539), .C(n5538), .Y(n5540) );
  NAND2X1 U4556 ( .A(\mem<17><0> ), .B(n4856), .Y(n5188) );
  AND2X2 U4557 ( .A(n4714), .B(n4715), .Y(n5207) );
  INVX1 U4558 ( .A(n5205), .Y(n4714) );
  INVX1 U4559 ( .A(n5206), .Y(n4715) );
  NAND3X1 U4560 ( .A(n5010), .B(n5020), .C(n4885), .Y(n4716) );
  INVX1 U4561 ( .A(n4716), .Y(n5133) );
  INVX4 U4562 ( .A(n5011), .Y(n5020) );
  OAI21X1 U4563 ( .A(n5621), .B(n3849), .C(n1186), .Y(n5622) );
  INVX1 U4564 ( .A(\mem<26><5> ), .Y(n5621) );
  AND2X2 U4565 ( .A(n4727), .B(n4717), .Y(n5515) );
  INVX1 U4566 ( .A(n5514), .Y(n4717) );
  OAI21X1 U4567 ( .A(n5506), .B(n4917), .C(n5505), .Y(n5514) );
  INVX1 U4568 ( .A(\mem<41><4> ), .Y(n5506) );
  OAI21X1 U4569 ( .A(n4718), .B(n4719), .C(n69), .Y(n4720) );
  INVX1 U4570 ( .A(\mem<56><6> ), .Y(n4718) );
  INVX1 U4571 ( .A(n4720), .Y(n5635) );
  AOI21X1 U4572 ( .A(\mem<33><6> ), .B(n3880), .C(n5628), .Y(n5636) );
  AND2X2 U4573 ( .A(n4721), .B(n4722), .Y(n5770) );
  INVX1 U4574 ( .A(n5764), .Y(n4721) );
  INVX1 U4575 ( .A(n5765), .Y(n4722) );
  AOI21X1 U4576 ( .A(n793), .B(n794), .C(n4696), .Y(\data_out<1> ) );
  NAND3X1 U4577 ( .A(n3991), .B(n2392), .C(n3118), .Y(n6917) );
  NAND3X1 U4578 ( .A(n3989), .B(n2390), .C(n3116), .Y(n6918) );
  NAND3X1 U4579 ( .A(n3987), .B(n2388), .C(n3114), .Y(n6919) );
  NAND3X1 U4580 ( .A(n3985), .B(n2386), .C(n3112), .Y(n6920) );
  NAND3X1 U4581 ( .A(n3983), .B(n2384), .C(n3110), .Y(n6921) );
  NAND3X1 U4582 ( .A(n3981), .B(n2382), .C(n3108), .Y(n6922) );
  NAND3X1 U4583 ( .A(n3979), .B(n2380), .C(n3106), .Y(n6923) );
  NAND3X1 U4584 ( .A(n3977), .B(n2378), .C(n3104), .Y(n6924) );
  NAND3X1 U4585 ( .A(n4977), .B(n3566), .C(n4667), .Y(n6291) );
  OAI21X1 U4586 ( .A(n5762), .B(n815), .C(n5761), .Y(n5765) );
  INVX1 U4587 ( .A(\mem<48><7> ), .Y(n5762) );
  AND2X2 U4588 ( .A(\mem<12><4> ), .B(n3654), .Y(n4723) );
  INVX1 U4589 ( .A(n4723), .Y(n5522) );
  INVX1 U4590 ( .A(n122), .Y(n4724) );
  INVX1 U4591 ( .A(n4858), .Y(n4725) );
  NAND3X1 U4592 ( .A(n847), .B(n3975), .C(n3796), .Y(n6925) );
  NAND3X1 U4593 ( .A(n845), .B(n3973), .C(n3794), .Y(n6926) );
  NAND3X1 U4594 ( .A(n843), .B(n3971), .C(n3792), .Y(n6927) );
  NAND3X1 U4595 ( .A(n841), .B(n3969), .C(n3790), .Y(n6928) );
  NAND3X1 U4596 ( .A(n839), .B(n3967), .C(n3788), .Y(n6929) );
  NAND3X1 U4597 ( .A(n837), .B(n3965), .C(n3786), .Y(n6930) );
  NAND3X1 U4598 ( .A(n835), .B(n3963), .C(n3784), .Y(n6931) );
  NAND3X1 U4599 ( .A(n833), .B(n3961), .C(n3782), .Y(n6932) );
  OAI21X1 U4600 ( .A(n5523), .B(n93), .C(n5522), .Y(n5526) );
  INVX1 U4601 ( .A(\mem<48><4> ), .Y(n5523) );
  OAI21X1 U4602 ( .A(n3565), .B(n4667), .C(n4977), .Y(n6293) );
  AND2X2 U4603 ( .A(n4832), .B(n4873), .Y(n4877) );
  INVX1 U4604 ( .A(n4668), .Y(n6289) );
  AND2X2 U4605 ( .A(n3574), .B(n6313), .Y(n4726) );
  INVX1 U4606 ( .A(n4726), .Y(n6311) );
  AOI21X1 U4607 ( .A(\mem<57><4> ), .B(n6303), .C(n1261), .Y(n4727) );
  INVX1 U4608 ( .A(n5603), .Y(n4728) );
  INVX1 U4609 ( .A(n5604), .Y(n4729) );
  INVX1 U4610 ( .A(n6223), .Y(n4730) );
  NAND3X1 U4611 ( .A(n67), .B(n4731), .C(n4732), .Y(n4733) );
  INVX1 U4612 ( .A(n5757), .Y(n4732) );
  INVX1 U4613 ( .A(n4733), .Y(n5758) );
  INVX1 U4614 ( .A(\mem<49><6> ), .Y(n4734) );
  INVX1 U4615 ( .A(n4884), .Y(n4735) );
  INVX1 U4616 ( .A(n777), .Y(n6298) );
  AND2X2 U4617 ( .A(n4736), .B(n4737), .Y(n5600) );
  INVX1 U4618 ( .A(n5598), .Y(n4736) );
  INVX1 U4619 ( .A(n5599), .Y(n4737) );
  INVX1 U4620 ( .A(n5681), .Y(n4738) );
  INVX1 U4621 ( .A(n5682), .Y(n4739) );
  OAI21X1 U4622 ( .A(n5671), .B(n3677), .C(n5670), .Y(n5682) );
  INVX1 U4623 ( .A(\mem<41><6> ), .Y(n5671) );
  INVX1 U4624 ( .A(n6286), .Y(n4740) );
  INVX1 U4625 ( .A(n5909), .Y(n4741) );
  INVX1 U4626 ( .A(n6353), .Y(n6350) );
  NOR3X1 U4627 ( .A(n5126), .B(n4913), .C(n4725), .Y(n4742) );
  INVX1 U4628 ( .A(n4742), .Y(n6361) );
  AOI21X1 U4629 ( .A(n4665), .B(n4857), .C(n4978), .Y(n4743) );
  INVX1 U4630 ( .A(n4743), .Y(n6365) );
  INVX1 U4631 ( .A(n6160), .Y(n4744) );
  AND2X2 U4632 ( .A(n4745), .B(n674), .Y(n5541) );
  INVX1 U4633 ( .A(n5540), .Y(n4745) );
  INVX1 U4634 ( .A(n5776), .Y(n4746) );
  INVX1 U4635 ( .A(n5775), .Y(n4747) );
  INVX1 U4636 ( .A(n5972), .Y(n4748) );
  AND2X2 U4637 ( .A(n3576), .B(\mem<25><5> ), .Y(n4749) );
  INVX1 U4638 ( .A(n4749), .Y(n5589) );
  OAI21X1 U4639 ( .A(n5590), .B(n4917), .C(n5589), .Y(n5599) );
  INVX1 U4640 ( .A(\mem<41><5> ), .Y(n5590) );
  NAND2X1 U4641 ( .A(\mem<17><1> ), .B(n4856), .Y(n5212) );
  INVX1 U4642 ( .A(\mem<24><4> ), .Y(n4750) );
  INVX1 U4643 ( .A(n3868), .Y(n4751) );
  OAI21X1 U4644 ( .A(n5680), .B(n104), .C(n5679), .Y(n5681) );
  INVX1 U4645 ( .A(\mem<57><6> ), .Y(n5680) );
  AOI21X1 U4646 ( .A(n4752), .B(n689), .C(n6404), .Y(n4753) );
  INVX1 U4647 ( .A(n5595), .Y(n4752) );
  INVX1 U4648 ( .A(n4753), .Y(n5596) );
  OAI21X1 U4649 ( .A(n5597), .B(n104), .C(n5596), .Y(n5598) );
  INVX1 U4650 ( .A(\mem<57><5> ), .Y(n5597) );
  INVX1 U4651 ( .A(n4861), .Y(n4754) );
  AOI21X1 U4652 ( .A(n3847), .B(\mem<15><2> ), .C(n5314), .Y(n5323) );
  INVX1 U4653 ( .A(\addr<14> ), .Y(n5112) );
  INVX1 U4654 ( .A(n5537), .Y(n4755) );
  INVX1 U4655 ( .A(n5536), .Y(n4756) );
  OAI21X1 U4656 ( .A(n4757), .B(n6345), .C(n4758), .Y(n4759) );
  INVX1 U4657 ( .A(\mem<33><5> ), .Y(n4757) );
  INVX1 U4658 ( .A(n5544), .Y(n4758) );
  INVX1 U4659 ( .A(n4759), .Y(n5554) );
  OAI21X1 U4660 ( .A(n5535), .B(n3849), .C(n1174), .Y(n5536) );
  INVX1 U4661 ( .A(\mem<26><4> ), .Y(n5535) );
  AND2X2 U4662 ( .A(n115), .B(n5187), .Y(n4856) );
  INVX4 U4663 ( .A(n3675), .Y(n6415) );
  NAND3X1 U4664 ( .A(n1285), .B(n802), .C(n704), .Y(n4760) );
  INVX1 U4665 ( .A(n4760), .Y(n5710) );
  INVX2 U4666 ( .A(n6362), .Y(n6360) );
  NAND3X1 U4667 ( .A(n4021), .B(n2744), .C(n3356), .Y(n6653) );
  NAND3X1 U4668 ( .A(n4019), .B(n2742), .C(n3354), .Y(n6654) );
  NAND3X1 U4669 ( .A(n4017), .B(n2740), .C(n3352), .Y(n6655) );
  NAND3X1 U4670 ( .A(n4015), .B(n2738), .C(n3350), .Y(n6656) );
  NAND3X1 U4671 ( .A(n4013), .B(n2736), .C(n3348), .Y(n6657) );
  NAND3X1 U4672 ( .A(n4011), .B(n2734), .C(n3346), .Y(n6658) );
  NAND3X1 U4673 ( .A(n4009), .B(n2732), .C(n3344), .Y(n6659) );
  NAND3X1 U4674 ( .A(n4007), .B(n2730), .C(n3342), .Y(n6660) );
  INVX1 U4675 ( .A(n5518), .Y(n4761) );
  INVX1 U4676 ( .A(n5519), .Y(n4762) );
  AND2X2 U4677 ( .A(n17), .B(\mem<49><4> ), .Y(n4763) );
  INVX1 U4678 ( .A(n4763), .Y(n5460) );
  AND2X2 U4679 ( .A(n4826), .B(n3673), .Y(n4764) );
  AND2X2 U4680 ( .A(n4898), .B(n4765), .Y(n4858) );
  INVX1 U4681 ( .A(n5115), .Y(n4765) );
  NAND2X1 U4682 ( .A(\mem<52><3> ), .B(n4877), .Y(n5381) );
  NOR3X1 U4683 ( .A(N181), .B(n5009), .C(n4885), .Y(n4766) );
  INVX1 U4684 ( .A(n4766), .Y(n5114) );
  NOR3X1 U4685 ( .A(N178), .B(n4811), .C(n4817), .Y(n4767) );
  INVX4 U4686 ( .A(n4767), .Y(n6404) );
  INVX1 U4687 ( .A(n5002), .Y(n4811) );
  AND2X2 U4688 ( .A(n4768), .B(n4769), .Y(n5211) );
  INVX1 U4689 ( .A(n5210), .Y(n4768) );
  INVX1 U4690 ( .A(n604), .Y(n4769) );
  OAI21X1 U4691 ( .A(n5774), .B(n3849), .C(n5773), .Y(n5775) );
  INVX1 U4692 ( .A(\mem<26><7> ), .Y(n5774) );
  OAI21X1 U4693 ( .A(n3871), .B(n5200), .C(n5199), .Y(n5201) );
  INVX1 U4694 ( .A(\mem<49><0> ), .Y(n5200) );
  AOI21X1 U4695 ( .A(n3847), .B(\mem<15><3> ), .C(n5402), .Y(n5410) );
  OAI21X1 U4696 ( .A(n3669), .B(n5382), .C(n5381), .Y(n5386) );
  INVX1 U4697 ( .A(\mem<50><3> ), .Y(n5382) );
  AND2X2 U4698 ( .A(n4911), .B(\mem<18><7> ), .Y(n4770) );
  INVX1 U4699 ( .A(n4770), .Y(n5771) );
  OAI21X1 U4700 ( .A(n5772), .B(n6344), .C(n5771), .Y(n5776) );
  INVX1 U4701 ( .A(\mem<34><7> ), .Y(n5772) );
  INVX1 U4702 ( .A(n5686), .Y(n4771) );
  INVX1 U4703 ( .A(n5687), .Y(n4772) );
  AND2X2 U4704 ( .A(n561), .B(n813), .Y(n6410) );
  NOR3X1 U4705 ( .A(n6350), .B(n3870), .C(n6358), .Y(n4773) );
  INVX1 U4706 ( .A(n4773), .Y(n6355) );
  NOR3X1 U4707 ( .A(n3854), .B(n117), .C(n4774), .Y(n4775) );
  INVX1 U4708 ( .A(n5133), .Y(n4774) );
  INVX1 U4709 ( .A(n4775), .Y(n6403) );
  NAND3X1 U4710 ( .A(n277), .B(n979), .C(n4380), .Y(n6669) );
  NAND3X1 U4711 ( .A(n275), .B(n977), .C(n4379), .Y(n6670) );
  NAND3X1 U4712 ( .A(n273), .B(n975), .C(n4377), .Y(n6671) );
  NAND3X1 U4713 ( .A(n271), .B(n973), .C(n4375), .Y(n6672) );
  NAND3X1 U4714 ( .A(n269), .B(n971), .C(n4372), .Y(n6673) );
  NAND3X1 U4715 ( .A(n267), .B(n969), .C(n4371), .Y(n6674) );
  NAND3X1 U4716 ( .A(n265), .B(n967), .C(n4369), .Y(n6675) );
  NAND3X1 U4717 ( .A(n263), .B(n965), .C(n4367), .Y(n6676) );
  INVX1 U4718 ( .A(n5438), .Y(n4776) );
  INVX1 U4719 ( .A(n5439), .Y(n4777) );
  INVX1 U4720 ( .A(n5433), .Y(n4778) );
  INVX1 U4721 ( .A(n5434), .Y(n4779) );
  NAND3X1 U4722 ( .A(n1283), .B(n5635), .C(n5636), .Y(n5687) );
  NAND3X1 U4723 ( .A(n1281), .B(n5553), .C(n5554), .Y(n5604) );
  INVX1 U4724 ( .A(n608), .Y(n4780) );
  NOR2X1 U4725 ( .A(n4782), .B(n3879), .Y(n4783) );
  INVX1 U4726 ( .A(\mem<33><1> ), .Y(n4782) );
  INVX1 U4727 ( .A(n4783), .Y(n5222) );
  AOI21X1 U4728 ( .A(n4784), .B(n658), .C(n6404), .Y(n4785) );
  INVX1 U4729 ( .A(n5430), .Y(n4784) );
  INVX1 U4730 ( .A(n4785), .Y(n5431) );
  INVX1 U4731 ( .A(n5353), .Y(n4786) );
  AND2X2 U4732 ( .A(n4787), .B(n4788), .Y(n5219) );
  INVX1 U4733 ( .A(n5217), .Y(n4787) );
  INVX1 U4734 ( .A(n5218), .Y(n4788) );
  INVX1 U4735 ( .A(n5290), .Y(n4789) );
  NAND3X1 U4736 ( .A(n4790), .B(n4791), .C(n4792), .Y(n4793) );
  INVX1 U4737 ( .A(n5366), .Y(n4790) );
  INVX1 U4738 ( .A(n5367), .Y(n4791) );
  INVX1 U4739 ( .A(n4872), .Y(n4792) );
  INVX1 U4740 ( .A(n4793), .Y(n5374) );
  INVX1 U4741 ( .A(n5227), .Y(n4794) );
  INVX1 U4742 ( .A(n5228), .Y(n4795) );
  NAND3X1 U4743 ( .A(n5350), .B(n4061), .C(n1264), .Y(n5353) );
  NAND3X1 U4744 ( .A(N180), .B(n5013), .C(n4885), .Y(n4796) );
  INVX1 U4745 ( .A(n4796), .Y(n5127) );
  NAND3X1 U4746 ( .A(n5471), .B(n5470), .C(n1279), .Y(n5519) );
  OAI21X1 U4747 ( .A(n5461), .B(n4678), .C(n5460), .Y(n5462) );
  INVX1 U4748 ( .A(\mem<9><4> ), .Y(n5461) );
  AND2X2 U4749 ( .A(n4797), .B(n4798), .Y(n5360) );
  INVX1 U4750 ( .A(n5358), .Y(n4797) );
  INVX1 U4751 ( .A(n5359), .Y(n4798) );
  NAND3X1 U4752 ( .A(n5287), .B(n2350), .C(n3096), .Y(n5290) );
  NAND3X1 U4753 ( .A(n4799), .B(n4800), .C(n4121), .Y(n5439) );
  INVX1 U4754 ( .A(n5379), .Y(n4799) );
  INVX1 U4755 ( .A(n5380), .Y(n4800) );
  INVX1 U4756 ( .A(n4863), .Y(n4801) );
  AOI21X1 U4757 ( .A(n4802), .B(n671), .C(n6404), .Y(n4803) );
  INVX1 U4758 ( .A(n5513), .Y(n4802) );
  NAND3X1 U4759 ( .A(n4804), .B(n4805), .C(n709), .Y(n4806) );
  INVX1 U4760 ( .A(n5759), .Y(n4804) );
  INVX1 U4761 ( .A(n5760), .Y(n4805) );
  INVX1 U4762 ( .A(n4806), .Y(n5782) );
  NAND3X1 U4763 ( .A(n4807), .B(n4808), .C(n4871), .Y(n4872) );
  INVX1 U4764 ( .A(n5371), .Y(n4807) );
  INVX1 U4765 ( .A(n5372), .Y(n4808) );
  AND2X2 U4766 ( .A(n4866), .B(n5192), .Y(n4809) );
  INVX1 U4767 ( .A(n3572), .Y(n4810) );
  INVX1 U4768 ( .A(n4910), .Y(n4812) );
  INVX1 U4769 ( .A(n6314), .Y(n4813) );
  INVX1 U4770 ( .A(n4825), .Y(n4814) );
  INVX1 U4771 ( .A(n3879), .Y(n4844) );
  OR2X2 U4772 ( .A(n82), .B(n5198), .Y(n4815) );
  INVX1 U4773 ( .A(n4953), .Y(n4818) );
  AND2X2 U4774 ( .A(n3861), .B(n5034), .Y(n4820) );
  INVX1 U4775 ( .A(n6401), .Y(n4821) );
  INVX1 U4776 ( .A(n4843), .Y(n4822) );
  INVX2 U4777 ( .A(n4955), .Y(n4954) );
  BUFX2 U4778 ( .A(n4835), .Y(n4824) );
  INVX1 U4779 ( .A(n4855), .Y(n4825) );
  INVX1 U4780 ( .A(n4856), .Y(n6388) );
  INVX1 U4781 ( .A(n6400), .Y(n4827) );
  INVX1 U4782 ( .A(n4827), .Y(n4828) );
  INVX1 U4783 ( .A(n3654), .Y(n4830) );
  NOR3X1 U4784 ( .A(n805), .B(n4621), .C(n3854), .Y(n4831) );
  INVX1 U4785 ( .A(n750), .Y(n4832) );
  OR2X2 U4786 ( .A(n4833), .B(n4843), .Y(n5199) );
  INVX1 U4787 ( .A(n3567), .Y(n6333) );
  INVX1 U4788 ( .A(n6410), .Y(n4968) );
  BUFX4 U4789 ( .A(n6404), .Y(n4834) );
  INVX1 U4790 ( .A(n4812), .Y(n4835) );
  OR2X2 U4791 ( .A(n4837), .B(n4829), .Y(n5761) );
  INVX4 U4792 ( .A(n6403), .Y(n4838) );
  INVX1 U4793 ( .A(n561), .Y(n4840) );
  NOR3X1 U4794 ( .A(n5017), .B(n5033), .C(n5010), .Y(n4842) );
  INVX1 U4795 ( .A(n4855), .Y(n4843) );
  AND2X2 U4796 ( .A(n122), .B(n4954), .Y(n4845) );
  INVX8 U4797 ( .A(n4845), .Y(n6344) );
  AND2X2 U4798 ( .A(n4954), .B(n4832), .Y(n4846) );
  INVX1 U4799 ( .A(n6312), .Y(n4847) );
  INVX1 U4800 ( .A(n4847), .Y(n4848) );
  INVX1 U4801 ( .A(n3576), .Y(n4849) );
  INVX1 U4802 ( .A(n4910), .Y(n4850) );
  INVX1 U4803 ( .A(n578), .Y(n4851) );
  INVX1 U4804 ( .A(n6414), .Y(n6413) );
  INVX1 U4805 ( .A(n81), .Y(n4971) );
  INVX1 U4806 ( .A(n4972), .Y(n4970) );
  AND2X2 U4807 ( .A(n3712), .B(n4853), .Y(n4884) );
  AND2X2 U4808 ( .A(n4981), .B(n582), .Y(n4910) );
  AND2X2 U4809 ( .A(n4981), .B(n818), .Y(n4855) );
  INVX1 U4810 ( .A(n4855), .Y(n6345) );
  INVX1 U4811 ( .A(n4865), .Y(n4981) );
  INVX1 U4812 ( .A(n6363), .Y(n4857) );
  INVX1 U4813 ( .A(n6344), .Y(n6343) );
  INVX1 U4814 ( .A(n5751), .Y(n4859) );
  INVX1 U4815 ( .A(n13), .Y(n6387) );
  INVX1 U4816 ( .A(n3874), .Y(n4913) );
  AND2X2 U4817 ( .A(n4913), .B(\mem<17><2> ), .Y(n4860) );
  INVX4 U4818 ( .A(n5013), .Y(n5011) );
  INVX1 U4819 ( .A(n4956), .Y(n4955) );
  AND2X2 U4820 ( .A(n4867), .B(n5203), .Y(n4861) );
  INVX1 U4821 ( .A(n6303), .Y(n4862) );
  AND2X2 U4822 ( .A(n573), .B(\mem<57><2> ), .Y(n4863) );
  AND2X2 U4823 ( .A(n4832), .B(n80), .Y(n4864) );
  INVX8 U4824 ( .A(n4864), .Y(n6414) );
  INVX1 U4825 ( .A(n561), .Y(n4865) );
  INVX2 U4826 ( .A(N181), .Y(n5013) );
  INVX8 U4827 ( .A(n5036), .Y(n5029) );
  INVX1 U4828 ( .A(n5011), .Y(n5019) );
  INVX1 U4829 ( .A(N180), .Y(n5010) );
  INVX1 U4830 ( .A(n568), .Y(n4866) );
  INVX1 U4831 ( .A(n561), .Y(n4980) );
  INVX1 U4832 ( .A(n3578), .Y(n4869) );
  INVX1 U4833 ( .A(n4869), .Y(n4870) );
  INVX1 U4834 ( .A(n5373), .Y(n4871) );
  INVX1 U4835 ( .A(\data_in<4> ), .Y(n5058) );
  INVX1 U4836 ( .A(\data_in<4> ), .Y(n5059) );
  INVX1 U4837 ( .A(\data_in<5> ), .Y(n5062) );
  INVX1 U4838 ( .A(\data_in<5> ), .Y(n5063) );
  INVX1 U4839 ( .A(n93), .Y(n6315) );
  INVX1 U4840 ( .A(n4877), .Y(n4874) );
  INVX1 U4841 ( .A(n4874), .Y(n4875) );
  INVX1 U4842 ( .A(n4874), .Y(n4876) );
  INVX1 U4843 ( .A(n819), .Y(n4878) );
  INVX2 U4844 ( .A(\data_in<3> ), .Y(n5054) );
  NAND3X1 U4845 ( .A(n5134), .B(n3861), .C(n4842), .Y(n4880) );
  INVX1 U4846 ( .A(n5023), .Y(n4883) );
  INVX1 U4847 ( .A(N182), .Y(n5023) );
  INVX1 U4848 ( .A(n804), .Y(n6347) );
  INVX1 U4849 ( .A(n4884), .Y(n6288) );
  NOR2X1 U4850 ( .A(n4886), .B(n566), .Y(n5717) );
  MUX2X1 U4851 ( .B(n6282), .A(n6283), .S(n4841), .Y(n6284) );
  INVX1 U4852 ( .A(n4820), .Y(n4888) );
  INVX1 U4853 ( .A(n4820), .Y(n4889) );
  INVX1 U4854 ( .A(n4895), .Y(n4890) );
  INVX1 U4855 ( .A(n4888), .Y(n4891) );
  INVX1 U4856 ( .A(n4900), .Y(n4892) );
  INVX1 U4857 ( .A(n4940), .Y(n4894) );
  INVX1 U4858 ( .A(n4941), .Y(n4895) );
  INVX1 U4859 ( .A(n4894), .Y(n4896) );
  INVX1 U4860 ( .A(n4894), .Y(n4897) );
  INVX1 U4861 ( .A(n4888), .Y(n4898) );
  INVX1 U4862 ( .A(n4895), .Y(n4899) );
  INVX1 U4863 ( .A(n4940), .Y(n4900) );
  INVX1 U4864 ( .A(n121), .Y(n4901) );
  INVX1 U4865 ( .A(n4941), .Y(n4902) );
  INVX1 U4866 ( .A(n4901), .Y(n4903) );
  INVX1 U4867 ( .A(n4900), .Y(n4904) );
  INVX1 U4868 ( .A(n4901), .Y(n4905) );
  INVX1 U4869 ( .A(n4902), .Y(n4906) );
  INVX1 U4870 ( .A(n127), .Y(n4907) );
  INVX1 U4871 ( .A(n127), .Y(n4908) );
  INVX1 U4872 ( .A(n4942), .Y(n4940) );
  INVX1 U4873 ( .A(\data_in<6> ), .Y(n5067) );
  INVX1 U4874 ( .A(\data_in<6> ), .Y(n5068) );
  INVX1 U4875 ( .A(n4873), .Y(n4909) );
  INVX1 U4876 ( .A(n6312), .Y(n4950) );
  INVX1 U4877 ( .A(n5126), .Y(n5167) );
  NOR3X1 U4878 ( .A(n4817), .B(n4628), .C(n15), .Y(n4912) );
  INVX1 U4879 ( .A(n4820), .Y(n4942) );
  INVX1 U4880 ( .A(\addr<11> ), .Y(n4914) );
  INVX1 U4881 ( .A(n4942), .Y(n4941) );
  INVX1 U4882 ( .A(n5019), .Y(n5018) );
  INVX1 U4883 ( .A(\data_in<2> ), .Y(n5050) );
  INVX1 U4884 ( .A(n4847), .Y(n4948) );
  INVX1 U4885 ( .A(n3652), .Y(n6303) );
  INVX1 U4886 ( .A(n4839), .Y(n5113) );
  INVX4 U4887 ( .A(n6361), .Y(n6363) );
  BUFX4 U4888 ( .A(n6299), .Y(n4922) );
  BUFX4 U4889 ( .A(n6376), .Y(n4935) );
  BUFX4 U4890 ( .A(n6396), .Y(n4937) );
  INVX8 U4891 ( .A(n5115), .Y(n4947) );
  INVX8 U4892 ( .A(n4979), .Y(n4973) );
  INVX8 U4893 ( .A(n4979), .Y(n4974) );
  INVX8 U4894 ( .A(n4979), .Y(n4975) );
  INVX8 U4895 ( .A(n4978), .Y(n4976) );
  INVX8 U4896 ( .A(n4978), .Y(n4977) );
  INVX8 U4897 ( .A(n6417), .Y(n4978) );
  INVX8 U4898 ( .A(n6417), .Y(n4979) );
  INVX8 U4899 ( .A(n4993), .Y(n4984) );
  INVX8 U4900 ( .A(n4993), .Y(n4985) );
  INVX8 U4901 ( .A(n4994), .Y(n4986) );
  INVX8 U4902 ( .A(n4994), .Y(n4987) );
  INVX8 U4903 ( .A(n4995), .Y(n4988) );
  INVX8 U4904 ( .A(n4995), .Y(n4989) );
  INVX8 U4905 ( .A(n4995), .Y(n4990) );
  INVX8 U4906 ( .A(n4996), .Y(n4991) );
  INVX8 U4907 ( .A(n4994), .Y(n4992) );
  INVX8 U4908 ( .A(N178), .Y(n4994) );
  INVX8 U4909 ( .A(N178), .Y(n4995) );
  INVX8 U4910 ( .A(n5005), .Y(n4997) );
  INVX8 U4911 ( .A(n5005), .Y(n4998) );
  INVX8 U4912 ( .A(n5005), .Y(n4999) );
  INVX8 U4913 ( .A(n5004), .Y(n5000) );
  INVX8 U4914 ( .A(n5004), .Y(n5001) );
  INVX8 U4915 ( .A(n5003), .Y(n5002) );
  INVX4 U4916 ( .A(N179), .Y(n5003) );
  INVX4 U4917 ( .A(N179), .Y(n5004) );
  INVX4 U4918 ( .A(N179), .Y(n5005) );
  INVX8 U4919 ( .A(n5009), .Y(n5006) );
  INVX8 U4920 ( .A(n5010), .Y(n5007) );
  INVX8 U4921 ( .A(n5009), .Y(n5008) );
  INVX8 U4922 ( .A(n5021), .Y(n5014) );
  INVX8 U4923 ( .A(n5021), .Y(n5015) );
  INVX8 U4924 ( .A(n5021), .Y(n5016) );
  INVX8 U4925 ( .A(n5020), .Y(n5017) );
  INVX8 U4926 ( .A(n5034), .Y(n5024) );
  INVX8 U4927 ( .A(n5034), .Y(n5025) );
  INVX8 U4928 ( .A(n5034), .Y(n5026) );
  INVX8 U4929 ( .A(n5035), .Y(n5027) );
  INVX8 U4930 ( .A(n5035), .Y(n5028) );
  INVX8 U4931 ( .A(n4885), .Y(n5033) );
  INVX8 U4932 ( .A(n5040), .Y(n5038) );
  INVX8 U4933 ( .A(n5040), .Y(n5039) );
  INVX8 U4934 ( .A(n5046), .Y(n5041) );
  INVX8 U4935 ( .A(n5046), .Y(n5042) );
  INVX8 U4936 ( .A(n5046), .Y(n5043) );
  INVX8 U4937 ( .A(n5046), .Y(n5044) );
  INVX8 U4938 ( .A(n5046), .Y(n5045) );
  INVX8 U4939 ( .A(\data_in<1> ), .Y(n5046) );
  INVX8 U4940 ( .A(n5054), .Y(n5052) );
  INVX8 U4941 ( .A(n5071), .Y(n5069) );
  INVX8 U4942 ( .A(n5071), .Y(n5070) );
  INVX8 U4943 ( .A(n5076), .Y(n5072) );
  INVX8 U4944 ( .A(n5076), .Y(n5073) );
  INVX8 U4945 ( .A(n5076), .Y(n5074) );
  INVX8 U4946 ( .A(n5080), .Y(n5077) );
  INVX8 U4947 ( .A(n5081), .Y(n5078) );
  INVX8 U4948 ( .A(n5086), .Y(n5082) );
  INVX8 U4949 ( .A(n5086), .Y(n5084) );
  INVX8 U4950 ( .A(n5091), .Y(n5089) );
  INVX8 U4951 ( .A(n5097), .Y(n5094) );
  INVX8 U4952 ( .A(n5097), .Y(n5095) );
  INVX8 U4953 ( .A(n5101), .Y(n5098) );
  INVX8 U4954 ( .A(n5101), .Y(n5099) );
  INVX8 U4955 ( .A(n5105), .Y(n5102) );
  INVX8 U4956 ( .A(n5106), .Y(n5103) );
  INVX8 U4957 ( .A(n5110), .Y(n5107) );
  INVX8 U4958 ( .A(n5111), .Y(n5108) );
  INVX4 U4959 ( .A(\data_in<15> ), .Y(n5110) );
  INVX4 U4960 ( .A(\data_in<15> ), .Y(n5111) );
  NOR3X1 U4961 ( .A(\addr<15> ), .B(n5114), .C(n5113), .Y(n5751) );
  OR2X2 U4962 ( .A(n5002), .B(n4992), .Y(n5198) );
  INVX2 U4963 ( .A(n5198), .Y(n5203) );
  OR2X2 U4964 ( .A(n5002), .B(n4995), .Y(n5126) );
  OR2X2 U4965 ( .A(n4669), .B(\addr<15> ), .Y(n5115) );
  NAND2X1 U4966 ( .A(\mem<20><0> ), .B(n6377), .Y(n5116) );
  OAI21X1 U4967 ( .A(n4), .B(n5117), .C(n5116), .Y(n5118) );
  AOI21X1 U4968 ( .A(\mem<42><0> ), .B(n6331), .C(n5118), .Y(n5125) );
  AOI22X1 U4969 ( .A(\mem<58><0> ), .B(n83), .C(\mem<28><0> ), .D(n6363), .Y(
        n5124) );
  OAI21X1 U4970 ( .A(n6344), .B(n5119), .C(n1134), .Y(n5123) );
  NAND2X1 U4971 ( .A(\mem<18><0> ), .B(n4911), .Y(n5120) );
  OAI21X1 U4972 ( .A(n6342), .B(n5121), .C(n5120), .Y(n5122) );
  NAND3X1 U4973 ( .A(n5134), .B(n3861), .C(n5127), .Y(n6390) );
  NOR2X1 U4974 ( .A(n137), .B(n5128), .Y(n5129) );
  AOI21X1 U4975 ( .A(\mem<11><0> ), .B(n4961), .C(n5129), .Y(n5139) );
  OR2X2 U4976 ( .A(n4669), .B(\addr<15> ), .Y(n5130) );
  AND2X2 U4977 ( .A(\mem<27><0> ), .B(n4853), .Y(n5131) );
  OAI21X1 U4978 ( .A(n2328), .B(n113), .C(n3891), .Y(n5132) );
  AOI21X1 U4979 ( .A(\mem<19><0> ), .B(n4957), .C(n5132), .Y(n5138) );
  OAI21X1 U4980 ( .A(n4953), .B(n5135), .C(n3893), .Y(n5136) );
  AOI21X1 U4981 ( .A(\mem<3><0> ), .B(n4838), .C(n5136), .Y(n5137) );
  AND2X2 U4982 ( .A(\addr<13> ), .B(\addr<12> ), .Y(n5140) );
  NAND3X1 U4983 ( .A(n3854), .B(\addr<14> ), .C(n5140), .Y(n5141) );
  NOR3X1 U4984 ( .A(n4993), .B(n4670), .C(n5003), .Y(n5142) );
  NOR2X1 U4985 ( .A(n4689), .B(n6420), .Y(n5144) );
  OAI21X1 U4986 ( .A(n3658), .B(n5145), .C(n3895), .Y(n5146) );
  NOR2X1 U4987 ( .A(n131), .B(n5147), .Y(n5148) );
  AOI21X1 U4988 ( .A(\mem<15><0> ), .B(n4961), .C(n5148), .Y(n5156) );
  NAND2X1 U4989 ( .A(\mem<63><0> ), .B(n4946), .Y(n5150) );
  AND2X2 U4990 ( .A(\mem<31><0> ), .B(n4765), .Y(n5149) );
  OAI21X1 U4991 ( .A(n5150), .B(n4945), .C(n3897), .Y(n5151) );
  AOI21X1 U4992 ( .A(\mem<23><0> ), .B(n4959), .C(n5151), .Y(n5155) );
  OAI21X1 U4993 ( .A(n4953), .B(n5152), .C(n3899), .Y(n5153) );
  AOI21X1 U4994 ( .A(\mem<7><0> ), .B(n4838), .C(n5153), .Y(n5154) );
  NOR2X1 U4995 ( .A(n141), .B(n5157), .Y(n5158) );
  AOI21X1 U4996 ( .A(\mem<13><0> ), .B(n4961), .C(n5158), .Y(n5166) );
  NAND2X1 U4997 ( .A(\mem<61><0> ), .B(n4946), .Y(n5160) );
  AND2X2 U4998 ( .A(\mem<29><0> ), .B(n4853), .Y(n5159) );
  OAI21X1 U4999 ( .A(n5160), .B(n4945), .C(n3901), .Y(n5161) );
  AOI21X1 U5000 ( .A(\mem<21><0> ), .B(n4957), .C(n5161), .Y(n5165) );
  OAI21X1 U5001 ( .A(n4953), .B(n5162), .C(n1136), .Y(n5163) );
  AOI21X1 U5002 ( .A(\mem<5><0> ), .B(n4838), .C(n5163), .Y(n5164) );
  AOI22X1 U5003 ( .A(n4964), .B(n733), .C(n4966), .D(n599), .Y(n5184) );
  NAND3X1 U5004 ( .A(n5192), .B(n153), .C(n55), .Y(n6334) );
  NAND2X1 U5005 ( .A(\mem<40><0> ), .B(n4680), .Y(n5168) );
  OAI21X1 U5006 ( .A(n4829), .B(n5169), .C(n5168), .Y(n5182) );
  NOR2X1 U5007 ( .A(n93), .B(n5170), .Y(n5181) );
  AND2X2 U5008 ( .A(\mem<62><0> ), .B(n4853), .Y(n5171) );
  AND2X2 U5009 ( .A(\mem<30><0> ), .B(n4853), .Y(n5172) );
  NAND3X1 U5010 ( .A(n1273), .B(n2356), .C(n4063), .Y(n5176) );
  NAND2X1 U5011 ( .A(\mem<46><0> ), .B(n150), .Y(n5173) );
  OAI21X1 U5012 ( .A(n4963), .B(n5174), .C(n5173), .Y(n5175) );
  OAI21X1 U5013 ( .A(n4953), .B(n5177), .C(n1138), .Y(n5178) );
  AOI21X1 U5014 ( .A(\mem<6><0> ), .B(n4838), .C(n5178), .Y(n5179) );
  AOI21X1 U5015 ( .A(n4055), .B(n5179), .C(n4834), .Y(n5180) );
  NOR3X1 U5016 ( .A(n5182), .B(n5181), .C(n3569), .Y(n5183) );
  NAND3X1 U5017 ( .A(n5183), .B(n5185), .C(n3095), .Y(n5186) );
  AOI22X1 U5018 ( .A(\mem<8><0> ), .B(n6402), .C(\mem<9><0> ), .D(n3863), .Y(
        n5197) );
  OAI21X1 U5019 ( .A(n6370), .B(n5189), .C(n5188), .Y(n5190) );
  AOI21X1 U5020 ( .A(\mem<4><0> ), .B(n6413), .C(n5190), .Y(n5196) );
  OAI21X1 U5021 ( .A(n806), .B(n5191), .C(n165), .Y(n5195) );
  OAI21X1 U5022 ( .A(n120), .B(n5193), .C(n3681), .Y(n5194) );
  AOI22X1 U5023 ( .A(\mem<32><0> ), .B(n804), .C(\mem<25><0> ), .D(n3856), .Y(
        n5209) );
  OAI21X1 U5024 ( .A(n4879), .B(n5202), .C(n167), .Y(n5206) );
  OAI21X1 U5025 ( .A(n3652), .B(n5204), .C(n3903), .Y(n5205) );
  NAND3X1 U5026 ( .A(n5209), .B(n5207), .C(n5208), .Y(n5210) );
  AOI21X1 U5027 ( .A(n1808), .B(n5211), .C(n4697), .Y(\data_out<0> ) );
  OAI21X1 U5028 ( .A(n6370), .B(n5213), .C(n5212), .Y(n5214) );
  AOI21X1 U5029 ( .A(\mem<4><1> ), .B(n6413), .C(n5214), .Y(n5220) );
  OAI21X1 U5030 ( .A(n6304), .B(n5215), .C(n169), .Y(n5218) );
  OAI21X1 U5031 ( .A(n3567), .B(n5216), .C(n3683), .Y(n5217) );
  AOI22X1 U5032 ( .A(\mem<32><1> ), .B(n804), .C(\mem<25><1> ), .D(n6368), .Y(
        n5230) );
  OAI21X1 U5033 ( .A(n4850), .B(n5223), .C(n5222), .Y(n5224) );
  AOI21X1 U5034 ( .A(\mem<26><1> ), .B(n6366), .C(n5224), .Y(n5229) );
  OAI21X1 U5035 ( .A(n4879), .B(n5225), .C(n171), .Y(n5228) );
  OAI21X1 U5036 ( .A(n3652), .B(n5226), .C(n3905), .Y(n5227) );
  NAND2X1 U5037 ( .A(\mem<20><1> ), .B(n6377), .Y(n5231) );
  OAI21X1 U5038 ( .A(n4887), .B(n5232), .C(n5231), .Y(n5233) );
  AOI21X1 U5039 ( .A(\mem<42><1> ), .B(n6331), .C(n5233), .Y(n5240) );
  AOI22X1 U5040 ( .A(\mem<58><1> ), .B(n84), .C(\mem<28><1> ), .D(n6363), .Y(
        n5239) );
  OAI21X1 U5041 ( .A(n6344), .B(n5234), .C(n1140), .Y(n5238) );
  NAND2X1 U5042 ( .A(\mem<18><1> ), .B(n4911), .Y(n5235) );
  OAI21X1 U5043 ( .A(n6342), .B(n5236), .C(n5235), .Y(n5237) );
  NOR2X1 U5044 ( .A(n138), .B(n5241), .Y(n5242) );
  AOI21X1 U5045 ( .A(\mem<11><1> ), .B(n4961), .C(n5242), .Y(n5249) );
  NAND2X1 U5046 ( .A(\mem<59><1> ), .B(n4946), .Y(n5244) );
  AND2X2 U5047 ( .A(\mem<27><1> ), .B(n4765), .Y(n5243) );
  OAI21X1 U5048 ( .A(n5244), .B(n4945), .C(n1142), .Y(n5245) );
  OAI21X1 U5049 ( .A(n4953), .B(n5246), .C(n3907), .Y(n5247) );
  AOI21X1 U5050 ( .A(\mem<3><1> ), .B(n4838), .C(n5247), .Y(n5248) );
  NOR2X1 U5051 ( .A(n4688), .B(n6421), .Y(n5250) );
  OAI21X1 U5052 ( .A(n3658), .B(n5251), .C(n3909), .Y(n5252) );
  AOI21X1 U5053 ( .A(n6415), .B(n618), .C(n5252), .Y(n5289) );
  NOR2X1 U5054 ( .A(n137), .B(n5253), .Y(n5254) );
  AOI21X1 U5055 ( .A(\mem<15><1> ), .B(n3847), .C(n5254), .Y(n5262) );
  NAND2X1 U5056 ( .A(\mem<63><1> ), .B(n4946), .Y(n5256) );
  AND2X2 U5057 ( .A(\mem<31><1> ), .B(n4853), .Y(n5255) );
  OAI21X1 U5058 ( .A(n5256), .B(n4945), .C(n1144), .Y(n5257) );
  AOI21X1 U5059 ( .A(\mem<23><1> ), .B(n4957), .C(n5257), .Y(n5261) );
  OAI21X1 U5060 ( .A(n4953), .B(n5258), .C(n3911), .Y(n5259) );
  AOI21X1 U5061 ( .A(\mem<7><1> ), .B(n4838), .C(n5259), .Y(n5260) );
  NOR2X1 U5062 ( .A(n135), .B(n5263), .Y(n5264) );
  AOI21X1 U5063 ( .A(\mem<13><1> ), .B(n4961), .C(n5264), .Y(n5272) );
  NAND2X1 U5064 ( .A(\mem<61><1> ), .B(n4946), .Y(n5266) );
  AND2X2 U5065 ( .A(\mem<29><1> ), .B(n4853), .Y(n5265) );
  OAI21X1 U5066 ( .A(n5266), .B(n113), .C(n1146), .Y(n5267) );
  AOI21X1 U5067 ( .A(\mem<21><1> ), .B(n4959), .C(n5267), .Y(n5271) );
  OAI21X1 U5068 ( .A(n4953), .B(n5268), .C(n3913), .Y(n5269) );
  AOI21X1 U5069 ( .A(\mem<5><1> ), .B(n4838), .C(n5269), .Y(n5270) );
  AOI22X1 U5070 ( .A(n4964), .B(n622), .C(n4967), .D(n627), .Y(n5288) );
  OAI21X1 U5071 ( .A(n4830), .B(n5273), .C(n173), .Y(n5286) );
  NOR2X1 U5072 ( .A(n93), .B(n5274), .Y(n5285) );
  AND2X2 U5073 ( .A(\mem<62><1> ), .B(n4765), .Y(n5275) );
  AND2X2 U5074 ( .A(\mem<30><1> ), .B(n4853), .Y(n5276) );
  NAND3X1 U5075 ( .A(n1275), .B(n2358), .C(n3098), .Y(n5280) );
  NAND2X1 U5076 ( .A(\mem<46><1> ), .B(n151), .Y(n5277) );
  OAI21X1 U5077 ( .A(n4673), .B(n5278), .C(n5277), .Y(n5279) );
  OAI21X1 U5078 ( .A(n4953), .B(n5281), .C(n3915), .Y(n5282) );
  AOI21X1 U5079 ( .A(\mem<6><1> ), .B(n4838), .C(n5282), .Y(n5283) );
  AOI21X1 U5080 ( .A(n4057), .B(n5283), .C(n4834), .Y(n5284) );
  NOR3X1 U5081 ( .A(n5286), .B(n5285), .C(n3570), .Y(n5287) );
  NAND2X1 U5082 ( .A(\mem<20><2> ), .B(n6377), .Y(n5291) );
  OAI21X1 U5083 ( .A(n4887), .B(n5292), .C(n5291), .Y(n5293) );
  AOI21X1 U5084 ( .A(\mem<42><2> ), .B(n6331), .C(n5293), .Y(n5299) );
  AOI22X1 U5085 ( .A(\mem<58><2> ), .B(n83), .C(\mem<28><2> ), .D(n6363), .Y(
        n5298) );
  OAI21X1 U5086 ( .A(n6344), .B(n5294), .C(n175), .Y(n5297) );
  OAI21X1 U5087 ( .A(n6342), .B(n5295), .C(n177), .Y(n5296) );
  NOR2X1 U5088 ( .A(n4951), .B(n5300), .Y(n5301) );
  AOI21X1 U5089 ( .A(\mem<11><2> ), .B(n4961), .C(n5301), .Y(n5309) );
  NAND2X1 U5090 ( .A(\mem<59><2> ), .B(n4946), .Y(n5303) );
  AND2X2 U5091 ( .A(\mem<27><2> ), .B(n4947), .Y(n5302) );
  OAI21X1 U5092 ( .A(n5303), .B(n4945), .C(n1148), .Y(n5304) );
  AOI21X1 U5093 ( .A(\mem<19><2> ), .B(n4959), .C(n5304), .Y(n5308) );
  OAI21X1 U5094 ( .A(n4953), .B(n5305), .C(n3917), .Y(n5306) );
  AOI21X1 U5095 ( .A(\mem<3><2> ), .B(n4838), .C(n5306), .Y(n5307) );
  NOR2X1 U5096 ( .A(n4687), .B(n6422), .Y(n5310) );
  OAI21X1 U5097 ( .A(n5649), .B(n5311), .C(n3919), .Y(n5312) );
  AOI21X1 U5098 ( .A(n6415), .B(n731), .C(n5312), .Y(n5352) );
  NOR2X1 U5099 ( .A(n135), .B(n5313), .Y(n5314) );
  NAND2X1 U5100 ( .A(\mem<63><2> ), .B(n4946), .Y(n5316) );
  AND2X2 U5101 ( .A(\mem<31><2> ), .B(n4947), .Y(n5315) );
  OAI21X1 U5102 ( .A(n5316), .B(n4945), .C(n1150), .Y(n5317) );
  AOI21X1 U5103 ( .A(\mem<23><2> ), .B(n4958), .C(n5317), .Y(n5322) );
  NAND2X1 U5104 ( .A(\mem<55><2> ), .B(n4948), .Y(n5318) );
  OAI21X1 U5105 ( .A(n4953), .B(n5319), .C(n5318), .Y(n5320) );
  AOI21X1 U5106 ( .A(\mem<7><2> ), .B(n4838), .C(n5320), .Y(n5321) );
  NOR2X1 U5107 ( .A(n4951), .B(n5324), .Y(n5325) );
  AOI21X1 U5108 ( .A(\mem<13><2> ), .B(n4962), .C(n5325), .Y(n5333) );
  NAND2X1 U5109 ( .A(\mem<61><2> ), .B(n4946), .Y(n5327) );
  AND2X2 U5110 ( .A(\mem<29><2> ), .B(n4947), .Y(n5326) );
  OAI21X1 U5111 ( .A(n5327), .B(n4945), .C(n1152), .Y(n5328) );
  AOI21X1 U5112 ( .A(\mem<21><2> ), .B(n4959), .C(n5328), .Y(n5332) );
  OAI21X1 U5113 ( .A(n4953), .B(n5329), .C(n3921), .Y(n5330) );
  AOI21X1 U5114 ( .A(\mem<5><2> ), .B(n4838), .C(n5330), .Y(n5331) );
  AOI22X1 U5115 ( .A(n4964), .B(n735), .C(n4966), .D(n637), .Y(n5351) );
  NAND2X1 U5116 ( .A(\mem<40><2> ), .B(n4680), .Y(n5334) );
  OAI21X1 U5117 ( .A(n4830), .B(n5335), .C(n5334), .Y(n5349) );
  NOR2X1 U5118 ( .A(n96), .B(n5336), .Y(n5348) );
  AND2X2 U5119 ( .A(\mem<62><2> ), .B(n4947), .Y(n5337) );
  AND2X2 U5120 ( .A(\mem<30><2> ), .B(n4947), .Y(n5338) );
  NAND3X1 U5121 ( .A(n1277), .B(n2360), .C(n4065), .Y(n5342) );
  NAND2X1 U5122 ( .A(\mem<46><2> ), .B(n149), .Y(n5339) );
  OAI21X1 U5123 ( .A(n4963), .B(n5340), .C(n5339), .Y(n5341) );
  NAND2X1 U5124 ( .A(\mem<54><2> ), .B(n4949), .Y(n5343) );
  OAI21X1 U5125 ( .A(n125), .B(n5344), .C(n5343), .Y(n5345) );
  AOI21X1 U5126 ( .A(\mem<6><2> ), .B(n4838), .C(n5345), .Y(n5346) );
  AOI21X1 U5127 ( .A(n4059), .B(n5346), .C(n4834), .Y(n5347) );
  NOR3X1 U5128 ( .A(n5349), .B(n5348), .C(n3571), .Y(n5350) );
  OAI21X1 U5129 ( .A(n566), .B(n5354), .C(n1132), .Y(n5355) );
  AOI21X1 U5130 ( .A(\mem<32><2> ), .B(n804), .C(n5355), .Y(n5362) );
  OAI21X1 U5131 ( .A(n4917), .B(n5356), .C(n796), .Y(n5359) );
  OAI21X1 U5132 ( .A(n3575), .B(n5357), .C(n1154), .Y(n5358) );
  NAND3X1 U5133 ( .A(n5362), .B(n5361), .C(n5360), .Y(n5373) );
  OAI21X1 U5134 ( .A(n4918), .B(n5363), .C(n1156), .Y(n5367) );
  NAND2X1 U5135 ( .A(\mem<8><2> ), .B(n6402), .Y(n5364) );
  OAI21X1 U5136 ( .A(n3669), .B(n5365), .C(n5364), .Y(n5366) );
  OAI21X1 U5137 ( .A(n6313), .B(n5368), .C(n156), .Y(n5372) );
  AOI22X1 U5138 ( .A(\mem<16><2> ), .B(n4816), .C(\mem<10><2> ), .D(n6399), 
        .Y(n5369) );
  OAI21X1 U5139 ( .A(n4879), .B(n5370), .C(n5369), .Y(n5371) );
  AOI21X1 U5140 ( .A(n795), .B(n5374), .C(n4697), .Y(\data_out<2> ) );
  NAND2X1 U5141 ( .A(\mem<17><3> ), .B(n6387), .Y(n5375) );
  OAI21X1 U5142 ( .A(n4719), .B(n5376), .C(n5375), .Y(n5380) );
  AOI22X1 U5143 ( .A(\mem<49><3> ), .B(n17), .C(\mem<33><3> ), .D(n4822), .Y(
        n5377) );
  OAI21X1 U5144 ( .A(n3862), .B(n5378), .C(n5377), .Y(n5379) );
  NAND2X1 U5145 ( .A(\mem<32><3> ), .B(n804), .Y(n5383) );
  OAI21X1 U5146 ( .A(n3578), .B(n5384), .C(n5383), .Y(n5385) );
  NOR2X1 U5147 ( .A(n134), .B(n5387), .Y(n5388) );
  AOI21X1 U5148 ( .A(\mem<11><3> ), .B(n4961), .C(n5388), .Y(n5397) );
  NAND2X1 U5149 ( .A(\mem<59><3> ), .B(n4946), .Y(n5390) );
  AND2X2 U5150 ( .A(\mem<27><3> ), .B(n4947), .Y(n5389) );
  OAI21X1 U5151 ( .A(n5390), .B(n4945), .C(n1158), .Y(n5391) );
  AOI21X1 U5152 ( .A(\mem<19><3> ), .B(n4957), .C(n5391), .Y(n5396) );
  NAND2X1 U5153 ( .A(\mem<51><3> ), .B(n4851), .Y(n5392) );
  OAI21X1 U5154 ( .A(n4953), .B(n5393), .C(n5392), .Y(n5394) );
  AOI21X1 U5155 ( .A(\mem<3><3> ), .B(n4838), .C(n5394), .Y(n5395) );
  NOR2X1 U5156 ( .A(n4689), .B(n6423), .Y(n5398) );
  OAI21X1 U5157 ( .A(n5649), .B(n5399), .C(n3923), .Y(n5400) );
  AOI21X1 U5158 ( .A(n6415), .B(n642), .C(n5400), .Y(n5437) );
  NOR2X1 U5159 ( .A(n134), .B(n5401), .Y(n5402) );
  AND2X2 U5160 ( .A(\mem<31><3> ), .B(n4947), .Y(n5403) );
  OAI21X1 U5161 ( .A(n305), .B(n4945), .C(n1160), .Y(n5404) );
  AOI21X1 U5162 ( .A(\mem<23><3> ), .B(n4958), .C(n5404), .Y(n5409) );
  NAND2X1 U5163 ( .A(\mem<55><3> ), .B(n4851), .Y(n5405) );
  OAI21X1 U5164 ( .A(n4955), .B(n5406), .C(n5405), .Y(n5407) );
  AOI21X1 U5165 ( .A(\mem<7><3> ), .B(n4838), .C(n5407), .Y(n5408) );
  NOR2X1 U5166 ( .A(n140), .B(n5411), .Y(n5412) );
  AOI21X1 U5167 ( .A(\mem<13><3> ), .B(n4961), .C(n5412), .Y(n5421) );
  NAND2X1 U5168 ( .A(\mem<61><3> ), .B(n4946), .Y(n5414) );
  AND2X2 U5169 ( .A(\mem<29><3> ), .B(n4947), .Y(n5413) );
  OAI21X1 U5170 ( .A(n5414), .B(n4945), .C(n1162), .Y(n5415) );
  AOI21X1 U5171 ( .A(\mem<21><3> ), .B(n4957), .C(n5415), .Y(n5420) );
  NAND2X1 U5172 ( .A(\mem<53><3> ), .B(n4848), .Y(n5416) );
  OAI21X1 U5173 ( .A(n125), .B(n5417), .C(n5416), .Y(n5418) );
  AOI21X1 U5174 ( .A(\mem<5><3> ), .B(n4838), .C(n5418), .Y(n5419) );
  AOI22X1 U5175 ( .A(n3661), .B(n647), .C(n4966), .D(n652), .Y(n5436) );
  NAND2X1 U5176 ( .A(\mem<25><3> ), .B(n4916), .Y(n5422) );
  OAI21X1 U5177 ( .A(n3881), .B(n5423), .C(n5422), .Y(n5434) );
  AND2X2 U5178 ( .A(\mem<62><3> ), .B(n4947), .Y(n5425) );
  NAND2X1 U5179 ( .A(\mem<30><3> ), .B(n4946), .Y(n5424) );
  AOI21X1 U5180 ( .A(n4944), .B(n5425), .C(n821), .Y(n5429) );
  NOR2X1 U5181 ( .A(n131), .B(n5426), .Y(n5427) );
  AOI21X1 U5182 ( .A(\mem<14><3> ), .B(n3847), .C(n5427), .Y(n5428) );
  NAND3X1 U5183 ( .A(n1266), .B(n3721), .C(n5428), .Y(n5430) );
  OAI21X1 U5184 ( .A(n4862), .B(n5432), .C(n5431), .Y(n5433) );
  NAND3X1 U5185 ( .A(n3687), .B(n2347), .C(n5435), .Y(n5438) );
  OAI21X1 U5186 ( .A(n6342), .B(n5440), .C(n1164), .Y(n5441) );
  AOI21X1 U5187 ( .A(\mem<28><3> ), .B(n6363), .C(n5441), .Y(n5449) );
  AOI21X1 U5188 ( .A(\mem<60><3> ), .B(n3665), .C(n5442), .Y(n5448) );
  OAI21X1 U5189 ( .A(n815), .B(n5444), .C(n5443), .Y(n5447) );
  INVX2 U5190 ( .A(\mem<20><3> ), .Y(n5445) );
  OAI21X1 U5191 ( .A(n3662), .B(n5445), .C(n3925), .Y(n5446) );
  NAND2X1 U5192 ( .A(\mem<24><3> ), .B(n3867), .Y(n5450) );
  OAI21X1 U5193 ( .A(n6414), .B(n5451), .C(n5450), .Y(n5452) );
  INVX2 U5194 ( .A(n4878), .Y(n6416) );
  AOI22X1 U5195 ( .A(\mem<10><3> ), .B(n6399), .C(\mem<2><3> ), .D(n6416), .Y(
        n5459) );
  NAND2X1 U5196 ( .A(\mem<18><3> ), .B(n577), .Y(n5453) );
  OAI21X1 U5197 ( .A(n6344), .B(n5454), .C(n5453), .Y(n5458) );
  NAND2X1 U5198 ( .A(\mem<44><3> ), .B(n4868), .Y(n5455) );
  AOI21X1 U5199 ( .A(n1810), .B(n764), .C(n4697), .Y(\data_out<3> ) );
  AOI21X1 U5200 ( .A(\mem<33><4> ), .B(n4844), .C(n5462), .Y(n5471) );
  NAND2X1 U5201 ( .A(\mem<52><4> ), .B(n4876), .Y(n5463) );
  OAI21X1 U5202 ( .A(n3669), .B(n5464), .C(n5463), .Y(n5468) );
  NAND2X1 U5203 ( .A(\mem<32><4> ), .B(n804), .Y(n5465) );
  OAI21X1 U5204 ( .A(n3578), .B(n5466), .C(n5465), .Y(n5467) );
  NOR2X1 U5205 ( .A(n131), .B(n5472), .Y(n5473) );
  AOI21X1 U5206 ( .A(\mem<11><4> ), .B(n4961), .C(n5473), .Y(n5481) );
  NAND2X1 U5207 ( .A(\mem<59><4> ), .B(n4946), .Y(n5475) );
  AND2X2 U5208 ( .A(\mem<27><4> ), .B(n4947), .Y(n5474) );
  OAI21X1 U5209 ( .A(n5475), .B(n4945), .C(n1166), .Y(n5476) );
  AOI21X1 U5210 ( .A(\mem<19><4> ), .B(n4957), .C(n5476), .Y(n5480) );
  OAI21X1 U5211 ( .A(n4953), .B(n5477), .C(n3927), .Y(n5478) );
  AOI21X1 U5212 ( .A(\mem<3><4> ), .B(n4838), .C(n5478), .Y(n5479) );
  NOR2X1 U5213 ( .A(n4690), .B(n6424), .Y(n5482) );
  OAI21X1 U5214 ( .A(n3658), .B(n5483), .C(n3929), .Y(n5484) );
  AOI21X1 U5215 ( .A(n6415), .B(n660), .C(n5484), .Y(n5517) );
  NOR2X1 U5216 ( .A(n4951), .B(n5485), .Y(n5486) );
  AOI21X1 U5217 ( .A(\mem<15><4> ), .B(n4961), .C(n5486), .Y(n5494) );
  NAND2X1 U5218 ( .A(\mem<63><4> ), .B(n4946), .Y(n5488) );
  AND2X2 U5219 ( .A(\mem<31><4> ), .B(n4947), .Y(n5487) );
  OAI21X1 U5220 ( .A(n5488), .B(n4945), .C(n1168), .Y(n5489) );
  NAND2X1 U5221 ( .A(\mem<55><4> ), .B(n4949), .Y(n5490) );
  OAI21X1 U5222 ( .A(n4953), .B(n5491), .C(n5490), .Y(n5492) );
  AOI21X1 U5223 ( .A(\mem<7><4> ), .B(n4838), .C(n5492), .Y(n5493) );
  NOR2X1 U5224 ( .A(n140), .B(n5495), .Y(n5496) );
  AOI21X1 U5225 ( .A(\mem<13><4> ), .B(n4962), .C(n5496), .Y(n5504) );
  NAND2X1 U5226 ( .A(\mem<61><4> ), .B(n4946), .Y(n5498) );
  AND2X2 U5227 ( .A(\mem<29><4> ), .B(n4947), .Y(n5497) );
  OAI21X1 U5228 ( .A(n5498), .B(n4945), .C(n1170), .Y(n5499) );
  AOI21X1 U5229 ( .A(\mem<21><4> ), .B(n4957), .C(n5499), .Y(n5503) );
  OAI21X1 U5230 ( .A(n4953), .B(n5500), .C(n3931), .Y(n5501) );
  AOI21X1 U5231 ( .A(\mem<5><4> ), .B(n4838), .C(n5501), .Y(n5502) );
  AOI22X1 U5232 ( .A(n4964), .B(n737), .C(n4966), .D(n665), .Y(n5516) );
  NAND2X1 U5233 ( .A(\mem<25><4> ), .B(n3564), .Y(n5505) );
  AND2X2 U5234 ( .A(\mem<62><4> ), .B(n4947), .Y(n5508) );
  NAND2X1 U5235 ( .A(\mem<30><4> ), .B(n4946), .Y(n5507) );
  AOI21X1 U5236 ( .A(n4944), .B(n5508), .C(n823), .Y(n5512) );
  NOR2X1 U5237 ( .A(n138), .B(n5509), .Y(n5510) );
  AOI21X1 U5238 ( .A(\mem<14><4> ), .B(n3847), .C(n5510), .Y(n5511) );
  NAND3X1 U5239 ( .A(n1267), .B(n3723), .C(n5511), .Y(n5513) );
  NAND3X1 U5240 ( .A(n1265), .B(n2351), .C(n5515), .Y(n5518) );
  OAI21X1 U5241 ( .A(n6342), .B(n5520), .C(n1172), .Y(n5521) );
  AOI21X1 U5242 ( .A(\mem<28><4> ), .B(n6363), .C(n5521), .Y(n5530) );
  OAI21X1 U5243 ( .A(n6378), .B(n5524), .C(n3933), .Y(n5525) );
  NOR2X1 U5244 ( .A(n6332), .B(n5527), .Y(n5528) );
  AOI21X1 U5245 ( .A(\mem<60><4> ), .B(n3665), .C(n5528), .Y(n5529) );
  OAI21X1 U5246 ( .A(n6414), .B(n5531), .C(n68), .Y(n5532) );
  NAND2X1 U5247 ( .A(\mem<18><4> ), .B(n4911), .Y(n5533) );
  OAI21X1 U5248 ( .A(n6344), .B(n5534), .C(n5533), .Y(n5537) );
  AOI22X1 U5249 ( .A(\mem<10><4> ), .B(n6399), .C(\mem<2><4> ), .D(n6416), .Y(
        n5538) );
  AOI21X1 U5250 ( .A(n790), .B(n5541), .C(n4697), .Y(\data_out<4> ) );
  NAND2X1 U5251 ( .A(\mem<49><5> ), .B(n4835), .Y(n5542) );
  OAI21X1 U5252 ( .A(n3862), .B(n5543), .C(n5542), .Y(n5544) );
  NAND2X1 U5253 ( .A(\mem<52><5> ), .B(n4875), .Y(n5545) );
  OAI21X1 U5254 ( .A(n3669), .B(n5546), .C(n5545), .Y(n5550) );
  NAND2X1 U5255 ( .A(\mem<32><5> ), .B(n804), .Y(n5547) );
  OAI21X1 U5256 ( .A(n3578), .B(n5548), .C(n5547), .Y(n5549) );
  NOR2X1 U5257 ( .A(n13), .B(n5551), .Y(n5552) );
  AOI21X1 U5258 ( .A(\mem<56><5> ), .B(n4682), .C(n5552), .Y(n5553) );
  NOR2X1 U5259 ( .A(n141), .B(n5555), .Y(n5556) );
  AOI21X1 U5260 ( .A(\mem<11><5> ), .B(n4962), .C(n5556), .Y(n5564) );
  NAND2X1 U5261 ( .A(\mem<59><5> ), .B(n4946), .Y(n5558) );
  AND2X2 U5262 ( .A(\mem<27><5> ), .B(n4947), .Y(n5557) );
  OAI21X1 U5263 ( .A(n5558), .B(n4945), .C(n1176), .Y(n5559) );
  AOI21X1 U5264 ( .A(\mem<19><5> ), .B(n4957), .C(n5559), .Y(n5563) );
  OAI21X1 U5265 ( .A(n4953), .B(n5560), .C(n3935), .Y(n5561) );
  AOI21X1 U5266 ( .A(\mem<3><5> ), .B(n4838), .C(n5561), .Y(n5562) );
  NOR2X1 U5267 ( .A(n4688), .B(n6425), .Y(n5565) );
  OAI21X1 U5268 ( .A(n3658), .B(n5566), .C(n3937), .Y(n5567) );
  AOI21X1 U5269 ( .A(n6415), .B(n678), .C(n5567), .Y(n5602) );
  NOR2X1 U5270 ( .A(n129), .B(n5568), .Y(n5569) );
  AOI21X1 U5271 ( .A(\mem<15><5> ), .B(n4961), .C(n5569), .Y(n5578) );
  NAND2X1 U5272 ( .A(\mem<63><5> ), .B(n4946), .Y(n5571) );
  AND2X2 U5273 ( .A(\mem<31><5> ), .B(n4947), .Y(n5570) );
  OAI21X1 U5274 ( .A(n5571), .B(n58), .C(n1178), .Y(n5572) );
  AOI21X1 U5275 ( .A(\mem<23><5> ), .B(n4957), .C(n5572), .Y(n5577) );
  NAND2X1 U5276 ( .A(\mem<55><5> ), .B(n4948), .Y(n5573) );
  OAI21X1 U5277 ( .A(n4953), .B(n5574), .C(n5573), .Y(n5575) );
  AOI21X1 U5278 ( .A(\mem<7><5> ), .B(n4838), .C(n5575), .Y(n5576) );
  NOR2X1 U5279 ( .A(n130), .B(n5579), .Y(n5580) );
  AOI21X1 U5280 ( .A(\mem<13><5> ), .B(n4961), .C(n5580), .Y(n5588) );
  NAND2X1 U5281 ( .A(\mem<61><5> ), .B(n4946), .Y(n5582) );
  AND2X2 U5282 ( .A(\mem<29><5> ), .B(n4947), .Y(n5581) );
  OAI21X1 U5283 ( .A(n5582), .B(n113), .C(n1180), .Y(n5583) );
  AOI21X1 U5284 ( .A(\mem<21><5> ), .B(n4957), .C(n5583), .Y(n5587) );
  OAI21X1 U5285 ( .A(n4953), .B(n5584), .C(n3939), .Y(n5585) );
  AOI21X1 U5286 ( .A(\mem<5><5> ), .B(n4838), .C(n5585), .Y(n5586) );
  AOI22X1 U5287 ( .A(n4964), .B(n739), .C(n4966), .D(n683), .Y(n5601) );
  AND2X2 U5288 ( .A(\mem<62><5> ), .B(n4947), .Y(n5592) );
  NAND2X1 U5289 ( .A(\mem<30><5> ), .B(n4946), .Y(n5591) );
  AOI21X1 U5290 ( .A(n4944), .B(n5592), .C(n825), .Y(n5594) );
  AOI21X1 U5291 ( .A(\mem<14><5> ), .B(n3847), .C(n4625), .Y(n5593) );
  NAND3X1 U5292 ( .A(n1269), .B(n3725), .C(n5593), .Y(n5595) );
  NAND3X1 U5293 ( .A(n1268), .B(n2348), .C(n5600), .Y(n5603) );
  OAI21X1 U5294 ( .A(n6342), .B(n5605), .C(n1182), .Y(n5606) );
  AOI21X1 U5295 ( .A(\mem<28><5> ), .B(n6363), .C(n5606), .Y(n5615) );
  NAND2X1 U5296 ( .A(\mem<12><5> ), .B(n3654), .Y(n5607) );
  OAI21X1 U5297 ( .A(n6378), .B(n5609), .C(n1184), .Y(n5610) );
  NOR2X1 U5298 ( .A(n6332), .B(n5612), .Y(n5613) );
  AOI21X1 U5299 ( .A(\mem<60><5> ), .B(n3665), .C(n5613), .Y(n5614) );
  NAND2X1 U5300 ( .A(\mem<24><5> ), .B(n3868), .Y(n5616) );
  OAI21X1 U5301 ( .A(n6414), .B(n5617), .C(n5616), .Y(n5618) );
  AOI21X1 U5302 ( .A(\mem<16><5> ), .B(n4816), .C(n5618), .Y(n5626) );
  NAND2X1 U5303 ( .A(\mem<18><5> ), .B(n4911), .Y(n5619) );
  OAI21X1 U5304 ( .A(n6344), .B(n5620), .C(n5619), .Y(n5623) );
  AOI22X1 U5305 ( .A(\mem<10><5> ), .B(n6399), .C(\mem<2><5> ), .D(n6416), .Y(
        n5624) );
  AOI21X1 U5306 ( .A(n1812), .B(n769), .C(n4697), .Y(\data_out<5> ) );
  OAI21X1 U5307 ( .A(n4677), .B(n5627), .C(n71), .Y(n5628) );
  OAI21X1 U5308 ( .A(n3669), .B(n5629), .C(n1188), .Y(n5633) );
  NAND2X1 U5309 ( .A(\mem<32><6> ), .B(n804), .Y(n5630) );
  OAI21X1 U5310 ( .A(n3578), .B(n5631), .C(n5630), .Y(n5632) );
  NOR2X1 U5311 ( .A(n138), .B(n5637), .Y(n5638) );
  AOI21X1 U5312 ( .A(\mem<11><6> ), .B(n4961), .C(n5638), .Y(n5646) );
  AND2X2 U5313 ( .A(\mem<27><6> ), .B(n4947), .Y(n5639) );
  OAI21X1 U5314 ( .A(n307), .B(n113), .C(n1190), .Y(n5640) );
  AOI21X1 U5315 ( .A(\mem<19><6> ), .B(n4957), .C(n5640), .Y(n5645) );
  NAND2X1 U5316 ( .A(\mem<51><6> ), .B(n4848), .Y(n5641) );
  OAI21X1 U5317 ( .A(n4953), .B(n5642), .C(n5641), .Y(n5643) );
  AOI21X1 U5318 ( .A(\mem<3><6> ), .B(n4838), .C(n5643), .Y(n5644) );
  NOR2X1 U5319 ( .A(n4687), .B(n6426), .Y(n5647) );
  OAI21X1 U5320 ( .A(n3658), .B(n5648), .C(n3941), .Y(n5650) );
  AOI21X1 U5321 ( .A(n6415), .B(n691), .C(n5650), .Y(n5685) );
  NOR2X1 U5322 ( .A(n142), .B(n5651), .Y(n5652) );
  AOI21X1 U5323 ( .A(\mem<15><6> ), .B(n4961), .C(n5652), .Y(n5660) );
  AND2X2 U5324 ( .A(\mem<31><6> ), .B(n4853), .Y(n5653) );
  OAI21X1 U5325 ( .A(n2330), .B(n113), .C(n3943), .Y(n5654) );
  AOI21X1 U5326 ( .A(\mem<23><6> ), .B(n4957), .C(n5654), .Y(n5659) );
  NAND2X1 U5327 ( .A(\mem<55><6> ), .B(n4949), .Y(n5655) );
  OAI21X1 U5328 ( .A(n4953), .B(n5656), .C(n5655), .Y(n5657) );
  AOI21X1 U5329 ( .A(\mem<7><6> ), .B(n4838), .C(n5657), .Y(n5658) );
  NOR2X1 U5330 ( .A(n137), .B(n5661), .Y(n5662) );
  AOI21X1 U5331 ( .A(\mem<13><6> ), .B(n4961), .C(n5662), .Y(n5669) );
  AND2X2 U5332 ( .A(\mem<29><6> ), .B(n4853), .Y(n5663) );
  OAI21X1 U5333 ( .A(n2332), .B(n113), .C(n3945), .Y(n5664) );
  NAND2X1 U5334 ( .A(\mem<53><6> ), .B(n4848), .Y(n5665) );
  OAI21X1 U5335 ( .A(n4953), .B(n5666), .C(n5665), .Y(n5667) );
  AOI21X1 U5336 ( .A(\mem<5><6> ), .B(n4838), .C(n5667), .Y(n5668) );
  AOI22X1 U5337 ( .A(n4964), .B(n741), .C(n4966), .D(n696), .Y(n5684) );
  NAND2X1 U5338 ( .A(\mem<25><6> ), .B(n4916), .Y(n5670) );
  AND2X2 U5339 ( .A(\mem<62><6> ), .B(n4853), .Y(n5673) );
  NAND2X1 U5340 ( .A(\mem<30><6> ), .B(n4946), .Y(n5672) );
  AOI21X1 U5341 ( .A(n4944), .B(n5673), .C(n827), .Y(n5677) );
  NOR2X1 U5342 ( .A(n133), .B(n5674), .Y(n5675) );
  AOI21X1 U5343 ( .A(\mem<14><6> ), .B(n3847), .C(n5675), .Y(n5676) );
  NAND3X1 U5344 ( .A(n1271), .B(n3727), .C(n5676), .Y(n5678) );
  NAND3X1 U5345 ( .A(n1270), .B(n5683), .C(n2349), .Y(n5686) );
  OAI21X1 U5346 ( .A(n6342), .B(n5688), .C(n1192), .Y(n5689) );
  AOI21X1 U5347 ( .A(\mem<28><6> ), .B(n6363), .C(n5689), .Y(n5698) );
  NAND2X1 U5348 ( .A(\mem<12><6> ), .B(n3654), .Y(n5690) );
  OAI21X1 U5349 ( .A(n93), .B(n5691), .C(n5690), .Y(n5694) );
  OAI21X1 U5350 ( .A(n6378), .B(n5692), .C(n1194), .Y(n5693) );
  NOR2X1 U5351 ( .A(n6332), .B(n5695), .Y(n5696) );
  AOI21X1 U5352 ( .A(\mem<60><6> ), .B(n3665), .C(n5696), .Y(n5697) );
  NAND2X1 U5353 ( .A(\mem<24><6> ), .B(n3868), .Y(n5699) );
  OAI21X1 U5354 ( .A(n6414), .B(n5700), .C(n5699), .Y(n5701) );
  AOI21X1 U5355 ( .A(\mem<16><6> ), .B(n4816), .C(n5701), .Y(n5709) );
  NAND2X1 U5356 ( .A(\mem<18><6> ), .B(n4911), .Y(n5702) );
  OAI21X1 U5357 ( .A(n6344), .B(n5703), .C(n5702), .Y(n5707) );
  NAND2X1 U5358 ( .A(\mem<44><6> ), .B(n574), .Y(n5704) );
  OAI21X1 U5359 ( .A(n3849), .B(n5705), .C(n5704), .Y(n5706) );
  AOI22X1 U5360 ( .A(\mem<10><6> ), .B(n6399), .C(\mem<2><6> ), .D(n6416), .Y(
        n5708) );
  AOI21X1 U5361 ( .A(n791), .B(n5710), .C(n4697), .Y(\data_out<6> ) );
  NAND2X1 U5362 ( .A(\mem<52><7> ), .B(n4876), .Y(n5711) );
  OAI21X1 U5363 ( .A(n3669), .B(n5712), .C(n5711), .Y(n5716) );
  NAND2X1 U5364 ( .A(\mem<32><7> ), .B(n804), .Y(n5713) );
  OAI21X1 U5365 ( .A(n3578), .B(n5714), .C(n5713), .Y(n5715) );
  AOI21X1 U5366 ( .A(\mem<17><7> ), .B(n6387), .C(n5717), .Y(n5722) );
  NAND2X1 U5367 ( .A(\mem<49><7> ), .B(n4813), .Y(n5718) );
  OAI21X1 U5368 ( .A(n4677), .B(n5719), .C(n5718), .Y(n5720) );
  AOI21X1 U5369 ( .A(\mem<33><7> ), .B(n4844), .C(n5720), .Y(n5721) );
  NAND2X1 U5370 ( .A(\mem<11><7> ), .B(n4962), .Y(n5723) );
  NAND3X1 U5371 ( .A(\mem<27><7> ), .B(n4946), .C(n4896), .Y(n5725) );
  NAND3X1 U5372 ( .A(\mem<59><7> ), .B(n4946), .C(n4944), .Y(n5724) );
  NOR3X1 U5373 ( .A(n743), .B(n713), .C(n830), .Y(n5728) );
  NOR2X1 U5374 ( .A(n4690), .B(n6428), .Y(n5726) );
  OAI21X1 U5375 ( .A(n4675), .B(n5728), .C(n5727), .Y(n5760) );
  NAND2X1 U5376 ( .A(\mem<63><7> ), .B(n4947), .Y(n5730) );
  NAND3X1 U5377 ( .A(\mem<31><7> ), .B(n4946), .C(n4891), .Y(n5729) );
  OAI21X1 U5378 ( .A(n5730), .B(n4943), .C(n5729), .Y(n5731) );
  AOI21X1 U5379 ( .A(\mem<23><7> ), .B(n4959), .C(n5731), .Y(n5737) );
  NAND2X1 U5380 ( .A(\mem<55><7> ), .B(n4949), .Y(n5732) );
  OAI21X1 U5381 ( .A(n4953), .B(n5733), .C(n5732), .Y(n5734) );
  AOI21X1 U5382 ( .A(\mem<7><7> ), .B(n4971), .C(n5734), .Y(n5736) );
  AOI22X1 U5383 ( .A(\mem<47><7> ), .B(n152), .C(\mem<15><7> ), .D(n4961), .Y(
        n5735) );
  NAND2X1 U5384 ( .A(\mem<61><7> ), .B(n4946), .Y(n5739) );
  NAND3X1 U5385 ( .A(\mem<29><7> ), .B(n4946), .C(n4893), .Y(n5738) );
  OAI21X1 U5386 ( .A(n5739), .B(n113), .C(n5738), .Y(n5740) );
  AOI21X1 U5387 ( .A(\mem<21><7> ), .B(n4959), .C(n5740), .Y(n5745) );
  OAI21X1 U5388 ( .A(n4953), .B(n5741), .C(n179), .Y(n5742) );
  AOI21X1 U5389 ( .A(\mem<5><7> ), .B(n4970), .C(n5742), .Y(n5744) );
  AOI22X1 U5390 ( .A(\mem<45><7> ), .B(n149), .C(\mem<13><7> ), .D(n4962), .Y(
        n5743) );
  NAND2X1 U5391 ( .A(\mem<25><7> ), .B(n6368), .Y(n5746) );
  OAI21X1 U5392 ( .A(n3881), .B(n5747), .C(n5746), .Y(n5757) );
  NAND2X1 U5393 ( .A(\mem<30><7> ), .B(n4946), .Y(n5750) );
  NAND3X1 U5394 ( .A(\mem<62><7> ), .B(n4765), .C(n4944), .Y(n5749) );
  OAI21X1 U5395 ( .A(n5750), .B(n4908), .C(n5749), .Y(n5753) );
  NAND3X1 U5396 ( .A(n181), .B(n4071), .C(n3959), .Y(n5752) );
  NAND2X1 U5397 ( .A(\mem<54><7> ), .B(n4949), .Y(n5754) );
  AOI21X1 U5398 ( .A(n153), .B(\mem<38><7> ), .C(n1263), .Y(n5755) );
  AOI21X1 U5399 ( .A(n1814), .B(n5755), .C(n4834), .Y(n5756) );
  NAND3X1 U5400 ( .A(n3957), .B(n4069), .C(n5758), .Y(n5759) );
  OAI21X1 U5401 ( .A(n6378), .B(n5763), .C(n3947), .Y(n5764) );
  AND2X2 U5402 ( .A(\mem<60><7> ), .B(n3665), .Y(n5766) );
  OAI21X1 U5403 ( .A(n6342), .B(n5767), .C(n1196), .Y(n5768) );
  AOI21X1 U5404 ( .A(\mem<28><7> ), .B(n6363), .C(n5768), .Y(n5769) );
  NAND2X1 U5405 ( .A(\mem<44><7> ), .B(n574), .Y(n5773) );
  AOI22X1 U5406 ( .A(\mem<2><7> ), .B(n6416), .C(\mem<10><7> ), .D(n6399), .Y(
        n5781) );
  NAND2X1 U5407 ( .A(\mem<24><7> ), .B(n3868), .Y(n5777) );
  OAI21X1 U5408 ( .A(n6414), .B(n5778), .C(n5777), .Y(n5779) );
  AOI21X1 U5409 ( .A(\mem<16><7> ), .B(n4816), .C(n5779), .Y(n5780) );
  AOI21X1 U5410 ( .A(n5782), .B(n763), .C(n4697), .Y(\data_out<7> ) );
  MUX2X1 U5411 ( .B(\mem<0><0> ), .A(\mem<32><0> ), .S(n5033), .Y(n5784) );
  MUX2X1 U5412 ( .B(\mem<2><0> ), .A(\mem<34><0> ), .S(n5033), .Y(n5783) );
  MUX2X1 U5413 ( .B(n5784), .A(n5783), .S(n4992), .Y(n5788) );
  MUX2X1 U5414 ( .B(\mem<4><0> ), .A(\mem<36><0> ), .S(n5033), .Y(n5786) );
  MUX2X1 U5415 ( .B(\mem<6><0> ), .A(\mem<38><0> ), .S(n5033), .Y(n5785) );
  MUX2X1 U5416 ( .B(n5786), .A(n5785), .S(n4992), .Y(n5787) );
  MUX2X1 U5417 ( .B(n5788), .A(n5787), .S(n5002), .Y(n5796) );
  MUX2X1 U5418 ( .B(\mem<8><0> ), .A(\mem<40><0> ), .S(n5033), .Y(n5790) );
  MUX2X1 U5419 ( .B(\mem<10><0> ), .A(\mem<42><0> ), .S(n5033), .Y(n5789) );
  MUX2X1 U5420 ( .B(n5790), .A(n5789), .S(n4992), .Y(n5794) );
  MUX2X1 U5421 ( .B(\mem<12><0> ), .A(\mem<44><0> ), .S(n5033), .Y(n5792) );
  MUX2X1 U5422 ( .B(\mem<14><0> ), .A(\mem<46><0> ), .S(n5032), .Y(n5791) );
  MUX2X1 U5423 ( .B(n5792), .A(n5791), .S(n4992), .Y(n5793) );
  MUX2X1 U5424 ( .B(n5794), .A(n5793), .S(n5002), .Y(n5795) );
  MUX2X1 U5425 ( .B(n5796), .A(n5795), .S(n5008), .Y(n5812) );
  MUX2X1 U5426 ( .B(\mem<16><0> ), .A(\mem<48><0> ), .S(n5032), .Y(n5798) );
  MUX2X1 U5427 ( .B(\mem<18><0> ), .A(\mem<50><0> ), .S(n5032), .Y(n5797) );
  MUX2X1 U5428 ( .B(n5798), .A(n5797), .S(n4992), .Y(n5802) );
  MUX2X1 U5429 ( .B(\mem<20><0> ), .A(\mem<52><0> ), .S(n5032), .Y(n5800) );
  MUX2X1 U5430 ( .B(\mem<22><0> ), .A(\mem<54><0> ), .S(n5032), .Y(n5799) );
  MUX2X1 U5431 ( .B(n5800), .A(n5799), .S(n4992), .Y(n5801) );
  MUX2X1 U5432 ( .B(n5802), .A(n5801), .S(n5002), .Y(n5810) );
  MUX2X1 U5433 ( .B(\mem<24><0> ), .A(\mem<56><0> ), .S(n5032), .Y(n5804) );
  MUX2X1 U5434 ( .B(\mem<26><0> ), .A(\mem<58><0> ), .S(n5032), .Y(n5803) );
  MUX2X1 U5435 ( .B(n5804), .A(n5803), .S(n4992), .Y(n5808) );
  MUX2X1 U5436 ( .B(\mem<28><0> ), .A(\mem<60><0> ), .S(n5032), .Y(n5806) );
  MUX2X1 U5437 ( .B(\mem<30><0> ), .A(\mem<62><0> ), .S(n5032), .Y(n5805) );
  MUX2X1 U5438 ( .B(n5806), .A(n5805), .S(n4992), .Y(n5807) );
  MUX2X1 U5439 ( .B(n5808), .A(n5807), .S(n5002), .Y(n5809) );
  MUX2X1 U5440 ( .B(n5810), .A(n5809), .S(n5008), .Y(n5811) );
  MUX2X1 U5441 ( .B(n5812), .A(n5811), .S(n5017), .Y(n5844) );
  MUX2X1 U5442 ( .B(\mem<1><0> ), .A(\mem<33><0> ), .S(n5032), .Y(n5814) );
  MUX2X1 U5443 ( .B(\mem<3><0> ), .A(\mem<35><0> ), .S(n5032), .Y(n5813) );
  MUX2X1 U5444 ( .B(n5814), .A(n5813), .S(n4991), .Y(n5818) );
  MUX2X1 U5445 ( .B(\mem<5><0> ), .A(\mem<37><0> ), .S(n5032), .Y(n5816) );
  MUX2X1 U5446 ( .B(\mem<7><0> ), .A(\mem<39><0> ), .S(n5031), .Y(n5815) );
  MUX2X1 U5447 ( .B(n5816), .A(n5815), .S(n4991), .Y(n5817) );
  MUX2X1 U5448 ( .B(n5818), .A(n5817), .S(n5001), .Y(n5826) );
  MUX2X1 U5449 ( .B(\mem<9><0> ), .A(\mem<41><0> ), .S(n5031), .Y(n5820) );
  MUX2X1 U5450 ( .B(\mem<11><0> ), .A(\mem<43><0> ), .S(n5031), .Y(n5819) );
  MUX2X1 U5451 ( .B(n5820), .A(n5819), .S(n4991), .Y(n5824) );
  MUX2X1 U5452 ( .B(\mem<13><0> ), .A(\mem<45><0> ), .S(n5031), .Y(n5822) );
  MUX2X1 U5453 ( .B(\mem<15><0> ), .A(\mem<47><0> ), .S(n5031), .Y(n5821) );
  MUX2X1 U5454 ( .B(n5822), .A(n5821), .S(n4991), .Y(n5823) );
  MUX2X1 U5455 ( .B(n5824), .A(n5823), .S(n5001), .Y(n5825) );
  MUX2X1 U5456 ( .B(n5826), .A(n5825), .S(n5008), .Y(n5842) );
  MUX2X1 U5457 ( .B(\mem<17><0> ), .A(\mem<49><0> ), .S(n5031), .Y(n5828) );
  MUX2X1 U5458 ( .B(\mem<19><0> ), .A(\mem<51><0> ), .S(n5031), .Y(n5827) );
  MUX2X1 U5459 ( .B(n5828), .A(n5827), .S(n4991), .Y(n5832) );
  MUX2X1 U5460 ( .B(\mem<21><0> ), .A(\mem<53><0> ), .S(n5031), .Y(n5830) );
  MUX2X1 U5461 ( .B(\mem<23><0> ), .A(\mem<55><0> ), .S(n5031), .Y(n5829) );
  MUX2X1 U5462 ( .B(n5830), .A(n5829), .S(n4991), .Y(n5831) );
  MUX2X1 U5463 ( .B(n5832), .A(n5831), .S(n5001), .Y(n5840) );
  MUX2X1 U5464 ( .B(\mem<25><0> ), .A(\mem<57><0> ), .S(n5031), .Y(n5834) );
  MUX2X1 U5465 ( .B(\mem<27><0> ), .A(\mem<59><0> ), .S(n5031), .Y(n5833) );
  MUX2X1 U5466 ( .B(n5834), .A(n5833), .S(n4991), .Y(n5838) );
  MUX2X1 U5467 ( .B(\mem<29><0> ), .A(\mem<61><0> ), .S(n5031), .Y(n5836) );
  MUX2X1 U5468 ( .B(\mem<31><0> ), .A(\mem<63><0> ), .S(n5029), .Y(n5835) );
  MUX2X1 U5469 ( .B(n5836), .A(n5835), .S(n4991), .Y(n5837) );
  MUX2X1 U5470 ( .B(n5838), .A(n5837), .S(n5001), .Y(n5839) );
  MUX2X1 U5471 ( .B(n5840), .A(n5839), .S(n5008), .Y(n5841) );
  MUX2X1 U5472 ( .B(n5842), .A(n5841), .S(n5017), .Y(n5843) );
  MUX2X1 U5473 ( .B(n5844), .A(n5843), .S(n114), .Y(n5845) );
  AND2X2 U5474 ( .A(n5845), .B(n5846), .Y(\data_out<8> ) );
  MUX2X1 U5475 ( .B(\mem<0><1> ), .A(\mem<32><1> ), .S(n5025), .Y(n5848) );
  MUX2X1 U5476 ( .B(\mem<2><1> ), .A(\mem<34><1> ), .S(n5030), .Y(n5847) );
  MUX2X1 U5477 ( .B(n5848), .A(n5847), .S(n4991), .Y(n5852) );
  MUX2X1 U5478 ( .B(\mem<4><1> ), .A(\mem<36><1> ), .S(n5029), .Y(n5850) );
  MUX2X1 U5479 ( .B(\mem<6><1> ), .A(\mem<38><1> ), .S(n5029), .Y(n5849) );
  MUX2X1 U5480 ( .B(n5850), .A(n5849), .S(n4991), .Y(n5851) );
  MUX2X1 U5481 ( .B(n5852), .A(n5851), .S(n5001), .Y(n5860) );
  MUX2X1 U5482 ( .B(\mem<8><1> ), .A(\mem<40><1> ), .S(n5030), .Y(n5854) );
  MUX2X1 U5483 ( .B(\mem<10><1> ), .A(\mem<42><1> ), .S(n5030), .Y(n5853) );
  MUX2X1 U5484 ( .B(n5854), .A(n5853), .S(n4991), .Y(n5858) );
  MUX2X1 U5485 ( .B(\mem<12><1> ), .A(\mem<44><1> ), .S(n5025), .Y(n5856) );
  MUX2X1 U5486 ( .B(\mem<14><1> ), .A(\mem<46><1> ), .S(n5029), .Y(n5855) );
  MUX2X1 U5487 ( .B(n5856), .A(n5855), .S(n4991), .Y(n5857) );
  MUX2X1 U5488 ( .B(n5858), .A(n5857), .S(n5001), .Y(n5859) );
  MUX2X1 U5489 ( .B(n5860), .A(n5859), .S(n5008), .Y(n5876) );
  MUX2X1 U5490 ( .B(\mem<16><1> ), .A(\mem<48><1> ), .S(n5029), .Y(n5862) );
  MUX2X1 U5491 ( .B(\mem<18><1> ), .A(\mem<50><1> ), .S(n5024), .Y(n5861) );
  MUX2X1 U5492 ( .B(n5862), .A(n5861), .S(n4989), .Y(n5866) );
  MUX2X1 U5493 ( .B(\mem<20><1> ), .A(\mem<52><1> ), .S(n5029), .Y(n5864) );
  MUX2X1 U5494 ( .B(\mem<22><1> ), .A(\mem<54><1> ), .S(n5029), .Y(n5863) );
  MUX2X1 U5495 ( .B(n5864), .A(n5863), .S(n4990), .Y(n5865) );
  MUX2X1 U5496 ( .B(n5866), .A(n5865), .S(n5001), .Y(n5874) );
  MUX2X1 U5497 ( .B(\mem<24><1> ), .A(\mem<56><1> ), .S(n5029), .Y(n5868) );
  MUX2X1 U5498 ( .B(\mem<26><1> ), .A(\mem<58><1> ), .S(n5029), .Y(n5867) );
  MUX2X1 U5499 ( .B(n5868), .A(n5867), .S(n4987), .Y(n5872) );
  MUX2X1 U5500 ( .B(\mem<28><1> ), .A(\mem<60><1> ), .S(n5029), .Y(n5870) );
  MUX2X1 U5501 ( .B(\mem<30><1> ), .A(\mem<62><1> ), .S(n5029), .Y(n5869) );
  MUX2X1 U5502 ( .B(n5870), .A(n5869), .S(n4989), .Y(n5871) );
  MUX2X1 U5503 ( .B(n5872), .A(n5871), .S(n5001), .Y(n5873) );
  MUX2X1 U5504 ( .B(n5874), .A(n5873), .S(n5008), .Y(n5875) );
  MUX2X1 U5505 ( .B(n5876), .A(n5875), .S(n5017), .Y(n5908) );
  MUX2X1 U5506 ( .B(\mem<1><1> ), .A(\mem<33><1> ), .S(n5030), .Y(n5878) );
  MUX2X1 U5507 ( .B(\mem<3><1> ), .A(\mem<35><1> ), .S(n5030), .Y(n5877) );
  MUX2X1 U5508 ( .B(n5878), .A(n5877), .S(n4990), .Y(n5882) );
  MUX2X1 U5509 ( .B(\mem<5><1> ), .A(\mem<37><1> ), .S(n5029), .Y(n5880) );
  MUX2X1 U5510 ( .B(\mem<7><1> ), .A(\mem<39><1> ), .S(n5024), .Y(n5879) );
  MUX2X1 U5511 ( .B(n5880), .A(n5879), .S(n4990), .Y(n5881) );
  MUX2X1 U5512 ( .B(n5882), .A(n5881), .S(n5001), .Y(n5890) );
  MUX2X1 U5513 ( .B(\mem<9><1> ), .A(\mem<41><1> ), .S(n5030), .Y(n5884) );
  MUX2X1 U5514 ( .B(\mem<11><1> ), .A(\mem<43><1> ), .S(n5030), .Y(n5883) );
  MUX2X1 U5515 ( .B(n5884), .A(n5883), .S(n4987), .Y(n5888) );
  MUX2X1 U5516 ( .B(\mem<13><1> ), .A(\mem<45><1> ), .S(n5024), .Y(n5886) );
  MUX2X1 U5517 ( .B(\mem<15><1> ), .A(\mem<47><1> ), .S(n5029), .Y(n5885) );
  MUX2X1 U5518 ( .B(n5886), .A(n5885), .S(n4990), .Y(n5887) );
  MUX2X1 U5519 ( .B(n5888), .A(n5887), .S(n5001), .Y(n5889) );
  MUX2X1 U5520 ( .B(n5890), .A(n5889), .S(n5008), .Y(n5906) );
  MUX2X1 U5521 ( .B(\mem<17><1> ), .A(\mem<49><1> ), .S(n5025), .Y(n5892) );
  MUX2X1 U5522 ( .B(\mem<19><1> ), .A(\mem<51><1> ), .S(n5029), .Y(n5891) );
  MUX2X1 U5523 ( .B(n5892), .A(n5891), .S(n4987), .Y(n5896) );
  MUX2X1 U5524 ( .B(\mem<21><1> ), .A(\mem<53><1> ), .S(n5026), .Y(n5894) );
  MUX2X1 U5525 ( .B(\mem<23><1> ), .A(\mem<55><1> ), .S(n5024), .Y(n5893) );
  MUX2X1 U5526 ( .B(n5894), .A(n5893), .S(n4987), .Y(n5895) );
  MUX2X1 U5527 ( .B(n5896), .A(n5895), .S(n5001), .Y(n5904) );
  MUX2X1 U5528 ( .B(\mem<25><1> ), .A(\mem<57><1> ), .S(n5025), .Y(n5898) );
  MUX2X1 U5529 ( .B(\mem<27><1> ), .A(\mem<59><1> ), .S(n5029), .Y(n5897) );
  MUX2X1 U5530 ( .B(n5898), .A(n5897), .S(n4987), .Y(n5902) );
  MUX2X1 U5531 ( .B(\mem<29><1> ), .A(\mem<61><1> ), .S(n5029), .Y(n5900) );
  MUX2X1 U5532 ( .B(\mem<31><1> ), .A(\mem<63><1> ), .S(n5027), .Y(n5899) );
  MUX2X1 U5533 ( .B(n5900), .A(n5899), .S(n4990), .Y(n5901) );
  MUX2X1 U5534 ( .B(n5902), .A(n5901), .S(n5001), .Y(n5903) );
  MUX2X1 U5535 ( .B(n5904), .A(n5903), .S(n5008), .Y(n5905) );
  MUX2X1 U5536 ( .B(n5906), .A(n5905), .S(n5017), .Y(n5907) );
  MUX2X1 U5537 ( .B(n5908), .A(n5907), .S(n55), .Y(n5909) );
  MUX2X1 U5538 ( .B(\mem<0><2> ), .A(\mem<32><2> ), .S(n5029), .Y(n5911) );
  MUX2X1 U5539 ( .B(\mem<2><2> ), .A(\mem<34><2> ), .S(n5029), .Y(n5910) );
  MUX2X1 U5540 ( .B(n5911), .A(n5910), .S(n4990), .Y(n5915) );
  MUX2X1 U5541 ( .B(\mem<4><2> ), .A(\mem<36><2> ), .S(n5029), .Y(n5913) );
  MUX2X1 U5542 ( .B(\mem<6><2> ), .A(\mem<38><2> ), .S(n5028), .Y(n5912) );
  MUX2X1 U5543 ( .B(n5913), .A(n5912), .S(n4990), .Y(n5914) );
  MUX2X1 U5544 ( .B(n5915), .A(n5914), .S(n5000), .Y(n5923) );
  MUX2X1 U5545 ( .B(\mem<8><2> ), .A(\mem<40><2> ), .S(n5028), .Y(n5917) );
  MUX2X1 U5546 ( .B(\mem<10><2> ), .A(\mem<42><2> ), .S(n5028), .Y(n5916) );
  MUX2X1 U5547 ( .B(n5917), .A(n5916), .S(n4990), .Y(n5921) );
  MUX2X1 U5548 ( .B(\mem<12><2> ), .A(\mem<44><2> ), .S(n5028), .Y(n5919) );
  MUX2X1 U5549 ( .B(\mem<14><2> ), .A(\mem<46><2> ), .S(n5028), .Y(n5918) );
  MUX2X1 U5550 ( .B(n5919), .A(n5918), .S(n4990), .Y(n5920) );
  MUX2X1 U5551 ( .B(n5921), .A(n5920), .S(n5000), .Y(n5922) );
  MUX2X1 U5552 ( .B(n5923), .A(n5922), .S(n5007), .Y(n5939) );
  MUX2X1 U5553 ( .B(\mem<16><2> ), .A(\mem<48><2> ), .S(n5028), .Y(n5925) );
  MUX2X1 U5554 ( .B(\mem<18><2> ), .A(\mem<50><2> ), .S(n5028), .Y(n5924) );
  MUX2X1 U5555 ( .B(n5925), .A(n5924), .S(n4990), .Y(n5929) );
  MUX2X1 U5556 ( .B(\mem<20><2> ), .A(\mem<52><2> ), .S(n5028), .Y(n5927) );
  MUX2X1 U5557 ( .B(\mem<22><2> ), .A(\mem<54><2> ), .S(n5028), .Y(n5926) );
  MUX2X1 U5558 ( .B(n5927), .A(n5926), .S(n4990), .Y(n5928) );
  MUX2X1 U5559 ( .B(n5929), .A(n5928), .S(n5000), .Y(n5937) );
  MUX2X1 U5560 ( .B(\mem<24><2> ), .A(\mem<56><2> ), .S(n5028), .Y(n5931) );
  MUX2X1 U5561 ( .B(\mem<26><2> ), .A(\mem<58><2> ), .S(n5028), .Y(n5930) );
  MUX2X1 U5562 ( .B(n5931), .A(n5930), .S(n4990), .Y(n5935) );
  MUX2X1 U5563 ( .B(\mem<28><2> ), .A(\mem<60><2> ), .S(n5027), .Y(n5933) );
  MUX2X1 U5564 ( .B(\mem<30><2> ), .A(\mem<62><2> ), .S(n5027), .Y(n5932) );
  MUX2X1 U5565 ( .B(n5933), .A(n5932), .S(n4990), .Y(n5934) );
  MUX2X1 U5566 ( .B(n5935), .A(n5934), .S(n5000), .Y(n5936) );
  MUX2X1 U5567 ( .B(n5937), .A(n5936), .S(n5007), .Y(n5938) );
  MUX2X1 U5568 ( .B(n5939), .A(n5938), .S(n5017), .Y(n5971) );
  MUX2X1 U5569 ( .B(\mem<1><2> ), .A(\mem<33><2> ), .S(n5027), .Y(n5941) );
  MUX2X1 U5570 ( .B(\mem<3><2> ), .A(\mem<35><2> ), .S(n5027), .Y(n5940) );
  MUX2X1 U5571 ( .B(n5941), .A(n5940), .S(n4990), .Y(n5945) );
  MUX2X1 U5572 ( .B(\mem<5><2> ), .A(\mem<37><2> ), .S(n5027), .Y(n5943) );
  MUX2X1 U5573 ( .B(\mem<7><2> ), .A(\mem<39><2> ), .S(n5027), .Y(n5942) );
  MUX2X1 U5574 ( .B(n5943), .A(n5942), .S(n4990), .Y(n5944) );
  MUX2X1 U5575 ( .B(n5945), .A(n5944), .S(n5000), .Y(n5953) );
  MUX2X1 U5576 ( .B(\mem<9><2> ), .A(\mem<41><2> ), .S(n5027), .Y(n5947) );
  MUX2X1 U5577 ( .B(\mem<11><2> ), .A(\mem<43><2> ), .S(n5028), .Y(n5946) );
  MUX2X1 U5578 ( .B(n5947), .A(n5946), .S(n4990), .Y(n5951) );
  MUX2X1 U5579 ( .B(\mem<13><2> ), .A(\mem<45><2> ), .S(n5027), .Y(n5949) );
  MUX2X1 U5580 ( .B(\mem<15><2> ), .A(\mem<47><2> ), .S(n5027), .Y(n5948) );
  MUX2X1 U5581 ( .B(n5949), .A(n5948), .S(n4990), .Y(n5950) );
  MUX2X1 U5582 ( .B(n5951), .A(n5950), .S(n5000), .Y(n5952) );
  MUX2X1 U5583 ( .B(n5953), .A(n5952), .S(n5007), .Y(n5969) );
  MUX2X1 U5584 ( .B(\mem<17><2> ), .A(\mem<49><2> ), .S(n5027), .Y(n5955) );
  MUX2X1 U5585 ( .B(\mem<19><2> ), .A(\mem<51><2> ), .S(n5027), .Y(n5954) );
  MUX2X1 U5586 ( .B(n5955), .A(n5954), .S(n4989), .Y(n5959) );
  MUX2X1 U5587 ( .B(\mem<21><2> ), .A(\mem<53><2> ), .S(n5026), .Y(n5957) );
  MUX2X1 U5588 ( .B(\mem<23><2> ), .A(\mem<55><2> ), .S(n5026), .Y(n5956) );
  MUX2X1 U5589 ( .B(n5957), .A(n5956), .S(n4989), .Y(n5958) );
  MUX2X1 U5590 ( .B(n5959), .A(n5958), .S(n5000), .Y(n5967) );
  MUX2X1 U5591 ( .B(\mem<25><2> ), .A(\mem<57><2> ), .S(n5026), .Y(n5961) );
  MUX2X1 U5592 ( .B(\mem<27><2> ), .A(\mem<59><2> ), .S(n5028), .Y(n5960) );
  MUX2X1 U5593 ( .B(n5961), .A(n5960), .S(n4989), .Y(n5965) );
  MUX2X1 U5594 ( .B(\mem<29><2> ), .A(\mem<61><2> ), .S(n5032), .Y(n5963) );
  MUX2X1 U5595 ( .B(\mem<31><2> ), .A(\mem<63><2> ), .S(n5024), .Y(n5962) );
  MUX2X1 U5596 ( .B(n5963), .A(n5962), .S(n4989), .Y(n5964) );
  MUX2X1 U5597 ( .B(n5965), .A(n5964), .S(n5000), .Y(n5966) );
  MUX2X1 U5598 ( .B(n5967), .A(n5966), .S(n5007), .Y(n5968) );
  MUX2X1 U5599 ( .B(n5969), .A(n5968), .S(n5017), .Y(n5970) );
  MUX2X1 U5600 ( .B(n5971), .A(n5970), .S(n4882), .Y(n5972) );
  MUX2X1 U5601 ( .B(\mem<0><3> ), .A(\mem<32><3> ), .S(n5032), .Y(n5974) );
  MUX2X1 U5602 ( .B(\mem<2><3> ), .A(\mem<34><3> ), .S(n5031), .Y(n5973) );
  MUX2X1 U5603 ( .B(n5974), .A(n5973), .S(n4989), .Y(n5978) );
  MUX2X1 U5604 ( .B(\mem<4><3> ), .A(\mem<36><3> ), .S(n5026), .Y(n5976) );
  MUX2X1 U5605 ( .B(\mem<6><3> ), .A(\mem<38><3> ), .S(n5031), .Y(n5975) );
  MUX2X1 U5606 ( .B(n5976), .A(n5975), .S(n4989), .Y(n5977) );
  MUX2X1 U5607 ( .B(n5978), .A(n5977), .S(n5000), .Y(n5986) );
  MUX2X1 U5608 ( .B(\mem<8><3> ), .A(\mem<40><3> ), .S(n5031), .Y(n5980) );
  MUX2X1 U5609 ( .B(\mem<10><3> ), .A(\mem<42><3> ), .S(n5032), .Y(n5979) );
  MUX2X1 U5610 ( .B(n5980), .A(n5979), .S(n4989), .Y(n5984) );
  MUX2X1 U5611 ( .B(\mem<12><3> ), .A(\mem<44><3> ), .S(n5032), .Y(n5982) );
  MUX2X1 U5612 ( .B(\mem<14><3> ), .A(\mem<46><3> ), .S(n5028), .Y(n5981) );
  MUX2X1 U5613 ( .B(n5982), .A(n5981), .S(n4989), .Y(n5983) );
  MUX2X1 U5614 ( .B(n5984), .A(n5983), .S(n5000), .Y(n5985) );
  MUX2X1 U5615 ( .B(n5986), .A(n5985), .S(n5007), .Y(n6002) );
  MUX2X1 U5616 ( .B(\mem<16><3> ), .A(\mem<48><3> ), .S(n5031), .Y(n5988) );
  MUX2X1 U5617 ( .B(\mem<18><3> ), .A(\mem<50><3> ), .S(n5026), .Y(n5987) );
  MUX2X1 U5618 ( .B(n5988), .A(n5987), .S(n4989), .Y(n5992) );
  MUX2X1 U5619 ( .B(\mem<20><3> ), .A(\mem<52><3> ), .S(n5028), .Y(n5990) );
  MUX2X1 U5620 ( .B(\mem<22><3> ), .A(\mem<54><3> ), .S(n5027), .Y(n5989) );
  MUX2X1 U5621 ( .B(n5990), .A(n5989), .S(n4989), .Y(n5991) );
  MUX2X1 U5622 ( .B(n5992), .A(n5991), .S(n5000), .Y(n6000) );
  MUX2X1 U5623 ( .B(\mem<24><3> ), .A(\mem<56><3> ), .S(n5026), .Y(n5994) );
  MUX2X1 U5624 ( .B(\mem<26><3> ), .A(\mem<58><3> ), .S(n5026), .Y(n5993) );
  MUX2X1 U5625 ( .B(n5994), .A(n5993), .S(n4989), .Y(n5998) );
  MUX2X1 U5626 ( .B(\mem<28><3> ), .A(\mem<60><3> ), .S(n5026), .Y(n5996) );
  MUX2X1 U5627 ( .B(\mem<30><3> ), .A(\mem<62><3> ), .S(n5026), .Y(n5995) );
  MUX2X1 U5628 ( .B(n5996), .A(n5995), .S(n4989), .Y(n5997) );
  MUX2X1 U5629 ( .B(n5998), .A(n5997), .S(n5000), .Y(n5999) );
  MUX2X1 U5630 ( .B(n6000), .A(n5999), .S(n5007), .Y(n6001) );
  MUX2X1 U5631 ( .B(n6002), .A(n6001), .S(n5017), .Y(n6034) );
  MUX2X1 U5632 ( .B(\mem<1><3> ), .A(\mem<33><3> ), .S(n5032), .Y(n6004) );
  MUX2X1 U5633 ( .B(\mem<3><3> ), .A(\mem<35><3> ), .S(n5032), .Y(n6003) );
  MUX2X1 U5634 ( .B(n6004), .A(n6003), .S(n4988), .Y(n6008) );
  MUX2X1 U5635 ( .B(\mem<5><3> ), .A(\mem<37><3> ), .S(n5026), .Y(n6006) );
  MUX2X1 U5636 ( .B(\mem<7><3> ), .A(\mem<39><3> ), .S(n5026), .Y(n6005) );
  MUX2X1 U5637 ( .B(n6006), .A(n6005), .S(n4988), .Y(n6007) );
  MUX2X1 U5638 ( .B(n6008), .A(n6007), .S(n4999), .Y(n6016) );
  MUX2X1 U5639 ( .B(\mem<9><3> ), .A(\mem<41><3> ), .S(n5032), .Y(n6010) );
  MUX2X1 U5640 ( .B(\mem<11><3> ), .A(\mem<43><3> ), .S(n5031), .Y(n6009) );
  MUX2X1 U5641 ( .B(n6010), .A(n6009), .S(n4988), .Y(n6014) );
  MUX2X1 U5642 ( .B(\mem<13><3> ), .A(\mem<45><3> ), .S(n5026), .Y(n6012) );
  MUX2X1 U5643 ( .B(\mem<15><3> ), .A(\mem<47><3> ), .S(n5026), .Y(n6011) );
  MUX2X1 U5644 ( .B(n6012), .A(n6011), .S(n4988), .Y(n6013) );
  MUX2X1 U5645 ( .B(n6014), .A(n6013), .S(n4999), .Y(n6015) );
  MUX2X1 U5646 ( .B(n6016), .A(n6015), .S(n5007), .Y(n6032) );
  MUX2X1 U5647 ( .B(\mem<17><3> ), .A(\mem<49><3> ), .S(n5027), .Y(n6018) );
  MUX2X1 U5648 ( .B(\mem<19><3> ), .A(\mem<51><3> ), .S(n5027), .Y(n6017) );
  MUX2X1 U5649 ( .B(n6018), .A(n6017), .S(n4988), .Y(n6022) );
  MUX2X1 U5650 ( .B(\mem<21><3> ), .A(\mem<53><3> ), .S(n5026), .Y(n6020) );
  MUX2X1 U5651 ( .B(\mem<23><3> ), .A(\mem<55><3> ), .S(n5024), .Y(n6019) );
  MUX2X1 U5652 ( .B(n6020), .A(n6019), .S(n4988), .Y(n6021) );
  MUX2X1 U5653 ( .B(n6022), .A(n6021), .S(n4999), .Y(n6030) );
  MUX2X1 U5654 ( .B(\mem<25><3> ), .A(\mem<57><3> ), .S(n5027), .Y(n6024) );
  MUX2X1 U5655 ( .B(\mem<27><3> ), .A(\mem<59><3> ), .S(n5028), .Y(n6023) );
  MUX2X1 U5656 ( .B(n6024), .A(n6023), .S(n4988), .Y(n6028) );
  MUX2X1 U5657 ( .B(\mem<29><3> ), .A(\mem<61><3> ), .S(n5025), .Y(n6026) );
  MUX2X1 U5658 ( .B(\mem<31><3> ), .A(\mem<63><3> ), .S(n5025), .Y(n6025) );
  MUX2X1 U5659 ( .B(n6026), .A(n6025), .S(n4988), .Y(n6027) );
  MUX2X1 U5660 ( .B(n6028), .A(n6027), .S(n4999), .Y(n6029) );
  MUX2X1 U5661 ( .B(n6030), .A(n6029), .S(n5007), .Y(n6031) );
  MUX2X1 U5662 ( .B(n6032), .A(n6031), .S(n5017), .Y(n6033) );
  MUX2X1 U5663 ( .B(n6034), .A(n6033), .S(n99), .Y(n6035) );
  MUX2X1 U5664 ( .B(\mem<0><4> ), .A(\mem<32><4> ), .S(n5025), .Y(n6037) );
  MUX2X1 U5665 ( .B(\mem<2><4> ), .A(\mem<34><4> ), .S(n5025), .Y(n6036) );
  MUX2X1 U5666 ( .B(n6037), .A(n6036), .S(n4988), .Y(n6041) );
  MUX2X1 U5667 ( .B(\mem<4><4> ), .A(\mem<36><4> ), .S(n5025), .Y(n6039) );
  MUX2X1 U5668 ( .B(\mem<6><4> ), .A(\mem<38><4> ), .S(n5025), .Y(n6038) );
  MUX2X1 U5669 ( .B(n6039), .A(n6038), .S(n4988), .Y(n6040) );
  MUX2X1 U5670 ( .B(n6041), .A(n6040), .S(n4999), .Y(n6049) );
  MUX2X1 U5671 ( .B(\mem<8><4> ), .A(\mem<40><4> ), .S(n5025), .Y(n6043) );
  MUX2X1 U5672 ( .B(\mem<10><4> ), .A(\mem<42><4> ), .S(n5025), .Y(n6042) );
  MUX2X1 U5673 ( .B(n6043), .A(n6042), .S(n4988), .Y(n6047) );
  MUX2X1 U5674 ( .B(\mem<12><4> ), .A(\mem<44><4> ), .S(n5025), .Y(n6045) );
  MUX2X1 U5675 ( .B(\mem<14><4> ), .A(\mem<46><4> ), .S(n5025), .Y(n6044) );
  MUX2X1 U5676 ( .B(n6045), .A(n6044), .S(n4987), .Y(n6046) );
  MUX2X1 U5677 ( .B(n6047), .A(n6046), .S(n4999), .Y(n6048) );
  MUX2X1 U5678 ( .B(n6049), .A(n6048), .S(n5007), .Y(n6065) );
  MUX2X1 U5679 ( .B(\mem<16><4> ), .A(\mem<48><4> ), .S(n5025), .Y(n6051) );
  MUX2X1 U5680 ( .B(\mem<18><4> ), .A(\mem<50><4> ), .S(n5025), .Y(n6050) );
  MUX2X1 U5681 ( .B(n6051), .A(n6050), .S(n4987), .Y(n6055) );
  MUX2X1 U5682 ( .B(\mem<20><4> ), .A(\mem<52><4> ), .S(n5027), .Y(n6053) );
  MUX2X1 U5683 ( .B(\mem<22><4> ), .A(\mem<54><4> ), .S(n5027), .Y(n6052) );
  MUX2X1 U5684 ( .B(n6053), .A(n6052), .S(n4987), .Y(n6054) );
  MUX2X1 U5685 ( .B(n6055), .A(n6054), .S(n4999), .Y(n6063) );
  MUX2X1 U5686 ( .B(\mem<24><4> ), .A(\mem<56><4> ), .S(n5027), .Y(n6057) );
  MUX2X1 U5687 ( .B(\mem<26><4> ), .A(\mem<58><4> ), .S(n5031), .Y(n6056) );
  MUX2X1 U5688 ( .B(n6057), .A(n6056), .S(n4987), .Y(n6061) );
  MUX2X1 U5689 ( .B(\mem<28><4> ), .A(\mem<60><4> ), .S(n5027), .Y(n6059) );
  MUX2X1 U5690 ( .B(\mem<30><4> ), .A(\mem<62><4> ), .S(n5027), .Y(n6058) );
  MUX2X1 U5691 ( .B(n6059), .A(n6058), .S(n4987), .Y(n6060) );
  MUX2X1 U5692 ( .B(n6061), .A(n6060), .S(n4999), .Y(n6062) );
  MUX2X1 U5693 ( .B(n6063), .A(n6062), .S(n5007), .Y(n6064) );
  MUX2X1 U5694 ( .B(n6065), .A(n6064), .S(n5017), .Y(n6097) );
  MUX2X1 U5695 ( .B(\mem<1><4> ), .A(\mem<33><4> ), .S(n5028), .Y(n6067) );
  MUX2X1 U5696 ( .B(\mem<3><4> ), .A(\mem<35><4> ), .S(n5032), .Y(n6066) );
  MUX2X1 U5697 ( .B(n6067), .A(n6066), .S(n4987), .Y(n6071) );
  MUX2X1 U5698 ( .B(\mem<5><4> ), .A(\mem<37><4> ), .S(n5027), .Y(n6069) );
  MUX2X1 U5699 ( .B(\mem<7><4> ), .A(\mem<39><4> ), .S(n5024), .Y(n6068) );
  MUX2X1 U5700 ( .B(n6069), .A(n6068), .S(n4987), .Y(n6070) );
  MUX2X1 U5701 ( .B(n6071), .A(n6070), .S(n4999), .Y(n6079) );
  MUX2X1 U5702 ( .B(\mem<9><4> ), .A(\mem<41><4> ), .S(n5028), .Y(n6073) );
  MUX2X1 U5703 ( .B(\mem<11><4> ), .A(\mem<43><4> ), .S(n5028), .Y(n6072) );
  MUX2X1 U5704 ( .B(n6073), .A(n6072), .S(n4987), .Y(n6077) );
  MUX2X1 U5705 ( .B(\mem<13><4> ), .A(\mem<45><4> ), .S(n5024), .Y(n6075) );
  MUX2X1 U5706 ( .B(\mem<15><4> ), .A(\mem<47><4> ), .S(n5024), .Y(n6074) );
  MUX2X1 U5707 ( .B(n6075), .A(n6074), .S(n4987), .Y(n6076) );
  MUX2X1 U5708 ( .B(n6077), .A(n6076), .S(n4999), .Y(n6078) );
  MUX2X1 U5709 ( .B(n6079), .A(n6078), .S(n5007), .Y(n6095) );
  MUX2X1 U5710 ( .B(\mem<17><4> ), .A(\mem<49><4> ), .S(n5024), .Y(n6081) );
  MUX2X1 U5711 ( .B(\mem<19><4> ), .A(\mem<51><4> ), .S(n5024), .Y(n6080) );
  MUX2X1 U5712 ( .B(n6081), .A(n6080), .S(n4987), .Y(n6085) );
  MUX2X1 U5713 ( .B(\mem<21><4> ), .A(\mem<53><4> ), .S(n5024), .Y(n6083) );
  MUX2X1 U5714 ( .B(\mem<23><4> ), .A(\mem<55><4> ), .S(n5024), .Y(n6082) );
  MUX2X1 U5715 ( .B(n6083), .A(n6082), .S(n4987), .Y(n6084) );
  MUX2X1 U5716 ( .B(n6085), .A(n6084), .S(n4999), .Y(n6093) );
  MUX2X1 U5717 ( .B(\mem<25><4> ), .A(\mem<57><4> ), .S(n5024), .Y(n6087) );
  MUX2X1 U5718 ( .B(\mem<27><4> ), .A(\mem<59><4> ), .S(n5024), .Y(n6086) );
  MUX2X1 U5719 ( .B(n6087), .A(n6086), .S(n4987), .Y(n6091) );
  MUX2X1 U5720 ( .B(\mem<29><4> ), .A(\mem<61><4> ), .S(n5024), .Y(n6089) );
  MUX2X1 U5721 ( .B(\mem<31><4> ), .A(\mem<63><4> ), .S(n5024), .Y(n6088) );
  MUX2X1 U5722 ( .B(n6089), .A(n6088), .S(n4986), .Y(n6090) );
  MUX2X1 U5723 ( .B(n6091), .A(n6090), .S(n4998), .Y(n6092) );
  MUX2X1 U5724 ( .B(n6093), .A(n6092), .S(n5006), .Y(n6094) );
  MUX2X1 U5725 ( .B(n6095), .A(n6094), .S(n5017), .Y(n6096) );
  MUX2X1 U5726 ( .B(n6097), .A(n6096), .S(n54), .Y(n6098) );
  MUX2X1 U5727 ( .B(\mem<0><5> ), .A(\mem<16><5> ), .S(n5018), .Y(n6100) );
  MUX2X1 U5728 ( .B(\mem<2><5> ), .A(\mem<18><5> ), .S(n5016), .Y(n6099) );
  MUX2X1 U5729 ( .B(n6100), .A(n6099), .S(n4986), .Y(n6104) );
  MUX2X1 U5730 ( .B(\mem<4><5> ), .A(\mem<20><5> ), .S(n5014), .Y(n6102) );
  MUX2X1 U5731 ( .B(\mem<6><5> ), .A(\mem<22><5> ), .S(n5016), .Y(n6101) );
  MUX2X1 U5732 ( .B(n6102), .A(n6101), .S(n4986), .Y(n6103) );
  MUX2X1 U5733 ( .B(n6104), .A(n6103), .S(n4998), .Y(n6112) );
  MUX2X1 U5734 ( .B(\mem<8><5> ), .A(\mem<24><5> ), .S(n5016), .Y(n6106) );
  MUX2X1 U5735 ( .B(\mem<10><5> ), .A(\mem<26><5> ), .S(n5015), .Y(n6105) );
  MUX2X1 U5736 ( .B(n6106), .A(n6105), .S(n4986), .Y(n6110) );
  MUX2X1 U5737 ( .B(\mem<12><5> ), .A(\mem<28><5> ), .S(n5015), .Y(n6108) );
  MUX2X1 U5738 ( .B(\mem<14><5> ), .A(\mem<30><5> ), .S(n5014), .Y(n6107) );
  MUX2X1 U5739 ( .B(n6108), .A(n6107), .S(n4986), .Y(n6109) );
  MUX2X1 U5740 ( .B(n6110), .A(n6109), .S(n4998), .Y(n6111) );
  MUX2X1 U5741 ( .B(n6112), .A(n6111), .S(n5006), .Y(n6128) );
  MUX2X1 U5742 ( .B(\mem<1><5> ), .A(\mem<17><5> ), .S(n5016), .Y(n6114) );
  MUX2X1 U5743 ( .B(\mem<3><5> ), .A(\mem<19><5> ), .S(n5015), .Y(n6113) );
  MUX2X1 U5744 ( .B(n6114), .A(n6113), .S(n4986), .Y(n6118) );
  MUX2X1 U5745 ( .B(\mem<5><5> ), .A(\mem<21><5> ), .S(n5015), .Y(n6116) );
  MUX2X1 U5746 ( .B(\mem<7><5> ), .A(\mem<23><5> ), .S(n5014), .Y(n6115) );
  MUX2X1 U5747 ( .B(n6116), .A(n6115), .S(n4986), .Y(n6117) );
  MUX2X1 U5748 ( .B(n6118), .A(n6117), .S(n4998), .Y(n6126) );
  MUX2X1 U5749 ( .B(\mem<9><5> ), .A(\mem<25><5> ), .S(n5016), .Y(n6120) );
  MUX2X1 U5750 ( .B(\mem<11><5> ), .A(\mem<27><5> ), .S(n5015), .Y(n6119) );
  MUX2X1 U5751 ( .B(n6120), .A(n6119), .S(n4986), .Y(n6124) );
  MUX2X1 U5752 ( .B(\mem<13><5> ), .A(\mem<29><5> ), .S(n5016), .Y(n6122) );
  MUX2X1 U5753 ( .B(\mem<15><5> ), .A(\mem<31><5> ), .S(n5014), .Y(n6121) );
  MUX2X1 U5754 ( .B(n6122), .A(n6121), .S(n4986), .Y(n6123) );
  MUX2X1 U5755 ( .B(n6124), .A(n6123), .S(n4998), .Y(n6125) );
  MUX2X1 U5756 ( .B(n6126), .A(n6125), .S(n5006), .Y(n6127) );
  MUX2X1 U5757 ( .B(\mem<32><5> ), .A(\mem<48><5> ), .S(n5014), .Y(n6130) );
  MUX2X1 U5758 ( .B(\mem<34><5> ), .A(\mem<50><5> ), .S(n5016), .Y(n6129) );
  MUX2X1 U5759 ( .B(n6130), .A(n6129), .S(n4986), .Y(n6134) );
  MUX2X1 U5760 ( .B(\mem<36><5> ), .A(\mem<52><5> ), .S(n5016), .Y(n6132) );
  MUX2X1 U5761 ( .B(\mem<38><5> ), .A(\mem<54><5> ), .S(n5014), .Y(n6131) );
  MUX2X1 U5762 ( .B(n6132), .A(n6131), .S(n4986), .Y(n6133) );
  MUX2X1 U5763 ( .B(n6134), .A(n6133), .S(n4998), .Y(n6142) );
  MUX2X1 U5764 ( .B(\mem<40><5> ), .A(\mem<56><5> ), .S(n5016), .Y(n6136) );
  MUX2X1 U5765 ( .B(\mem<42><5> ), .A(\mem<58><5> ), .S(n5015), .Y(n6135) );
  MUX2X1 U5766 ( .B(n6136), .A(n6135), .S(n4986), .Y(n6140) );
  MUX2X1 U5767 ( .B(\mem<44><5> ), .A(\mem<60><5> ), .S(n5015), .Y(n6138) );
  MUX2X1 U5768 ( .B(\mem<46><5> ), .A(\mem<62><5> ), .S(n5015), .Y(n6137) );
  MUX2X1 U5769 ( .B(n6138), .A(n6137), .S(n4985), .Y(n6139) );
  MUX2X1 U5770 ( .B(n6140), .A(n6139), .S(n4998), .Y(n6141) );
  MUX2X1 U5771 ( .B(n6142), .A(n6141), .S(n5006), .Y(n6158) );
  MUX2X1 U5772 ( .B(\mem<33><5> ), .A(\mem<49><5> ), .S(n5014), .Y(n6144) );
  MUX2X1 U5773 ( .B(\mem<35><5> ), .A(\mem<51><5> ), .S(n5014), .Y(n6143) );
  MUX2X1 U5774 ( .B(n6144), .A(n6143), .S(n4985), .Y(n6148) );
  MUX2X1 U5775 ( .B(\mem<37><5> ), .A(\mem<53><5> ), .S(n5014), .Y(n6146) );
  MUX2X1 U5776 ( .B(\mem<39><5> ), .A(\mem<55><5> ), .S(n5016), .Y(n6145) );
  MUX2X1 U5777 ( .B(n6146), .A(n6145), .S(n4985), .Y(n6147) );
  MUX2X1 U5778 ( .B(n6148), .A(n6147), .S(n4998), .Y(n6156) );
  MUX2X1 U5779 ( .B(\mem<41><5> ), .A(\mem<57><5> ), .S(n5015), .Y(n6150) );
  MUX2X1 U5780 ( .B(\mem<43><5> ), .A(\mem<59><5> ), .S(n5018), .Y(n6149) );
  MUX2X1 U5781 ( .B(n6150), .A(n6149), .S(n4985), .Y(n6154) );
  MUX2X1 U5782 ( .B(\mem<45><5> ), .A(\mem<61><5> ), .S(n5014), .Y(n6152) );
  MUX2X1 U5783 ( .B(\mem<47><5> ), .A(\mem<63><5> ), .S(n5016), .Y(n6151) );
  MUX2X1 U5784 ( .B(n6152), .A(n6151), .S(n4985), .Y(n6153) );
  MUX2X1 U5785 ( .B(n6154), .A(n6153), .S(n4998), .Y(n6155) );
  MUX2X1 U5786 ( .B(n6156), .A(n6155), .S(n5006), .Y(n6157) );
  MUX2X1 U5787 ( .B(n6159), .A(n801), .S(n5024), .Y(n6160) );
  MUX2X1 U5788 ( .B(\mem<0><6> ), .A(\mem<16><6> ), .S(n5016), .Y(n6162) );
  MUX2X1 U5789 ( .B(\mem<2><6> ), .A(\mem<18><6> ), .S(n5014), .Y(n6161) );
  MUX2X1 U5790 ( .B(n6162), .A(n6161), .S(n4985), .Y(n6166) );
  MUX2X1 U5791 ( .B(\mem<4><6> ), .A(\mem<20><6> ), .S(n5015), .Y(n6164) );
  MUX2X1 U5792 ( .B(\mem<6><6> ), .A(\mem<22><6> ), .S(n5014), .Y(n6163) );
  MUX2X1 U5793 ( .B(n6164), .A(n6163), .S(n4985), .Y(n6165) );
  MUX2X1 U5794 ( .B(n6166), .A(n6165), .S(n4998), .Y(n6174) );
  MUX2X1 U5795 ( .B(\mem<8><6> ), .A(\mem<24><6> ), .S(n5016), .Y(n6168) );
  MUX2X1 U5796 ( .B(\mem<10><6> ), .A(\mem<26><6> ), .S(n5016), .Y(n6167) );
  MUX2X1 U5797 ( .B(n6168), .A(n6167), .S(n4985), .Y(n6172) );
  MUX2X1 U5798 ( .B(\mem<12><6> ), .A(\mem<28><6> ), .S(n5016), .Y(n6170) );
  MUX2X1 U5799 ( .B(\mem<14><6> ), .A(\mem<30><6> ), .S(n5016), .Y(n6169) );
  MUX2X1 U5800 ( .B(n6170), .A(n6169), .S(n4985), .Y(n6171) );
  MUX2X1 U5801 ( .B(n6172), .A(n6171), .S(n4998), .Y(n6173) );
  MUX2X1 U5802 ( .B(n6174), .A(n6173), .S(n5006), .Y(n6190) );
  MUX2X1 U5803 ( .B(\mem<1><6> ), .A(\mem<17><6> ), .S(n5016), .Y(n6176) );
  MUX2X1 U5804 ( .B(\mem<3><6> ), .A(\mem<19><6> ), .S(n5016), .Y(n6175) );
  MUX2X1 U5805 ( .B(n6176), .A(n6175), .S(n4985), .Y(n6180) );
  MUX2X1 U5806 ( .B(\mem<5><6> ), .A(\mem<21><6> ), .S(n5016), .Y(n6178) );
  MUX2X1 U5807 ( .B(\mem<7><6> ), .A(\mem<23><6> ), .S(n5016), .Y(n6177) );
  MUX2X1 U5808 ( .B(n6178), .A(n6177), .S(n4985), .Y(n6179) );
  MUX2X1 U5809 ( .B(n6180), .A(n6179), .S(n4998), .Y(n6188) );
  MUX2X1 U5810 ( .B(\mem<9><6> ), .A(\mem<25><6> ), .S(n5016), .Y(n6182) );
  MUX2X1 U5811 ( .B(\mem<11><6> ), .A(\mem<27><6> ), .S(n5016), .Y(n6181) );
  MUX2X1 U5812 ( .B(n6182), .A(n6181), .S(n4985), .Y(n6186) );
  MUX2X1 U5813 ( .B(\mem<13><6> ), .A(\mem<29><6> ), .S(n5016), .Y(n6184) );
  MUX2X1 U5814 ( .B(\mem<15><6> ), .A(\mem<31><6> ), .S(n5015), .Y(n6183) );
  MUX2X1 U5815 ( .B(n6184), .A(n6183), .S(n4984), .Y(n6185) );
  MUX2X1 U5816 ( .B(n6186), .A(n6185), .S(n4997), .Y(n6187) );
  MUX2X1 U5817 ( .B(n6188), .A(n6187), .S(n5006), .Y(n6189) );
  MUX2X1 U5818 ( .B(n6190), .A(n6189), .S(n4882), .Y(n6222) );
  MUX2X1 U5819 ( .B(\mem<32><6> ), .A(\mem<48><6> ), .S(n5015), .Y(n6192) );
  MUX2X1 U5820 ( .B(\mem<34><6> ), .A(\mem<50><6> ), .S(n5015), .Y(n6191) );
  MUX2X1 U5821 ( .B(n6192), .A(n6191), .S(n4984), .Y(n6196) );
  MUX2X1 U5822 ( .B(\mem<36><6> ), .A(\mem<52><6> ), .S(n5015), .Y(n6194) );
  MUX2X1 U5823 ( .B(\mem<38><6> ), .A(\mem<54><6> ), .S(n5015), .Y(n6193) );
  MUX2X1 U5824 ( .B(n6194), .A(n6193), .S(n4984), .Y(n6195) );
  MUX2X1 U5825 ( .B(n6196), .A(n6195), .S(n4997), .Y(n6204) );
  MUX2X1 U5826 ( .B(\mem<40><6> ), .A(\mem<56><6> ), .S(n5015), .Y(n6198) );
  MUX2X1 U5827 ( .B(\mem<42><6> ), .A(\mem<58><6> ), .S(n5015), .Y(n6197) );
  MUX2X1 U5828 ( .B(n6198), .A(n6197), .S(n4984), .Y(n6202) );
  MUX2X1 U5829 ( .B(\mem<44><6> ), .A(\mem<60><6> ), .S(n5015), .Y(n6200) );
  MUX2X1 U5830 ( .B(\mem<46><6> ), .A(\mem<62><6> ), .S(n5015), .Y(n6199) );
  MUX2X1 U5831 ( .B(n6200), .A(n6199), .S(n4984), .Y(n6201) );
  MUX2X1 U5832 ( .B(n6202), .A(n6201), .S(n4997), .Y(n6203) );
  MUX2X1 U5833 ( .B(n6204), .A(n6203), .S(n5006), .Y(n6220) );
  MUX2X1 U5834 ( .B(\mem<33><6> ), .A(\mem<49><6> ), .S(n5015), .Y(n6206) );
  MUX2X1 U5835 ( .B(\mem<35><6> ), .A(\mem<51><6> ), .S(n5015), .Y(n6205) );
  MUX2X1 U5836 ( .B(n6206), .A(n6205), .S(n4984), .Y(n6210) );
  MUX2X1 U5837 ( .B(\mem<37><6> ), .A(\mem<53><6> ), .S(n5015), .Y(n6208) );
  MUX2X1 U5838 ( .B(\mem<39><6> ), .A(\mem<55><6> ), .S(n5016), .Y(n6207) );
  MUX2X1 U5839 ( .B(n6208), .A(n6207), .S(n4984), .Y(n6209) );
  MUX2X1 U5840 ( .B(n6210), .A(n6209), .S(n4997), .Y(n6218) );
  MUX2X1 U5841 ( .B(\mem<41><6> ), .A(\mem<57><6> ), .S(n5015), .Y(n6212) );
  MUX2X1 U5842 ( .B(\mem<43><6> ), .A(\mem<59><6> ), .S(n5014), .Y(n6211) );
  MUX2X1 U5843 ( .B(n6212), .A(n6211), .S(n4984), .Y(n6216) );
  MUX2X1 U5844 ( .B(\mem<45><6> ), .A(\mem<61><6> ), .S(n5015), .Y(n6214) );
  MUX2X1 U5845 ( .B(\mem<47><6> ), .A(\mem<63><6> ), .S(n5015), .Y(n6213) );
  MUX2X1 U5846 ( .B(n6214), .A(n6213), .S(n4984), .Y(n6215) );
  MUX2X1 U5847 ( .B(n6216), .A(n6215), .S(n4997), .Y(n6217) );
  MUX2X1 U5848 ( .B(n6218), .A(n6217), .S(n5006), .Y(n6219) );
  MUX2X1 U5849 ( .B(n6220), .A(n6219), .S(n65), .Y(n6221) );
  MUX2X1 U5850 ( .B(n6222), .A(n6221), .S(n5024), .Y(n6223) );
  MUX2X1 U5851 ( .B(\mem<0><7> ), .A(\mem<16><7> ), .S(n5016), .Y(n6225) );
  MUX2X1 U5852 ( .B(\mem<2><7> ), .A(\mem<18><7> ), .S(n5014), .Y(n6224) );
  MUX2X1 U5853 ( .B(n6225), .A(n6224), .S(n4984), .Y(n6229) );
  MUX2X1 U5854 ( .B(\mem<4><7> ), .A(\mem<20><7> ), .S(n5014), .Y(n6227) );
  MUX2X1 U5855 ( .B(\mem<6><7> ), .A(\mem<22><7> ), .S(n5014), .Y(n6226) );
  MUX2X1 U5856 ( .B(n6227), .A(n6226), .S(n4984), .Y(n6228) );
  MUX2X1 U5857 ( .B(n6229), .A(n6228), .S(n4997), .Y(n6237) );
  MUX2X1 U5858 ( .B(\mem<8><7> ), .A(\mem<24><7> ), .S(n5014), .Y(n6231) );
  MUX2X1 U5859 ( .B(\mem<10><7> ), .A(\mem<26><7> ), .S(n5015), .Y(n6230) );
  MUX2X1 U5860 ( .B(n6231), .A(n6230), .S(n4984), .Y(n6235) );
  MUX2X1 U5861 ( .B(\mem<12><7> ), .A(\mem<28><7> ), .S(n5016), .Y(n6233) );
  MUX2X1 U5862 ( .B(\mem<14><7> ), .A(\mem<30><7> ), .S(n5014), .Y(n6232) );
  MUX2X1 U5863 ( .B(n6233), .A(n6232), .S(n4990), .Y(n6234) );
  MUX2X1 U5864 ( .B(n6235), .A(n6234), .S(n4997), .Y(n6236) );
  MUX2X1 U5865 ( .B(n6237), .A(n6236), .S(n5006), .Y(n6253) );
  MUX2X1 U5866 ( .B(\mem<1><7> ), .A(\mem<17><7> ), .S(n5014), .Y(n6239) );
  MUX2X1 U5867 ( .B(\mem<3><7> ), .A(\mem<19><7> ), .S(n5014), .Y(n6238) );
  MUX2X1 U5868 ( .B(n6239), .A(n6238), .S(n4987), .Y(n6243) );
  MUX2X1 U5869 ( .B(\mem<5><7> ), .A(\mem<21><7> ), .S(n5014), .Y(n6241) );
  MUX2X1 U5870 ( .B(\mem<7><7> ), .A(\mem<23><7> ), .S(n5014), .Y(n6240) );
  MUX2X1 U5871 ( .B(n6241), .A(n6240), .S(n4987), .Y(n6242) );
  MUX2X1 U5872 ( .B(n6243), .A(n6242), .S(n4997), .Y(n6251) );
  MUX2X1 U5873 ( .B(\mem<9><7> ), .A(\mem<25><7> ), .S(n5014), .Y(n6245) );
  MUX2X1 U5874 ( .B(\mem<11><7> ), .A(\mem<27><7> ), .S(n5014), .Y(n6244) );
  MUX2X1 U5875 ( .B(n6245), .A(n6244), .S(n4990), .Y(n6249) );
  MUX2X1 U5876 ( .B(\mem<13><7> ), .A(\mem<29><7> ), .S(n5014), .Y(n6247) );
  MUX2X1 U5877 ( .B(\mem<15><7> ), .A(\mem<31><7> ), .S(n5014), .Y(n6246) );
  MUX2X1 U5878 ( .B(n6247), .A(n6246), .S(n4990), .Y(n6248) );
  MUX2X1 U5879 ( .B(n6249), .A(n6248), .S(n4997), .Y(n6250) );
  MUX2X1 U5880 ( .B(n6251), .A(n6250), .S(n5006), .Y(n6252) );
  MUX2X1 U5881 ( .B(n6253), .A(n6252), .S(n4881), .Y(n6285) );
  MUX2X1 U5882 ( .B(\mem<32><7> ), .A(\mem<48><7> ), .S(n5014), .Y(n6255) );
  MUX2X1 U5883 ( .B(\mem<34><7> ), .A(\mem<50><7> ), .S(n5014), .Y(n6254) );
  MUX2X1 U5884 ( .B(n6255), .A(n6254), .S(n4990), .Y(n6259) );
  MUX2X1 U5885 ( .B(\mem<36><7> ), .A(\mem<52><7> ), .S(n5014), .Y(n6257) );
  MUX2X1 U5886 ( .B(\mem<38><7> ), .A(\mem<54><7> ), .S(n5015), .Y(n6256) );
  MUX2X1 U5887 ( .B(n6257), .A(n6256), .S(n4987), .Y(n6258) );
  MUX2X1 U5888 ( .B(n6259), .A(n6258), .S(n4997), .Y(n6267) );
  MUX2X1 U5889 ( .B(\mem<40><7> ), .A(\mem<56><7> ), .S(n5016), .Y(n6261) );
  MUX2X1 U5890 ( .B(\mem<42><7> ), .A(\mem<58><7> ), .S(n5014), .Y(n6260) );
  MUX2X1 U5891 ( .B(n6261), .A(n6260), .S(n4987), .Y(n6265) );
  MUX2X1 U5892 ( .B(\mem<44><7> ), .A(\mem<60><7> ), .S(n5014), .Y(n6263) );
  MUX2X1 U5893 ( .B(\mem<46><7> ), .A(\mem<62><7> ), .S(n5016), .Y(n6262) );
  MUX2X1 U5894 ( .B(n6263), .A(n6262), .S(n4990), .Y(n6264) );
  MUX2X1 U5895 ( .B(n6265), .A(n6264), .S(n4997), .Y(n6266) );
  MUX2X1 U5896 ( .B(n6267), .A(n6266), .S(n5006), .Y(n6283) );
  MUX2X1 U5897 ( .B(\mem<33><7> ), .A(\mem<49><7> ), .S(n5015), .Y(n6269) );
  MUX2X1 U5898 ( .B(\mem<35><7> ), .A(\mem<51><7> ), .S(n5015), .Y(n6268) );
  MUX2X1 U5899 ( .B(n6269), .A(n6268), .S(n4989), .Y(n6273) );
  MUX2X1 U5900 ( .B(\mem<37><7> ), .A(\mem<53><7> ), .S(n5014), .Y(n6271) );
  MUX2X1 U5901 ( .B(\mem<39><7> ), .A(\mem<55><7> ), .S(n5016), .Y(n6270) );
  MUX2X1 U5902 ( .B(n6271), .A(n6270), .S(n4990), .Y(n6272) );
  MUX2X1 U5903 ( .B(n6273), .A(n6272), .S(n4997), .Y(n6281) );
  MUX2X1 U5904 ( .B(\mem<41><7> ), .A(\mem<57><7> ), .S(n5016), .Y(n6275) );
  MUX2X1 U5905 ( .B(\mem<43><7> ), .A(\mem<59><7> ), .S(n5015), .Y(n6274) );
  MUX2X1 U5906 ( .B(n6275), .A(n6274), .S(n4988), .Y(n6279) );
  MUX2X1 U5907 ( .B(\mem<45><7> ), .A(\mem<61><7> ), .S(n5014), .Y(n6277) );
  MUX2X1 U5908 ( .B(\mem<47><7> ), .A(\mem<63><7> ), .S(n5016), .Y(n6276) );
  MUX2X1 U5909 ( .B(n6277), .A(n6276), .S(n4988), .Y(n6278) );
  MUX2X1 U5910 ( .B(n6279), .A(n6278), .S(n4999), .Y(n6280) );
  MUX2X1 U5911 ( .B(n6281), .A(n6280), .S(n5007), .Y(n6282) );
  MUX2X1 U5912 ( .B(n6285), .A(n6284), .S(n5028), .Y(n6286) );
  INVX2 U5913 ( .A(n761), .Y(n6417) );
  OAI21X1 U5914 ( .A(n6288), .B(n60), .C(n771), .Y(n6287) );
  NAND3X1 U5915 ( .A(n183), .B(n2362), .C(n1287), .Y(n6940) );
  NAND3X1 U5916 ( .A(n185), .B(n2364), .C(n1289), .Y(n6939) );
  NAND3X1 U5917 ( .A(n1291), .B(n2366), .C(n3100), .Y(n6938) );
  NAND3X1 U5918 ( .A(n187), .B(n2368), .C(n1293), .Y(n6937) );
  NAND3X1 U5919 ( .A(n189), .B(n2370), .C(n1295), .Y(n6936) );
  NAND3X1 U5920 ( .A(n1297), .B(n2372), .C(n3102), .Y(n6935) );
  NAND3X1 U5921 ( .A(n191), .B(n2374), .C(n1299), .Y(n6934) );
  NAND3X1 U5922 ( .A(n193), .B(n2376), .C(n1301), .Y(n6933) );
  INVX2 U5923 ( .A(n1686), .Y(n6292) );
  OAI21X1 U5924 ( .A(n3565), .B(n775), .C(n4977), .Y(n6295) );
  INVX2 U5925 ( .A(n6295), .Y(n6294) );
  OAI21X1 U5926 ( .A(n3665), .B(n775), .C(n4977), .Y(n6296) );
  NAND3X1 U5927 ( .A(n195), .B(n4073), .C(n3993), .Y(n6916) );
  NAND3X1 U5928 ( .A(n197), .B(n4075), .C(n3995), .Y(n6915) );
  NAND3X1 U5929 ( .A(n199), .B(n4077), .C(n849), .Y(n6914) );
  NAND3X1 U5930 ( .A(n201), .B(n4079), .C(n3997), .Y(n6913) );
  NAND3X1 U5931 ( .A(n203), .B(n4081), .C(n3999), .Y(n6912) );
  NAND3X1 U5932 ( .A(n205), .B(n4083), .C(n851), .Y(n6911) );
  NAND3X1 U5933 ( .A(n207), .B(n4085), .C(n4001), .Y(n6910) );
  NAND3X1 U5934 ( .A(n209), .B(n4087), .C(n4003), .Y(n6909) );
  OAI21X1 U5935 ( .A(n3665), .B(n100), .C(n4977), .Y(n6299) );
  NAND3X1 U5936 ( .A(n211), .B(n855), .C(n853), .Y(n6908) );
  NAND3X1 U5937 ( .A(n213), .B(n859), .C(n857), .Y(n6907) );
  NAND3X1 U5938 ( .A(n215), .B(n863), .C(n861), .Y(n6906) );
  NAND3X1 U5939 ( .A(n217), .B(n867), .C(n865), .Y(n6905) );
  NAND3X1 U5940 ( .A(n219), .B(n871), .C(n869), .Y(n6904) );
  NAND3X1 U5941 ( .A(n221), .B(n875), .C(n873), .Y(n6903) );
  NAND3X1 U5942 ( .A(n223), .B(n4004), .C(n878), .Y(n6902) );
  NAND3X1 U5943 ( .A(n225), .B(n882), .C(n880), .Y(n6901) );
  OAI21X1 U5944 ( .A(n3864), .B(n777), .C(n4977), .Y(n6301) );
  INVX2 U5945 ( .A(n6301), .Y(n6300) );
  NAND3X1 U5946 ( .A(n4127), .B(n2394), .C(n3120), .Y(n6900) );
  NAND3X1 U5947 ( .A(n4129), .B(n2396), .C(n3122), .Y(n6899) );
  NAND3X1 U5948 ( .A(n4131), .B(n2398), .C(n3124), .Y(n6898) );
  NAND3X1 U5949 ( .A(n4133), .B(n2400), .C(n3126), .Y(n6897) );
  NAND3X1 U5950 ( .A(n4135), .B(n2402), .C(n3128), .Y(n6896) );
  NAND3X1 U5951 ( .A(n4137), .B(n2404), .C(n3130), .Y(n6895) );
  NAND3X1 U5952 ( .A(n4139), .B(n2406), .C(n3132), .Y(n6894) );
  NAND3X1 U5953 ( .A(n4141), .B(n2408), .C(n3134), .Y(n6893) );
  NAND3X1 U5954 ( .A(n884), .B(n1303), .C(n3136), .Y(n6892) );
  NAND3X1 U5955 ( .A(n886), .B(n1305), .C(n3138), .Y(n6891) );
  NAND3X1 U5956 ( .A(n1307), .B(n888), .C(n3140), .Y(n6890) );
  NAND3X1 U5957 ( .A(n1309), .B(n890), .C(n3142), .Y(n6889) );
  NAND3X1 U5958 ( .A(n1311), .B(n892), .C(n3144), .Y(n6888) );
  NAND3X1 U5959 ( .A(n1313), .B(n894), .C(n3146), .Y(n6887) );
  NAND3X1 U5960 ( .A(n1315), .B(n896), .C(n3148), .Y(n6886) );
  NAND3X1 U5961 ( .A(n1317), .B(n3729), .C(n309), .Y(n6885) );
  NAND3X1 U5962 ( .A(n898), .B(n4088), .C(n311), .Y(n6884) );
  NAND3X1 U5963 ( .A(n900), .B(n4090), .C(n313), .Y(n6883) );
  NAND3X1 U5964 ( .A(n902), .B(n4093), .C(n315), .Y(n6882) );
  NAND3X1 U5965 ( .A(n904), .B(n4095), .C(n317), .Y(n6881) );
  NAND3X1 U5966 ( .A(n227), .B(n4097), .C(n906), .Y(n6880) );
  NAND3X1 U5967 ( .A(n908), .B(n4099), .C(n319), .Y(n6879) );
  NAND3X1 U5968 ( .A(n4005), .B(n4101), .C(n321), .Y(n6878) );
  NAND3X1 U5969 ( .A(n911), .B(n4103), .C(n323), .Y(n6877) );
  NAND3X1 U5970 ( .A(n2410), .B(n1319), .C(n325), .Y(n6876) );
  NAND3X1 U5971 ( .A(n1321), .B(n2412), .C(n327), .Y(n6875) );
  NAND3X1 U5972 ( .A(n1323), .B(n2414), .C(n329), .Y(n6874) );
  NAND3X1 U5973 ( .A(n1325), .B(n2416), .C(n331), .Y(n6873) );
  NAND3X1 U5974 ( .A(n229), .B(n2418), .C(n1327), .Y(n6872) );
  NAND3X1 U5975 ( .A(n1329), .B(n2420), .C(n333), .Y(n6871) );
  NAND3X1 U5976 ( .A(n1331), .B(n2422), .C(n335), .Y(n6870) );
  NAND3X1 U5977 ( .A(n1333), .B(n2424), .C(n337), .Y(n6869) );
  OR2X2 U5978 ( .A(n6404), .B(n4909), .Y(n6306) );
  OAI21X1 U5979 ( .A(n10), .B(n3713), .C(n4977), .Y(n6307) );
  INVX2 U5980 ( .A(n6307), .Y(n6305) );
  NAND3X1 U5981 ( .A(n4143), .B(n2426), .C(n3150), .Y(n6868) );
  NAND3X1 U5982 ( .A(n4145), .B(n2428), .C(n3152), .Y(n6867) );
  NAND3X1 U5983 ( .A(n4147), .B(n2430), .C(n3154), .Y(n6866) );
  NAND3X1 U5984 ( .A(n4149), .B(n2432), .C(n3156), .Y(n6865) );
  NAND3X1 U5985 ( .A(n4151), .B(n2434), .C(n3158), .Y(n6864) );
  NAND3X1 U5986 ( .A(n4153), .B(n2436), .C(n3160), .Y(n6863) );
  NAND3X1 U5987 ( .A(n4155), .B(n2438), .C(n3162), .Y(n6862) );
  NAND3X1 U5988 ( .A(n4157), .B(n2440), .C(n3164), .Y(n6861) );
  OAI21X1 U5989 ( .A(n3573), .B(n6308), .C(n4977), .Y(n6310) );
  NAND3X1 U5990 ( .A(n4159), .B(n3731), .C(n3798), .Y(n6860) );
  NAND3X1 U5991 ( .A(n4161), .B(n3733), .C(n3800), .Y(n6859) );
  NAND3X1 U5992 ( .A(n4163), .B(n3735), .C(n913), .Y(n6858) );
  NAND3X1 U5993 ( .A(n4165), .B(n3737), .C(n3802), .Y(n6857) );
  NAND3X1 U5994 ( .A(n4167), .B(n3739), .C(n915), .Y(n6856) );
  NAND3X1 U5995 ( .A(n4169), .B(n3741), .C(n917), .Y(n6855) );
  NAND3X1 U5996 ( .A(n4171), .B(n3743), .C(n919), .Y(n6854) );
  NAND3X1 U5997 ( .A(n4173), .B(n3745), .C(n3804), .Y(n6853) );
  NAND3X1 U5998 ( .A(n1335), .B(n2442), .C(n339), .Y(n6852) );
  NAND3X1 U5999 ( .A(n1337), .B(n2444), .C(n341), .Y(n6851) );
  NAND3X1 U6000 ( .A(n1339), .B(n2446), .C(n343), .Y(n6850) );
  NAND3X1 U6001 ( .A(n1341), .B(n2448), .C(n345), .Y(n6849) );
  NAND3X1 U6002 ( .A(n231), .B(n2450), .C(n1343), .Y(n6848) );
  NAND3X1 U6003 ( .A(n1345), .B(n2452), .C(n347), .Y(n6847) );
  NAND3X1 U6004 ( .A(n1347), .B(n2454), .C(n349), .Y(n6846) );
  NAND3X1 U6005 ( .A(n1349), .B(n2456), .C(n351), .Y(n6845) );
  NAND3X1 U6006 ( .A(n1351), .B(n2458), .C(n353), .Y(n6844) );
  NAND3X1 U6007 ( .A(n1353), .B(n2460), .C(n355), .Y(n6843) );
  NAND3X1 U6008 ( .A(n1355), .B(n2462), .C(n357), .Y(n6842) );
  NAND3X1 U6009 ( .A(n1357), .B(n2464), .C(n359), .Y(n6841) );
  NAND3X1 U6010 ( .A(n233), .B(n2466), .C(n1359), .Y(n6840) );
  NAND3X1 U6011 ( .A(n1361), .B(n2468), .C(n361), .Y(n6839) );
  NAND3X1 U6012 ( .A(n1363), .B(n2470), .C(n363), .Y(n6838) );
  NAND3X1 U6013 ( .A(n1365), .B(n2472), .C(n365), .Y(n6837) );
  NAND3X1 U6014 ( .A(n4175), .B(n2474), .C(n3166), .Y(n6836) );
  NAND3X1 U6015 ( .A(n4177), .B(n2476), .C(n3168), .Y(n6835) );
  NAND3X1 U6016 ( .A(n4179), .B(n2478), .C(n3170), .Y(n6834) );
  NAND3X1 U6017 ( .A(n4181), .B(n2480), .C(n3172), .Y(n6833) );
  NAND3X1 U6018 ( .A(n4183), .B(n2482), .C(n3174), .Y(n6832) );
  NAND3X1 U6019 ( .A(n4185), .B(n2484), .C(n3176), .Y(n6831) );
  NAND3X1 U6020 ( .A(n4187), .B(n2486), .C(n3178), .Y(n6830) );
  NAND3X1 U6021 ( .A(n4189), .B(n2488), .C(n3180), .Y(n6829) );
  NAND3X1 U6022 ( .A(n3886), .B(n3884), .C(n235), .Y(n6828) );
  NAND2X1 U6023 ( .A(\mem<48><0> ), .B(n3594), .Y(n6316) );
  NAND3X1 U6024 ( .A(n6316), .B(n923), .C(n921), .Y(n6820) );
  NAND2X1 U6025 ( .A(\mem<48><1> ), .B(n3594), .Y(n6317) );
  NAND3X1 U6026 ( .A(n6317), .B(n927), .C(n925), .Y(n6819) );
  NAND2X1 U6027 ( .A(\mem<48><2> ), .B(n3594), .Y(n6318) );
  NAND3X1 U6028 ( .A(n6318), .B(n931), .C(n929), .Y(n6818) );
  NAND2X1 U6029 ( .A(\mem<48><3> ), .B(n3594), .Y(n6319) );
  NAND3X1 U6030 ( .A(n6319), .B(n935), .C(n933), .Y(n6817) );
  NAND2X1 U6031 ( .A(\mem<48><4> ), .B(n3594), .Y(n6320) );
  NAND3X1 U6032 ( .A(n6320), .B(n939), .C(n937), .Y(n6816) );
  NAND2X1 U6033 ( .A(\mem<48><5> ), .B(n3594), .Y(n6321) );
  NAND3X1 U6034 ( .A(n6321), .B(n943), .C(n941), .Y(n6815) );
  NAND2X1 U6035 ( .A(\mem<48><6> ), .B(n3594), .Y(n6322) );
  NAND3X1 U6036 ( .A(n6322), .B(n947), .C(n945), .Y(n6814) );
  NAND2X1 U6037 ( .A(\mem<48><7> ), .B(n3594), .Y(n6323) );
  NAND3X1 U6038 ( .A(n6323), .B(n951), .C(n949), .Y(n6813) );
  NAND3X1 U6039 ( .A(n2490), .B(n1367), .C(n367), .Y(n6812) );
  NAND3X1 U6040 ( .A(n1369), .B(n2492), .C(n369), .Y(n6811) );
  NAND3X1 U6041 ( .A(n1371), .B(n2494), .C(n371), .Y(n6810) );
  NAND3X1 U6042 ( .A(n1373), .B(n2496), .C(n373), .Y(n6809) );
  NAND3X1 U6043 ( .A(n237), .B(n2498), .C(n1375), .Y(n6808) );
  NAND3X1 U6044 ( .A(n1377), .B(n2500), .C(n375), .Y(n6807) );
  NAND3X1 U6045 ( .A(n1379), .B(n2502), .C(n377), .Y(n6806) );
  NAND3X1 U6046 ( .A(n1381), .B(n2504), .C(n379), .Y(n6805) );
  OR2X2 U6047 ( .A(n6404), .B(n142), .Y(n6326) );
  OAI21X1 U6048 ( .A(n6328), .B(n952), .C(n4977), .Y(n6327) );
  INVX2 U6049 ( .A(n6327), .Y(n6325) );
  NAND3X1 U6050 ( .A(n4191), .B(n2506), .C(n3182), .Y(n6804) );
  NAND3X1 U6051 ( .A(n4193), .B(n2508), .C(n3184), .Y(n6803) );
  NAND3X1 U6052 ( .A(n4195), .B(n2510), .C(n3186), .Y(n6802) );
  NAND3X1 U6053 ( .A(n4197), .B(n2512), .C(n3188), .Y(n6801) );
  NAND3X1 U6054 ( .A(n4199), .B(n2514), .C(n3190), .Y(n6800) );
  NAND3X1 U6055 ( .A(n4201), .B(n2516), .C(n3192), .Y(n6799) );
  NAND3X1 U6056 ( .A(n4203), .B(n2518), .C(n3194), .Y(n6798) );
  NAND3X1 U6057 ( .A(n4205), .B(n2520), .C(n3196), .Y(n6797) );
  NAND3X1 U6058 ( .A(n3198), .B(n2522), .C(n4207), .Y(n6796) );
  NAND3X1 U6059 ( .A(n3200), .B(n2524), .C(n4209), .Y(n6795) );
  NAND3X1 U6060 ( .A(n3202), .B(n2526), .C(n4211), .Y(n6794) );
  NAND3X1 U6061 ( .A(n4213), .B(n2528), .C(n3204), .Y(n6793) );
  NAND3X1 U6062 ( .A(n4215), .B(n2530), .C(n3206), .Y(n6792) );
  NAND3X1 U6063 ( .A(n4217), .B(n2532), .C(n3208), .Y(n6791) );
  NAND3X1 U6064 ( .A(n4219), .B(n2534), .C(n3210), .Y(n6790) );
  NAND3X1 U6065 ( .A(n3212), .B(n2536), .C(n4221), .Y(n6789) );
  NAND3X1 U6066 ( .A(n4223), .B(n2538), .C(n3214), .Y(n6788) );
  NAND3X1 U6067 ( .A(n4225), .B(n2540), .C(n3216), .Y(n6787) );
  NAND3X1 U6068 ( .A(n4227), .B(n2542), .C(n3218), .Y(n6786) );
  NAND3X1 U6069 ( .A(n4229), .B(n2544), .C(n3220), .Y(n6785) );
  NAND3X1 U6070 ( .A(n4231), .B(n2546), .C(n3222), .Y(n6784) );
  NAND3X1 U6071 ( .A(n4233), .B(n2548), .C(n3224), .Y(n6783) );
  NAND3X1 U6072 ( .A(n4235), .B(n2550), .C(n3226), .Y(n6782) );
  NAND3X1 U6073 ( .A(n4237), .B(n2552), .C(n3228), .Y(n6781) );
  NAND3X1 U6074 ( .A(n4239), .B(n2554), .C(n3230), .Y(n6780) );
  NAND3X1 U6075 ( .A(n4241), .B(n2556), .C(n3232), .Y(n6779) );
  NAND3X1 U6076 ( .A(n4243), .B(n2558), .C(n3234), .Y(n6778) );
  NAND3X1 U6077 ( .A(n4245), .B(n2560), .C(n3236), .Y(n6777) );
  NAND3X1 U6078 ( .A(n4247), .B(n2562), .C(n3238), .Y(n6776) );
  NAND3X1 U6079 ( .A(n4249), .B(n2564), .C(n3240), .Y(n6775) );
  NAND3X1 U6080 ( .A(n4251), .B(n2566), .C(n3242), .Y(n6774) );
  NAND3X1 U6081 ( .A(n4253), .B(n2568), .C(n3244), .Y(n6773) );
  NAND3X1 U6082 ( .A(n4255), .B(n2570), .C(n3246), .Y(n6772) );
  NAND3X1 U6083 ( .A(n4257), .B(n2572), .C(n3248), .Y(n6771) );
  NAND3X1 U6084 ( .A(n4259), .B(n2574), .C(n3250), .Y(n6770) );
  NAND3X1 U6085 ( .A(n4261), .B(n2576), .C(n3252), .Y(n6769) );
  NAND3X1 U6086 ( .A(n4263), .B(n2578), .C(n3254), .Y(n6768) );
  NAND3X1 U6087 ( .A(n4265), .B(n2580), .C(n3256), .Y(n6767) );
  NAND3X1 U6088 ( .A(n4267), .B(n2582), .C(n3258), .Y(n6766) );
  NAND3X1 U6089 ( .A(n4269), .B(n2584), .C(n3260), .Y(n6765) );
  NAND3X1 U6090 ( .A(n1383), .B(n2586), .C(n381), .Y(n6764) );
  NAND3X1 U6091 ( .A(n1385), .B(n2588), .C(n383), .Y(n6763) );
  NAND3X1 U6092 ( .A(n1387), .B(n2590), .C(n385), .Y(n6762) );
  NAND3X1 U6093 ( .A(n1389), .B(n2592), .C(n387), .Y(n6761) );
  NAND3X1 U6094 ( .A(n239), .B(n2594), .C(n1391), .Y(n6760) );
  NAND3X1 U6095 ( .A(n1393), .B(n2596), .C(n389), .Y(n6759) );
  NAND3X1 U6096 ( .A(n1395), .B(n2598), .C(n391), .Y(n6758) );
  NAND3X1 U6097 ( .A(n1397), .B(n2600), .C(n393), .Y(n6757) );
  NAND3X1 U6098 ( .A(n2602), .B(n1399), .C(n4271), .Y(n6756) );
  NAND3X1 U6099 ( .A(n1401), .B(n2604), .C(n4273), .Y(n6755) );
  NAND3X1 U6100 ( .A(n1403), .B(n2606), .C(n4275), .Y(n6754) );
  NAND3X1 U6101 ( .A(n1405), .B(n2608), .C(n4277), .Y(n6753) );
  NAND3X1 U6102 ( .A(n1407), .B(n2610), .C(n4279), .Y(n6752) );
  NAND3X1 U6103 ( .A(n1409), .B(n2612), .C(n4281), .Y(n6751) );
  NAND3X1 U6104 ( .A(n1411), .B(n2614), .C(n4283), .Y(n6750) );
  NAND3X1 U6105 ( .A(n1413), .B(n2616), .C(n4285), .Y(n6749) );
  NAND3X1 U6106 ( .A(n4287), .B(n2618), .C(n3262), .Y(n6748) );
  NAND3X1 U6107 ( .A(n4289), .B(n2620), .C(n3264), .Y(n6747) );
  NAND3X1 U6108 ( .A(n4291), .B(n2622), .C(n3266), .Y(n6746) );
  NAND3X1 U6109 ( .A(n4293), .B(n2624), .C(n3268), .Y(n6745) );
  NAND3X1 U6110 ( .A(n4295), .B(n2626), .C(n3270), .Y(n6744) );
  NAND3X1 U6111 ( .A(n4297), .B(n2628), .C(n3272), .Y(n6743) );
  NAND3X1 U6112 ( .A(n4299), .B(n2630), .C(n3274), .Y(n6742) );
  NAND3X1 U6113 ( .A(n4301), .B(n2632), .C(n3276), .Y(n6741) );
  OR2X2 U6114 ( .A(n6404), .B(n125), .Y(n6337) );
  OAI21X1 U6115 ( .A(n9), .B(n954), .C(n4976), .Y(n6338) );
  INVX2 U6116 ( .A(n6338), .Y(n6336) );
  NAND3X1 U6117 ( .A(n4303), .B(n2634), .C(n3278), .Y(n6740) );
  NAND3X1 U6118 ( .A(n4305), .B(n2636), .C(n3280), .Y(n6739) );
  NAND3X1 U6119 ( .A(n4307), .B(n2638), .C(n3282), .Y(n6738) );
  NAND3X1 U6120 ( .A(n4309), .B(n2640), .C(n3284), .Y(n6737) );
  NAND3X1 U6121 ( .A(n4311), .B(n2642), .C(n3286), .Y(n6736) );
  NAND3X1 U6122 ( .A(n4313), .B(n2644), .C(n3288), .Y(n6735) );
  NAND3X1 U6123 ( .A(n4315), .B(n2646), .C(n3290), .Y(n6734) );
  NAND3X1 U6124 ( .A(n4317), .B(n2648), .C(n3292), .Y(n6733) );
  OAI21X1 U6125 ( .A(n6339), .B(n955), .C(n4976), .Y(n6341) );
  NAND3X1 U6126 ( .A(n4319), .B(n2650), .C(n3294), .Y(n6732) );
  NAND3X1 U6127 ( .A(n4321), .B(n2652), .C(n3296), .Y(n6731) );
  NAND3X1 U6128 ( .A(n4323), .B(n2654), .C(n3298), .Y(n6730) );
  NAND3X1 U6129 ( .A(n4325), .B(n2656), .C(n3300), .Y(n6729) );
  NAND3X1 U6130 ( .A(n4327), .B(n2658), .C(n3302), .Y(n6728) );
  NAND3X1 U6131 ( .A(n4329), .B(n2660), .C(n3304), .Y(n6727) );
  NAND3X1 U6132 ( .A(n4331), .B(n2662), .C(n3306), .Y(n6726) );
  NAND3X1 U6133 ( .A(n4333), .B(n2664), .C(n3308), .Y(n6725) );
  NAND3X1 U6134 ( .A(n1415), .B(n2666), .C(n395), .Y(n6724) );
  NAND3X1 U6135 ( .A(n1417), .B(n2668), .C(n397), .Y(n6723) );
  NAND3X1 U6136 ( .A(n1419), .B(n2670), .C(n399), .Y(n6722) );
  NAND3X1 U6137 ( .A(n401), .B(n2672), .C(n1421), .Y(n6721) );
  NAND3X1 U6138 ( .A(n241), .B(n2674), .C(n1423), .Y(n6720) );
  NAND3X1 U6139 ( .A(n1425), .B(n2676), .C(n403), .Y(n6719) );
  NAND3X1 U6140 ( .A(n405), .B(n2678), .C(n1427), .Y(n6718) );
  NAND3X1 U6141 ( .A(n1429), .B(n2680), .C(n407), .Y(n6717) );
  NAND3X1 U6142 ( .A(n1431), .B(n2682), .C(n409), .Y(n6716) );
  NAND3X1 U6143 ( .A(n1433), .B(n2684), .C(n411), .Y(n6715) );
  NAND3X1 U6144 ( .A(n1435), .B(n2686), .C(n413), .Y(n6714) );
  NAND3X1 U6145 ( .A(n1437), .B(n2688), .C(n415), .Y(n6713) );
  NAND3X1 U6146 ( .A(n2690), .B(n243), .C(n1439), .Y(n6712) );
  NAND3X1 U6147 ( .A(n1441), .B(n2692), .C(n417), .Y(n6711) );
  NAND3X1 U6148 ( .A(n1443), .B(n2694), .C(n419), .Y(n6710) );
  NAND3X1 U6149 ( .A(n1445), .B(n2696), .C(n421), .Y(n6709) );
  NAND3X1 U6150 ( .A(n4335), .B(n2698), .C(n3310), .Y(n6708) );
  NAND3X1 U6151 ( .A(n4337), .B(n2700), .C(n3312), .Y(n6707) );
  NAND3X1 U6152 ( .A(n4339), .B(n2702), .C(n3314), .Y(n6706) );
  NAND3X1 U6153 ( .A(n4341), .B(n2704), .C(n3316), .Y(n6705) );
  NAND3X1 U6154 ( .A(n4343), .B(n2706), .C(n3318), .Y(n6704) );
  NAND3X1 U6155 ( .A(n4345), .B(n2708), .C(n3320), .Y(n6703) );
  NAND3X1 U6156 ( .A(n4347), .B(n2710), .C(n3322), .Y(n6702) );
  NAND3X1 U6157 ( .A(n4349), .B(n2712), .C(n3324), .Y(n6701) );
  NAND3X1 U6158 ( .A(n1447), .B(n2714), .C(n423), .Y(n6700) );
  NAND3X1 U6159 ( .A(n1449), .B(n2716), .C(n425), .Y(n6699) );
  NAND3X1 U6160 ( .A(n1451), .B(n2718), .C(n427), .Y(n6698) );
  NAND3X1 U6161 ( .A(n1453), .B(n2720), .C(n429), .Y(n6697) );
  NAND3X1 U6162 ( .A(n245), .B(n2722), .C(n1455), .Y(n6696) );
  NAND3X1 U6163 ( .A(n1457), .B(n2724), .C(n431), .Y(n6695) );
  NAND3X1 U6164 ( .A(n1459), .B(n2726), .C(n433), .Y(n6694) );
  NAND3X1 U6165 ( .A(n1461), .B(n2728), .C(n435), .Y(n6693) );
  OAI21X1 U6166 ( .A(n804), .B(n4814), .C(n4976), .Y(n6348) );
  NAND3X1 U6167 ( .A(n3689), .B(n4351), .C(n3326), .Y(n6692) );
  NAND3X1 U6168 ( .A(n3691), .B(n4353), .C(n3328), .Y(n6691) );
  NAND3X1 U6169 ( .A(n957), .B(n4355), .C(n3330), .Y(n6690) );
  NAND3X1 U6170 ( .A(n3693), .B(n4357), .C(n3332), .Y(n6689) );
  NAND3X1 U6171 ( .A(n959), .B(n4359), .C(n3334), .Y(n6688) );
  NAND3X1 U6172 ( .A(n961), .B(n4361), .C(n3336), .Y(n6687) );
  NAND3X1 U6173 ( .A(n963), .B(n4363), .C(n3338), .Y(n6686) );
  NAND3X1 U6174 ( .A(n3695), .B(n4365), .C(n3340), .Y(n6685) );
  OAI21X1 U6175 ( .A(n783), .B(n804), .C(n4977), .Y(n6351) );
  NAND3X1 U6176 ( .A(n247), .B(n3747), .C(n1463), .Y(n6684) );
  NAND3X1 U6177 ( .A(n249), .B(n3749), .C(n1465), .Y(n6683) );
  NAND3X1 U6178 ( .A(n251), .B(n3751), .C(n1467), .Y(n6682) );
  NAND3X1 U6179 ( .A(n253), .B(n3753), .C(n1469), .Y(n6681) );
  NAND3X1 U6180 ( .A(n255), .B(n3755), .C(n1471), .Y(n6680) );
  NAND3X1 U6181 ( .A(n257), .B(n3757), .C(n1473), .Y(n6679) );
  NAND3X1 U6182 ( .A(n259), .B(n3759), .C(n1475), .Y(n6678) );
  NAND3X1 U6183 ( .A(n261), .B(n3761), .C(n1477), .Y(n6677) );
  OR2X2 U6184 ( .A(n6352), .B(n6404), .Y(n6354) );
  OAI21X1 U6185 ( .A(n6358), .B(n6353), .C(n4976), .Y(n6357) );
  INVX2 U6186 ( .A(n6355), .Y(n6356) );
  NAND3X1 U6187 ( .A(n1479), .B(n3763), .C(n437), .Y(n6668) );
  NAND3X1 U6188 ( .A(n1481), .B(n3765), .C(n439), .Y(n6667) );
  NAND3X1 U6189 ( .A(n1483), .B(n3767), .C(n441), .Y(n6666) );
  NAND3X1 U6190 ( .A(n1485), .B(n3769), .C(n443), .Y(n6665) );
  NAND3X1 U6191 ( .A(n279), .B(n3771), .C(n1487), .Y(n6664) );
  NAND3X1 U6192 ( .A(n1489), .B(n3773), .C(n445), .Y(n6663) );
  NAND3X1 U6193 ( .A(n1491), .B(n3775), .C(n447), .Y(n6662) );
  NAND3X1 U6194 ( .A(n1493), .B(n3777), .C(n449), .Y(n6661) );
  OAI21X1 U6195 ( .A(n6363), .B(n28), .C(n4976), .Y(n6362) );
  NAND3X1 U6196 ( .A(n3358), .B(n2746), .C(n4383), .Y(n6652) );
  NAND3X1 U6197 ( .A(n4385), .B(n2748), .C(n3360), .Y(n6651) );
  NAND3X1 U6198 ( .A(n4387), .B(n2750), .C(n3362), .Y(n6650) );
  NAND3X1 U6199 ( .A(n4389), .B(n2752), .C(n3364), .Y(n6649) );
  NAND3X1 U6200 ( .A(n4391), .B(n2754), .C(n3366), .Y(n6648) );
  NAND3X1 U6201 ( .A(n4393), .B(n2756), .C(n3368), .Y(n6647) );
  NAND3X1 U6202 ( .A(n4395), .B(n2758), .C(n3370), .Y(n6646) );
  NAND3X1 U6203 ( .A(n4397), .B(n2760), .C(n3372), .Y(n6645) );
  NAND3X1 U6204 ( .A(n2762), .B(n1495), .C(n451), .Y(n6644) );
  NAND3X1 U6205 ( .A(n1497), .B(n2764), .C(n453), .Y(n6643) );
  NAND3X1 U6206 ( .A(n1499), .B(n2766), .C(n455), .Y(n6642) );
  NAND3X1 U6207 ( .A(n1501), .B(n2768), .C(n457), .Y(n6641) );
  NAND3X1 U6208 ( .A(n281), .B(n2770), .C(n1503), .Y(n6640) );
  NAND3X1 U6209 ( .A(n1505), .B(n2772), .C(n459), .Y(n6639) );
  NAND3X1 U6210 ( .A(n1507), .B(n2774), .C(n461), .Y(n6638) );
  NAND3X1 U6211 ( .A(n1509), .B(n2776), .C(n463), .Y(n6637) );
  NAND3X1 U6212 ( .A(n4105), .B(n4023), .C(n3806), .Y(n6636) );
  NAND3X1 U6213 ( .A(n4025), .B(n4107), .C(n3808), .Y(n6635) );
  NAND3X1 U6214 ( .A(n4026), .B(n4109), .C(n3810), .Y(n6634) );
  NAND3X1 U6215 ( .A(n4029), .B(n4111), .C(n3812), .Y(n6633) );
  NAND3X1 U6216 ( .A(n1511), .B(n4113), .C(n4031), .Y(n6632) );
  NAND3X1 U6217 ( .A(n4033), .B(n4115), .C(n3814), .Y(n6631) );
  NAND3X1 U6218 ( .A(n4035), .B(n4117), .C(n3816), .Y(n6630) );
  NAND3X1 U6219 ( .A(n4037), .B(n4119), .C(n3818), .Y(n6629) );
  NAND3X1 U6220 ( .A(n4039), .B(n981), .C(n3820), .Y(n6628) );
  NAND3X1 U6221 ( .A(n4041), .B(n983), .C(n3822), .Y(n6627) );
  NAND3X1 U6222 ( .A(n4043), .B(n985), .C(n3824), .Y(n6626) );
  NAND3X1 U6223 ( .A(n4045), .B(n987), .C(n3826), .Y(n6625) );
  NAND3X1 U6224 ( .A(n1513), .B(n989), .C(n4047), .Y(n6624) );
  NAND3X1 U6225 ( .A(n4049), .B(n991), .C(n3828), .Y(n6623) );
  NAND3X1 U6226 ( .A(n4050), .B(n993), .C(n3830), .Y(n6622) );
  NAND3X1 U6227 ( .A(n4053), .B(n995), .C(n3832), .Y(n6621) );
  NAND3X1 U6228 ( .A(n2778), .B(n1515), .C(n465), .Y(n6620) );
  NAND3X1 U6229 ( .A(n1517), .B(n2780), .C(n467), .Y(n6619) );
  NAND3X1 U6230 ( .A(n1519), .B(n2782), .C(n469), .Y(n6618) );
  NAND3X1 U6231 ( .A(n1521), .B(n2784), .C(n471), .Y(n6617) );
  NAND3X1 U6232 ( .A(n283), .B(n2786), .C(n1523), .Y(n6616) );
  NAND3X1 U6233 ( .A(n1525), .B(n2788), .C(n473), .Y(n6615) );
  NAND3X1 U6234 ( .A(n1527), .B(n2790), .C(n475), .Y(n6614) );
  NAND3X1 U6235 ( .A(n1529), .B(n2792), .C(n477), .Y(n6613) );
  OR2X2 U6236 ( .A(n4834), .B(n4854), .Y(n6372) );
  OAI21X1 U6237 ( .A(n6374), .B(n3559), .C(n4976), .Y(n6373) );
  NAND3X1 U6238 ( .A(n38), .B(n2794), .C(n3374), .Y(n6612) );
  NAND3X1 U6239 ( .A(n4399), .B(n2796), .C(n3376), .Y(n6611) );
  NAND3X1 U6240 ( .A(n4401), .B(n2798), .C(n3378), .Y(n6610) );
  NAND3X1 U6241 ( .A(n4403), .B(n2800), .C(n3380), .Y(n6609) );
  NAND3X1 U6242 ( .A(n4405), .B(n2802), .C(n3382), .Y(n6608) );
  NAND3X1 U6243 ( .A(n4407), .B(n2804), .C(n3384), .Y(n6607) );
  NAND3X1 U6244 ( .A(n4409), .B(n2806), .C(n3386), .Y(n6606) );
  NAND3X1 U6245 ( .A(n4411), .B(n2808), .C(n3388), .Y(n6605) );
  OAI21X1 U6246 ( .A(n51), .B(n12), .C(n4976), .Y(n6376) );
  NAND3X1 U6247 ( .A(n4413), .B(n2810), .C(n3390), .Y(n6604) );
  NAND3X1 U6248 ( .A(n4415), .B(n2812), .C(n3392), .Y(n6603) );
  NAND3X1 U6249 ( .A(n4417), .B(n2814), .C(n3394), .Y(n6602) );
  NAND3X1 U6250 ( .A(n4419), .B(n2816), .C(n3396), .Y(n6601) );
  NAND3X1 U6251 ( .A(n4421), .B(n2818), .C(n3398), .Y(n6600) );
  NAND3X1 U6252 ( .A(n4423), .B(n2820), .C(n3400), .Y(n6599) );
  NAND3X1 U6253 ( .A(n4425), .B(n2822), .C(n3402), .Y(n6598) );
  NAND3X1 U6254 ( .A(n4427), .B(n2824), .C(n3404), .Y(n6597) );
  NAND3X1 U6255 ( .A(n2826), .B(n1531), .C(n479), .Y(n6596) );
  NAND3X1 U6256 ( .A(n1533), .B(n2828), .C(n481), .Y(n6595) );
  NAND3X1 U6257 ( .A(n1535), .B(n2830), .C(n483), .Y(n6594) );
  NAND3X1 U6258 ( .A(n1537), .B(n2832), .C(n485), .Y(n6593) );
  NAND3X1 U6259 ( .A(n285), .B(n2834), .C(n1539), .Y(n6592) );
  NAND3X1 U6260 ( .A(n1541), .B(n2836), .C(n487), .Y(n6591) );
  NAND3X1 U6261 ( .A(n1543), .B(n2838), .C(n489), .Y(n6590) );
  NAND3X1 U6262 ( .A(n1545), .B(n2840), .C(n491), .Y(n6589) );
  NAND2X1 U6263 ( .A(\mem<19><0> ), .B(n3628), .Y(n6379) );
  NAND3X1 U6264 ( .A(n6379), .B(n1547), .C(n2842), .Y(n6588) );
  NAND2X1 U6265 ( .A(\mem<19><1> ), .B(n3628), .Y(n6380) );
  NAND3X1 U6266 ( .A(n6380), .B(n2844), .C(n1549), .Y(n6587) );
  NAND2X1 U6267 ( .A(\mem<19><2> ), .B(n3628), .Y(n6381) );
  NAND3X1 U6268 ( .A(n6381), .B(n2846), .C(n1551), .Y(n6586) );
  NAND2X1 U6269 ( .A(\mem<19><3> ), .B(n3628), .Y(n6382) );
  NAND3X1 U6270 ( .A(n6382), .B(n2848), .C(n1553), .Y(n6585) );
  NAND2X1 U6271 ( .A(\mem<19><4> ), .B(n3628), .Y(n6383) );
  NAND3X1 U6272 ( .A(n6383), .B(n2850), .C(n1555), .Y(n6584) );
  NAND2X1 U6273 ( .A(\mem<19><5> ), .B(n3628), .Y(n6384) );
  NAND3X1 U6274 ( .A(n6384), .B(n2852), .C(n1557), .Y(n6583) );
  NAND2X1 U6275 ( .A(\mem<19><6> ), .B(n3628), .Y(n6385) );
  NAND3X1 U6276 ( .A(n6385), .B(n2854), .C(n1559), .Y(n6582) );
  NAND2X1 U6277 ( .A(\mem<19><7> ), .B(n3628), .Y(n6386) );
  NAND3X1 U6278 ( .A(n6386), .B(n2856), .C(n1561), .Y(n6581) );
  NAND3X1 U6279 ( .A(n4429), .B(n2858), .C(n3406), .Y(n6580) );
  NAND3X1 U6280 ( .A(n4431), .B(n2860), .C(n3408), .Y(n6579) );
  NAND3X1 U6281 ( .A(n4433), .B(n2862), .C(n3410), .Y(n6578) );
  NAND3X1 U6282 ( .A(n4435), .B(n2864), .C(n3412), .Y(n6577) );
  NAND3X1 U6283 ( .A(n4437), .B(n2866), .C(n3414), .Y(n6576) );
  NAND3X1 U6284 ( .A(n4439), .B(n2868), .C(n3416), .Y(n6575) );
  NAND3X1 U6285 ( .A(n4441), .B(n2870), .C(n3418), .Y(n6574) );
  NAND3X1 U6286 ( .A(n4443), .B(n2872), .C(n3420), .Y(n6573) );
  NAND3X1 U6287 ( .A(n3834), .B(n997), .C(n4445), .Y(n6572) );
  NAND3X1 U6288 ( .A(n4447), .B(n999), .C(n3836), .Y(n6571) );
  NAND3X1 U6289 ( .A(n4449), .B(n1001), .C(n3838), .Y(n6570) );
  NAND3X1 U6290 ( .A(n4451), .B(n1003), .C(n3840), .Y(n6569) );
  NAND3X1 U6291 ( .A(n4453), .B(n1007), .C(n1005), .Y(n6568) );
  NAND3X1 U6292 ( .A(n4455), .B(n1010), .C(n3841), .Y(n6567) );
  NAND3X1 U6293 ( .A(n4457), .B(n1014), .C(n1012), .Y(n6566) );
  NAND3X1 U6294 ( .A(n4459), .B(n1016), .C(n3843), .Y(n6565) );
  NAND3X1 U6295 ( .A(n4461), .B(n3778), .C(n3422), .Y(n6564) );
  NAND3X1 U6296 ( .A(n4463), .B(n3779), .C(n3424), .Y(n6563) );
  NAND3X1 U6297 ( .A(n4465), .B(n1020), .C(n3426), .Y(n6562) );
  NAND3X1 U6298 ( .A(n1563), .B(n1022), .C(n4467), .Y(n6561) );
  NAND3X1 U6299 ( .A(n1565), .B(n1024), .C(n4469), .Y(n6560) );
  NAND3X1 U6300 ( .A(n1567), .B(n1026), .C(n4471), .Y(n6559) );
  NAND3X1 U6301 ( .A(n4473), .B(n1028), .C(n1569), .Y(n6558) );
  NAND3X1 U6302 ( .A(n1571), .B(n1030), .C(n4475), .Y(n6557) );
  NAND3X1 U6303 ( .A(n2874), .B(n1573), .C(n493), .Y(n6556) );
  NAND3X1 U6304 ( .A(n1575), .B(n2876), .C(n495), .Y(n6555) );
  NAND3X1 U6305 ( .A(n1577), .B(n2878), .C(n497), .Y(n6554) );
  NAND3X1 U6306 ( .A(n1579), .B(n2880), .C(n499), .Y(n6553) );
  NAND3X1 U6307 ( .A(n287), .B(n2882), .C(n1581), .Y(n6552) );
  NAND3X1 U6308 ( .A(n1583), .B(n2884), .C(n501), .Y(n6551) );
  NAND3X1 U6309 ( .A(n1585), .B(n2886), .C(n503), .Y(n6550) );
  NAND3X1 U6310 ( .A(n1587), .B(n2888), .C(n505), .Y(n6549) );
  OR2X2 U6311 ( .A(n6404), .B(n4963), .Y(n6392) );
  OAI21X1 U6312 ( .A(n6394), .B(n4659), .C(n4976), .Y(n6393) );
  INVX2 U6313 ( .A(n6393), .Y(n6391) );
  NAND3X1 U6314 ( .A(n4477), .B(n2890), .C(n3428), .Y(n6548) );
  NAND3X1 U6315 ( .A(n4479), .B(n2892), .C(n3430), .Y(n6547) );
  NAND3X1 U6316 ( .A(n4481), .B(n2894), .C(n3432), .Y(n6546) );
  NAND3X1 U6317 ( .A(n4483), .B(n2896), .C(n3434), .Y(n6545) );
  NAND3X1 U6318 ( .A(n4485), .B(n2898), .C(n3436), .Y(n6544) );
  NAND3X1 U6319 ( .A(n4487), .B(n2900), .C(n3438), .Y(n6543) );
  NAND3X1 U6320 ( .A(n4489), .B(n2902), .C(n3440), .Y(n6542) );
  NAND3X1 U6321 ( .A(n4491), .B(n2904), .C(n3442), .Y(n6541) );
  OAI21X1 U6322 ( .A(n6394), .B(n3718), .C(n4977), .Y(n6396) );
  NAND3X1 U6323 ( .A(n4493), .B(n2906), .C(n3444), .Y(n6540) );
  NAND3X1 U6324 ( .A(n4495), .B(n2908), .C(n3446), .Y(n6539) );
  NAND3X1 U6325 ( .A(n4497), .B(n2910), .C(n3448), .Y(n6538) );
  NAND3X1 U6326 ( .A(n4499), .B(n2912), .C(n3450), .Y(n6537) );
  NAND3X1 U6327 ( .A(n4501), .B(n2914), .C(n3452), .Y(n6536) );
  NAND3X1 U6328 ( .A(n4503), .B(n2916), .C(n3454), .Y(n6535) );
  NAND3X1 U6329 ( .A(n4505), .B(n2918), .C(n3456), .Y(n6534) );
  NAND3X1 U6330 ( .A(n4507), .B(n2920), .C(n3458), .Y(n6533) );
  NAND3X1 U6331 ( .A(n1589), .B(n2922), .C(n507), .Y(n6532) );
  NAND3X1 U6332 ( .A(n1591), .B(n2924), .C(n509), .Y(n6531) );
  NAND3X1 U6333 ( .A(n1593), .B(n2926), .C(n511), .Y(n6530) );
  NAND3X1 U6334 ( .A(n1595), .B(n2928), .C(n513), .Y(n6529) );
  NAND3X1 U6335 ( .A(n289), .B(n2930), .C(n1597), .Y(n6528) );
  NAND3X1 U6336 ( .A(n1599), .B(n2932), .C(n515), .Y(n6527) );
  NAND3X1 U6337 ( .A(n1601), .B(n2934), .C(n517), .Y(n6526) );
  NAND3X1 U6338 ( .A(n1603), .B(n2936), .C(n519), .Y(n6525) );
  NAND3X1 U6339 ( .A(n291), .B(n2938), .C(n1605), .Y(n6524) );
  NAND3X1 U6340 ( .A(n293), .B(n2940), .C(n1607), .Y(n6523) );
  NAND3X1 U6341 ( .A(n295), .B(n2942), .C(n1609), .Y(n6522) );
  NAND3X1 U6342 ( .A(n297), .B(n2944), .C(n1611), .Y(n6521) );
  NAND3X1 U6343 ( .A(n299), .B(n2946), .C(n1613), .Y(n6520) );
  NAND3X1 U6344 ( .A(n1615), .B(n2948), .C(n521), .Y(n6519) );
  NAND3X1 U6345 ( .A(n1617), .B(n2950), .C(n523), .Y(n6518) );
  NAND3X1 U6346 ( .A(n1619), .B(n2952), .C(n525), .Y(n6517) );
  NAND3X1 U6347 ( .A(n4509), .B(n2954), .C(n3460), .Y(n6516) );
  NAND3X1 U6348 ( .A(n4511), .B(n2956), .C(n3462), .Y(n6515) );
  NAND3X1 U6349 ( .A(n4513), .B(n2958), .C(n3464), .Y(n6514) );
  NAND3X1 U6350 ( .A(n4515), .B(n2960), .C(n3466), .Y(n6513) );
  NAND3X1 U6351 ( .A(n4517), .B(n2962), .C(n3468), .Y(n6512) );
  NAND3X1 U6352 ( .A(n4519), .B(n2964), .C(n3470), .Y(n6511) );
  NAND3X1 U6353 ( .A(n4521), .B(n2966), .C(n3472), .Y(n6510) );
  NAND3X1 U6354 ( .A(n4523), .B(n2968), .C(n3474), .Y(n6509) );
  NAND3X1 U6355 ( .A(n4525), .B(n2970), .C(n3476), .Y(n6508) );
  NAND3X1 U6356 ( .A(n4527), .B(n2972), .C(n3478), .Y(n6507) );
  NAND3X1 U6357 ( .A(n4529), .B(n2974), .C(n3480), .Y(n6506) );
  NAND3X1 U6358 ( .A(n4531), .B(n2976), .C(n3482), .Y(n6505) );
  NAND3X1 U6359 ( .A(n4533), .B(n2978), .C(n3484), .Y(n6504) );
  NAND3X1 U6360 ( .A(n4535), .B(n2980), .C(n3486), .Y(n6503) );
  NAND3X1 U6361 ( .A(n4537), .B(n2982), .C(n3488), .Y(n6502) );
  NAND3X1 U6362 ( .A(n4539), .B(n2984), .C(n3490), .Y(n6501) );
  NAND3X1 U6363 ( .A(n1621), .B(n2986), .C(n4541), .Y(n6500) );
  NAND3X1 U6364 ( .A(n1623), .B(n2988), .C(n4543), .Y(n6499) );
  NAND3X1 U6365 ( .A(n1625), .B(n2990), .C(n4545), .Y(n6498) );
  NAND3X1 U6366 ( .A(n1627), .B(n2992), .C(n4547), .Y(n6497) );
  NAND3X1 U6367 ( .A(n1629), .B(n2994), .C(n4549), .Y(n6496) );
  NAND3X1 U6368 ( .A(n1631), .B(n2996), .C(n4551), .Y(n6495) );
  NAND3X1 U6369 ( .A(n1633), .B(n2998), .C(n4553), .Y(n6494) );
  NAND3X1 U6370 ( .A(n4555), .B(n1635), .C(n3492), .Y(n6493) );
  NAND3X1 U6371 ( .A(n4557), .B(n3000), .C(n3494), .Y(n6492) );
  NAND3X1 U6372 ( .A(n4559), .B(n3002), .C(n3496), .Y(n6491) );
  NAND3X1 U6373 ( .A(n4561), .B(n3004), .C(n3498), .Y(n6490) );
  NAND3X1 U6374 ( .A(n4563), .B(n3006), .C(n3500), .Y(n6489) );
  NAND3X1 U6375 ( .A(n4565), .B(n3008), .C(n3502), .Y(n6488) );
  NAND3X1 U6376 ( .A(n4567), .B(n3010), .C(n3504), .Y(n6487) );
  NAND3X1 U6377 ( .A(n4569), .B(n3506), .C(n3012), .Y(n6486) );
  NAND3X1 U6378 ( .A(n4571), .B(n3014), .C(n3508), .Y(n6485) );
  OR2X2 U6379 ( .A(n6404), .B(n4972), .Y(n6407) );
  OAI21X1 U6380 ( .A(n8), .B(n3561), .C(n4977), .Y(n6408) );
  INVX2 U6381 ( .A(n6408), .Y(n6406) );
  NAND3X1 U6382 ( .A(n4573), .B(n3016), .C(n3510), .Y(n6484) );
  NAND3X1 U6383 ( .A(n4575), .B(n3018), .C(n3512), .Y(n6483) );
  NAND3X1 U6384 ( .A(n4577), .B(n3020), .C(n3514), .Y(n6482) );
  NAND3X1 U6385 ( .A(n4579), .B(n3022), .C(n3516), .Y(n6481) );
  NAND3X1 U6386 ( .A(n4581), .B(n3024), .C(n3518), .Y(n6480) );
  NAND3X1 U6387 ( .A(n4583), .B(n3026), .C(n3520), .Y(n6479) );
  NAND3X1 U6388 ( .A(n4585), .B(n3028), .C(n3522), .Y(n6478) );
  NAND3X1 U6389 ( .A(n4587), .B(n3030), .C(n3524), .Y(n6477) );
  OAI21X1 U6390 ( .A(n6409), .B(n1031), .C(n4977), .Y(n6412) );
  NAND3X1 U6391 ( .A(n4589), .B(n3032), .C(n3526), .Y(n6476) );
  NAND3X1 U6392 ( .A(n4591), .B(n3034), .C(n3528), .Y(n6475) );
  NAND3X1 U6393 ( .A(n4593), .B(n3036), .C(n3530), .Y(n6474) );
  NAND3X1 U6394 ( .A(n4595), .B(n3038), .C(n3532), .Y(n6473) );
  NAND3X1 U6395 ( .A(n4597), .B(n3040), .C(n3534), .Y(n6472) );
  NAND3X1 U6396 ( .A(n4599), .B(n3042), .C(n3536), .Y(n6471) );
  NAND3X1 U6397 ( .A(n4601), .B(n3044), .C(n3538), .Y(n6470) );
  NAND3X1 U6398 ( .A(n4603), .B(n3046), .C(n3540), .Y(n6469) );
  NAND3X1 U6399 ( .A(n3048), .B(n1637), .C(n527), .Y(n6468) );
  NAND3X1 U6400 ( .A(n1639), .B(n3050), .C(n529), .Y(n6467) );
  NAND3X1 U6401 ( .A(n1641), .B(n3052), .C(n531), .Y(n6466) );
  NAND3X1 U6402 ( .A(n1643), .B(n3054), .C(n533), .Y(n6465) );
  NAND3X1 U6403 ( .A(n301), .B(n3056), .C(n1645), .Y(n6464) );
  NAND3X1 U6404 ( .A(n1647), .B(n3058), .C(n535), .Y(n6463) );
  NAND3X1 U6405 ( .A(n1649), .B(n3060), .C(n537), .Y(n6462) );
  NAND3X1 U6406 ( .A(n1651), .B(n3062), .C(n539), .Y(n6461) );
  NAND3X1 U6407 ( .A(n3064), .B(n1653), .C(n541), .Y(n6460) );
  NAND3X1 U6408 ( .A(n1655), .B(n3066), .C(n543), .Y(n6459) );
  NAND3X1 U6409 ( .A(n1657), .B(n3068), .C(n545), .Y(n6458) );
  NAND3X1 U6410 ( .A(n1659), .B(n3070), .C(n547), .Y(n6457) );
  NAND3X1 U6411 ( .A(n303), .B(n3072), .C(n1661), .Y(n6456) );
  NAND3X1 U6412 ( .A(n1663), .B(n3074), .C(n549), .Y(n6455) );
  NAND3X1 U6413 ( .A(n1665), .B(n3076), .C(n551), .Y(n6454) );
  NAND3X1 U6414 ( .A(n1667), .B(n3078), .C(n553), .Y(n6453) );
  NAND3X1 U6415 ( .A(n4605), .B(n3080), .C(n3542), .Y(n6452) );
  NAND3X1 U6416 ( .A(n4607), .B(n3082), .C(n3544), .Y(n6451) );
  NAND3X1 U6417 ( .A(n4609), .B(n3084), .C(n3546), .Y(n6450) );
  NAND3X1 U6418 ( .A(n4611), .B(n3086), .C(n3548), .Y(n6449) );
  NAND3X1 U6419 ( .A(n4613), .B(n3088), .C(n3550), .Y(n6448) );
  NAND3X1 U6420 ( .A(n4615), .B(n3090), .C(n3552), .Y(n6447) );
  NAND3X1 U6421 ( .A(n4617), .B(n3092), .C(n3554), .Y(n6446) );
  NAND3X1 U6422 ( .A(n4619), .B(n3094), .C(n3556), .Y(n6445) );
  OAI21X1 U6423 ( .A(n4978), .B(n78), .C(n7), .Y(n6418) );
  NAND3X1 U6424 ( .A(n3697), .B(n1033), .C(n1669), .Y(n6444) );
  NAND3X1 U6425 ( .A(n1671), .B(n1035), .C(n3699), .Y(n6443) );
  NAND3X1 U6426 ( .A(n1673), .B(n1037), .C(n3701), .Y(n6442) );
  NAND3X1 U6427 ( .A(n1675), .B(n1039), .C(n3703), .Y(n6441) );
  NAND3X1 U6428 ( .A(n1677), .B(n1041), .C(n3705), .Y(n6440) );
  NAND3X1 U6429 ( .A(n1679), .B(n1043), .C(n3707), .Y(n6439) );
  NAND3X1 U6430 ( .A(n1045), .B(n1681), .C(n3709), .Y(n6438) );
  NAND3X1 U6431 ( .A(n1683), .B(n1047), .C(n3711), .Y(n6437) );
  MUX2X1 U6432 ( .B(n6420), .A(n5076), .S(n6427), .Y(n6436) );
  MUX2X1 U6433 ( .B(n6421), .A(n5080), .S(n6427), .Y(n6435) );
  MUX2X1 U6434 ( .B(n6422), .A(n5086), .S(n6427), .Y(n6434) );
  MUX2X1 U6435 ( .B(n6423), .A(n5093), .S(n6427), .Y(n6433) );
  MUX2X1 U6436 ( .B(n6424), .A(n5097), .S(n6427), .Y(n6432) );
  MUX2X1 U6437 ( .B(n6425), .A(n5101), .S(n6427), .Y(n6431) );
  MUX2X1 U6438 ( .B(n6426), .A(n5105), .S(n6427), .Y(n6430) );
  MUX2X1 U6439 ( .B(n6428), .A(n5110), .S(n6427), .Y(n6429) );
endmodule


module fetch ( .NextPC({\NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> , 
        \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> , 
        \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> , 
        \NextPC<1> , \NextPC<0> }), clk, rst, Halt, Rti, Exception, .Instr({
        \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> , 
        \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> , 
        \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , \Instr<0> 
        }), .IncPC({\IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , 
        \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , 
        \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> , 
        \IncPC<0> }) );
  input \NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> , \NextPC<11> ,
         \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> , \NextPC<6> ,
         \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> , \NextPC<1> ,
         \NextPC<0> , clk, rst, Halt, Rti, Exception;
  output \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> ,
         \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> ,
         \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> ,
         \Instr<0> , \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> ,
         \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> ,
         \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> ,
         \IncPC<1> , \IncPC<0> ;
  wire   \actualNextPC<15> , \actualNextPC<12> , \actualNextPC<11> ,
         \actualNextPC<10> , \actualNextPC<9> , \actualNextPC<8> ,
         \actualNextPC<7> , \actualNextPC<6> , \actualNextPC<5> ,
         \actualNextPC<4> , \actualNextPC<3> , \actualNextPC<2> ,
         \actualNextPC<1> , \actualNextPC<0> , \pc<15> , \pc<14> , \pc<13> ,
         \pc<12> , \pc<11> , \pc<10> , \pc<9> , \pc<8> , \pc<7> , \pc<6> ,
         \pc<5> , \pc<4> , \pc<3> , \pc<2> , \pc<1> , \pc<0> , \nextEPC<15> ,
         \nextEPC<14> , \nextEPC<13> , \nextEPC<12> , \nextEPC<11> ,
         \nextEPC<10> , \nextEPC<9> , \nextEPC<8> , \nextEPC<7> , \nextEPC<6> ,
         \nextEPC<5> , \nextEPC<4> , \nextEPC<3> , \nextEPC<2> , \nextEPC<1> ,
         \nextEPC<0> , \epc<15> , \epc<14> , \epc<13> , \epc<12> , \epc<11> ,
         \epc<10> , \epc<9> , \epc<8> , \epc<7> , \epc<6> , \epc<5> , \epc<4> ,
         \epc<3> , \epc<2> , \epc<1> , \epc<0> , nextExcptState, curExcptState,
         n36, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;

  XOR2X1 U38 ( .A(curExcptState), .B(Exception), .Y(n36) );
  OAI21X1 U39 ( .A(n127), .B(n171), .C(n51), .Y(\nextEPC<9> ) );
  OAI21X1 U41 ( .A(n127), .B(n170), .C(n49), .Y(\nextEPC<8> ) );
  OAI21X1 U43 ( .A(n127), .B(n169), .C(n47), .Y(\nextEPC<7> ) );
  OAI21X1 U45 ( .A(n127), .B(n168), .C(n45), .Y(\nextEPC<6> ) );
  OAI21X1 U47 ( .A(n127), .B(n167), .C(n43), .Y(\nextEPC<5> ) );
  OAI21X1 U49 ( .A(n127), .B(n166), .C(n41), .Y(\nextEPC<4> ) );
  OAI21X1 U51 ( .A(n127), .B(n165), .C(n39), .Y(\nextEPC<3> ) );
  OAI21X1 U53 ( .A(n127), .B(n164), .C(n37), .Y(\nextEPC<2> ) );
  OAI21X1 U55 ( .A(n127), .B(n163), .C(n34), .Y(\nextEPC<1> ) );
  OAI21X1 U57 ( .A(n127), .B(n177), .C(n32), .Y(\nextEPC<15> ) );
  OAI21X1 U59 ( .A(n127), .B(n176), .C(n30), .Y(\nextEPC<14> ) );
  OAI21X1 U61 ( .A(n127), .B(n175), .C(n28), .Y(\nextEPC<13> ) );
  OAI21X1 U63 ( .A(n128), .B(n174), .C(n26), .Y(\nextEPC<12> ) );
  OAI21X1 U65 ( .A(n128), .B(n173), .C(n24), .Y(\nextEPC<11> ) );
  OAI21X1 U67 ( .A(n128), .B(n172), .C(n22), .Y(\nextEPC<10> ) );
  OAI21X1 U69 ( .A(n128), .B(n162), .C(n20), .Y(\nextEPC<0> ) );
  dff_144 \pc_reg[0]  ( .q(\pc<0> ), .d(\actualNextPC<0> ), .clk(clk), .rst(
        n129) );
  dff_145 \pc_reg[1]  ( .q(\pc<1> ), .d(\actualNextPC<1> ), .clk(clk), .rst(
        n129) );
  dff_146 \pc_reg[2]  ( .q(\pc<2> ), .d(\actualNextPC<2> ), .clk(clk), .rst(
        n129) );
  dff_147 \pc_reg[3]  ( .q(\pc<3> ), .d(\actualNextPC<3> ), .clk(clk), .rst(
        n129) );
  dff_148 \pc_reg[4]  ( .q(\pc<4> ), .d(\actualNextPC<4> ), .clk(clk), .rst(
        n129) );
  dff_149 \pc_reg[5]  ( .q(\pc<5> ), .d(\actualNextPC<5> ), .clk(clk), .rst(
        n129) );
  dff_150 \pc_reg[6]  ( .q(\pc<6> ), .d(\actualNextPC<6> ), .clk(clk), .rst(
        n129) );
  dff_151 \pc_reg[7]  ( .q(\pc<7> ), .d(\actualNextPC<7> ), .clk(clk), .rst(
        n129) );
  dff_152 \pc_reg[8]  ( .q(\pc<8> ), .d(\actualNextPC<8> ), .clk(clk), .rst(
        n129) );
  dff_153 \pc_reg[9]  ( .q(\pc<9> ), .d(\actualNextPC<9> ), .clk(clk), .rst(
        n129) );
  dff_154 \pc_reg[10]  ( .q(\pc<10> ), .d(\actualNextPC<10> ), .clk(clk), 
        .rst(rst) );
  dff_155 \pc_reg[11]  ( .q(\pc<11> ), .d(\actualNextPC<11> ), .clk(clk), 
        .rst(rst) );
  dff_156 \pc_reg[12]  ( .q(\pc<12> ), .d(\actualNextPC<12> ), .clk(clk), 
        .rst(n129) );
  dff_157 \pc_reg[13]  ( .q(\pc<13> ), .d(n7), .clk(clk), .rst(rst) );
  dff_158 \pc_reg[14]  ( .q(\pc<14> ), .d(n5), .clk(clk), .rst(n129) );
  dff_159 \pc_reg[15]  ( .q(\pc<15> ), .d(\actualNextPC<15> ), .clk(clk), 
        .rst(rst) );
  dff_128 \epc_reg[0]  ( .q(\epc<0> ), .d(\nextEPC<0> ), .clk(clk), .rst(rst)
         );
  dff_129 \epc_reg[1]  ( .q(\epc<1> ), .d(\nextEPC<1> ), .clk(clk), .rst(rst)
         );
  dff_130 \epc_reg[2]  ( .q(\epc<2> ), .d(\nextEPC<2> ), .clk(clk), .rst(rst)
         );
  dff_131 \epc_reg[3]  ( .q(\epc<3> ), .d(\nextEPC<3> ), .clk(clk), .rst(rst)
         );
  dff_132 \epc_reg[4]  ( .q(\epc<4> ), .d(\nextEPC<4> ), .clk(clk), .rst(rst)
         );
  dff_133 \epc_reg[5]  ( .q(\epc<5> ), .d(\nextEPC<5> ), .clk(clk), .rst(rst)
         );
  dff_134 \epc_reg[6]  ( .q(\epc<6> ), .d(\nextEPC<6> ), .clk(clk), .rst(rst)
         );
  dff_135 \epc_reg[7]  ( .q(\epc<7> ), .d(\nextEPC<7> ), .clk(clk), .rst(rst)
         );
  dff_136 \epc_reg[8]  ( .q(\epc<8> ), .d(\nextEPC<8> ), .clk(clk), .rst(rst)
         );
  dff_137 \epc_reg[9]  ( .q(\epc<9> ), .d(\nextEPC<9> ), .clk(clk), .rst(rst)
         );
  dff_138 \epc_reg[10]  ( .q(\epc<10> ), .d(\nextEPC<10> ), .clk(clk), .rst(
        rst) );
  dff_139 \epc_reg[11]  ( .q(\epc<11> ), .d(\nextEPC<11> ), .clk(clk), .rst(
        rst) );
  dff_140 \epc_reg[12]  ( .q(\epc<12> ), .d(\nextEPC<12> ), .clk(clk), .rst(
        rst) );
  dff_141 \epc_reg[13]  ( .q(\epc<13> ), .d(\nextEPC<13> ), .clk(clk), .rst(
        rst) );
  dff_142 \epc_reg[14]  ( .q(\epc<14> ), .d(\nextEPC<14> ), .clk(clk), .rst(
        rst) );
  dff_143 \epc_reg[15]  ( .q(\epc<15> ), .d(\nextEPC<15> ), .clk(clk), .rst(
        rst) );
  dff_160 excpt_reg ( .q(curExcptState), .d(nextExcptState), .clk(clk), .rst(
        rst) );
  memory2c_1 instr_mem ( .data_out({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , 
        \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , 
        \Instr<1> , \Instr<0> }), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .addr({
        \pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , \pc<10> , \pc<9> , 
        \pc<8> , \pc<7> , \pc<6> , \pc<5> , \pc<4> , \pc<3> , \pc<2> , \pc<1> , 
        \pc<0> }), .enable(1'b1), .wr(1'b0), .createdump(1'b0), .clk(clk), 
        .rst(n129) );
  cla16_2 pc_inc ( .A({n122, n119, n113, n114, n124, n116, n17, n121, n112, n1, 
        n16, n118, n14, n15, n110, n18}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), 
        .Cin(1'b0), .S({\IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , 
        \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , 
        \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> , 
        \IncPC<0> }), .Cout() );
  INVX1 U3 ( .A(n125), .Y(n140) );
  INVX1 U4 ( .A(n125), .Y(n144) );
  INVX1 U5 ( .A(n130), .Y(n129) );
  INVX1 U6 ( .A(n125), .Y(n153) );
  INVX1 U7 ( .A(Rti), .Y(n161) );
  AND2X1 U8 ( .A(Rti), .B(curExcptState), .Y(n2) );
  OR2X1 U9 ( .A(n126), .B(Exception), .Y(n131) );
  INVX1 U10 ( .A(\epc<0> ), .Y(n162) );
  INVX1 U11 ( .A(\epc<1> ), .Y(n163) );
  INVX1 U12 ( .A(\epc<2> ), .Y(n164) );
  INVX1 U13 ( .A(\epc<3> ), .Y(n165) );
  INVX1 U14 ( .A(\epc<4> ), .Y(n166) );
  INVX1 U15 ( .A(\epc<5> ), .Y(n167) );
  INVX1 U16 ( .A(\epc<6> ), .Y(n168) );
  INVX1 U17 ( .A(\epc<7> ), .Y(n169) );
  INVX1 U18 ( .A(\epc<8> ), .Y(n170) );
  INVX1 U19 ( .A(\epc<9> ), .Y(n171) );
  INVX1 U20 ( .A(\epc<10> ), .Y(n172) );
  INVX1 U21 ( .A(\epc<11> ), .Y(n173) );
  INVX1 U22 ( .A(\epc<12> ), .Y(n174) );
  INVX1 U23 ( .A(\epc<15> ), .Y(n177) );
  AND2X1 U24 ( .A(n36), .B(n161), .Y(nextExcptState) );
  INVX1 U25 ( .A(n125), .Y(n151) );
  INVX1 U26 ( .A(n125), .Y(n149) );
  INVX1 U27 ( .A(n125), .Y(n147) );
  INVX1 U28 ( .A(n125), .Y(n134) );
  INVX1 U29 ( .A(n125), .Y(n142) );
  INVX1 U30 ( .A(rst), .Y(n130) );
  INVX1 U31 ( .A(\epc<14> ), .Y(n176) );
  INVX1 U32 ( .A(\epc<13> ), .Y(n175) );
  BUFX2 U33 ( .A(\pc<6> ), .Y(n1) );
  INVX1 U34 ( .A(n2), .Y(n3) );
  AND2X2 U35 ( .A(n53), .B(n8), .Y(n4) );
  INVX1 U36 ( .A(n4), .Y(n5) );
  AND2X2 U37 ( .A(n55), .B(n9), .Y(n6) );
  INVX1 U40 ( .A(n6), .Y(n7) );
  BUFX2 U42 ( .A(n137), .Y(n8) );
  BUFX2 U44 ( .A(n139), .Y(n9) );
  AND2X2 U46 ( .A(n133), .B(n132), .Y(n10) );
  INVX1 U48 ( .A(n10), .Y(n11) );
  AND2X2 U50 ( .A(n3), .B(n132), .Y(n12) );
  AND2X1 U52 ( .A(curExcptState), .B(n161), .Y(n13) );
  BUFX2 U54 ( .A(\pc<3> ), .Y(n14) );
  BUFX2 U56 ( .A(\pc<2> ), .Y(n15) );
  BUFX2 U58 ( .A(\pc<5> ), .Y(n16) );
  BUFX2 U60 ( .A(\pc<9> ), .Y(n17) );
  BUFX2 U62 ( .A(\pc<0> ), .Y(n18) );
  INVX1 U64 ( .A(n13), .Y(n128) );
  INVX1 U66 ( .A(n13), .Y(n127) );
  AND2X2 U68 ( .A(\IncPC<0> ), .B(n128), .Y(n19) );
  INVX1 U70 ( .A(n19), .Y(n20) );
  AND2X2 U71 ( .A(\IncPC<10> ), .B(n127), .Y(n21) );
  INVX1 U72 ( .A(n21), .Y(n22) );
  AND2X2 U73 ( .A(\IncPC<11> ), .B(n128), .Y(n23) );
  INVX1 U74 ( .A(n23), .Y(n24) );
  AND2X2 U75 ( .A(\IncPC<12> ), .B(n128), .Y(n25) );
  INVX1 U76 ( .A(n25), .Y(n26) );
  AND2X2 U77 ( .A(\IncPC<13> ), .B(n128), .Y(n27) );
  INVX1 U78 ( .A(n27), .Y(n28) );
  AND2X2 U79 ( .A(\IncPC<14> ), .B(n128), .Y(n29) );
  INVX1 U80 ( .A(n29), .Y(n30) );
  AND2X2 U81 ( .A(\IncPC<15> ), .B(n128), .Y(n31) );
  INVX1 U82 ( .A(n31), .Y(n32) );
  AND2X2 U83 ( .A(\IncPC<1> ), .B(n128), .Y(n33) );
  INVX1 U84 ( .A(n33), .Y(n34) );
  AND2X2 U85 ( .A(\IncPC<2> ), .B(n128), .Y(n35) );
  INVX1 U86 ( .A(n35), .Y(n37) );
  AND2X2 U87 ( .A(\IncPC<3> ), .B(n128), .Y(n38) );
  INVX1 U88 ( .A(n38), .Y(n39) );
  AND2X2 U89 ( .A(\IncPC<4> ), .B(n128), .Y(n40) );
  INVX1 U90 ( .A(n40), .Y(n41) );
  AND2X2 U91 ( .A(\IncPC<5> ), .B(n128), .Y(n42) );
  INVX1 U92 ( .A(n42), .Y(n43) );
  AND2X2 U93 ( .A(\IncPC<6> ), .B(n128), .Y(n44) );
  INVX1 U94 ( .A(n44), .Y(n45) );
  AND2X2 U95 ( .A(\IncPC<7> ), .B(n128), .Y(n46) );
  INVX1 U96 ( .A(n46), .Y(n47) );
  AND2X2 U97 ( .A(\IncPC<8> ), .B(n128), .Y(n48) );
  INVX1 U98 ( .A(n48), .Y(n49) );
  AND2X2 U99 ( .A(\IncPC<9> ), .B(n127), .Y(n50) );
  INVX1 U100 ( .A(n50), .Y(n51) );
  AND2X2 U101 ( .A(\IncPC<14> ), .B(n126), .Y(n52) );
  INVX1 U102 ( .A(n52), .Y(n53) );
  AND2X2 U103 ( .A(\IncPC<13> ), .B(n126), .Y(n54) );
  INVX1 U104 ( .A(n54), .Y(n55) );
  AND2X2 U105 ( .A(\NextPC<15> ), .B(n12), .Y(n56) );
  INVX1 U106 ( .A(n56), .Y(n57) );
  AND2X2 U107 ( .A(\NextPC<12> ), .B(n12), .Y(n58) );
  INVX1 U108 ( .A(n58), .Y(n59) );
  AND2X2 U109 ( .A(\NextPC<11> ), .B(n12), .Y(n60) );
  INVX1 U110 ( .A(n60), .Y(n61) );
  AND2X2 U111 ( .A(\NextPC<10> ), .B(n12), .Y(n62) );
  INVX1 U112 ( .A(n62), .Y(n63) );
  AND2X2 U113 ( .A(\NextPC<9> ), .B(n12), .Y(n64) );
  INVX1 U114 ( .A(n64), .Y(n65) );
  AND2X2 U115 ( .A(\NextPC<8> ), .B(n12), .Y(n66) );
  INVX1 U116 ( .A(n66), .Y(n67) );
  AND2X2 U117 ( .A(\NextPC<7> ), .B(n12), .Y(n68) );
  INVX1 U118 ( .A(n68), .Y(n69) );
  AND2X2 U119 ( .A(\NextPC<6> ), .B(n12), .Y(n70) );
  INVX1 U120 ( .A(n70), .Y(n71) );
  AND2X2 U121 ( .A(\NextPC<5> ), .B(n12), .Y(n72) );
  INVX1 U122 ( .A(n72), .Y(n73) );
  AND2X2 U123 ( .A(\NextPC<4> ), .B(n12), .Y(n74) );
  INVX1 U124 ( .A(n74), .Y(n75) );
  AND2X2 U125 ( .A(\NextPC<3> ), .B(n12), .Y(n76) );
  INVX1 U126 ( .A(n76), .Y(n77) );
  AND2X2 U127 ( .A(\NextPC<2> ), .B(n12), .Y(n78) );
  INVX1 U128 ( .A(n78), .Y(n79) );
  AND2X2 U129 ( .A(\NextPC<1> ), .B(n12), .Y(n80) );
  INVX1 U130 ( .A(n80), .Y(n81) );
  AND2X2 U131 ( .A(\NextPC<0> ), .B(n12), .Y(n82) );
  INVX1 U132 ( .A(n82), .Y(n83) );
  AND2X2 U133 ( .A(n126), .B(\IncPC<15> ), .Y(n84) );
  INVX1 U134 ( .A(n84), .Y(n85) );
  AND2X2 U135 ( .A(\IncPC<12> ), .B(n126), .Y(n86) );
  INVX1 U136 ( .A(n86), .Y(n87) );
  AND2X2 U137 ( .A(\IncPC<11> ), .B(n126), .Y(n88) );
  INVX1 U138 ( .A(n88), .Y(n89) );
  AND2X2 U139 ( .A(\IncPC<10> ), .B(n126), .Y(n90) );
  INVX1 U140 ( .A(n90), .Y(n91) );
  AND2X2 U141 ( .A(\IncPC<9> ), .B(n126), .Y(n92) );
  INVX1 U142 ( .A(n92), .Y(n93) );
  AND2X2 U143 ( .A(\IncPC<8> ), .B(n126), .Y(n94) );
  INVX1 U144 ( .A(n94), .Y(n95) );
  AND2X2 U145 ( .A(\IncPC<7> ), .B(n126), .Y(n96) );
  INVX1 U146 ( .A(n96), .Y(n97) );
  AND2X2 U147 ( .A(\IncPC<6> ), .B(n126), .Y(n98) );
  INVX1 U148 ( .A(n98), .Y(n99) );
  AND2X2 U149 ( .A(\IncPC<5> ), .B(n126), .Y(n100) );
  INVX1 U150 ( .A(n100), .Y(n101) );
  AND2X2 U151 ( .A(\IncPC<4> ), .B(n126), .Y(n102) );
  INVX1 U152 ( .A(n102), .Y(n103) );
  AND2X2 U153 ( .A(\IncPC<3> ), .B(n126), .Y(n104) );
  INVX1 U154 ( .A(n104), .Y(n105) );
  AND2X2 U155 ( .A(\IncPC<2> ), .B(n126), .Y(n106) );
  INVX1 U156 ( .A(n106), .Y(n107) );
  AND2X2 U157 ( .A(\IncPC<0> ), .B(n126), .Y(n108) );
  INVX1 U158 ( .A(n108), .Y(n109) );
  INVX1 U159 ( .A(n3), .Y(n133) );
  INVX1 U160 ( .A(n131), .Y(n132) );
  BUFX2 U161 ( .A(Halt), .Y(n126) );
  BUFX2 U162 ( .A(\pc<1> ), .Y(n110) );
  INVX1 U163 ( .A(\pc<7> ), .Y(n111) );
  INVX2 U164 ( .A(n111), .Y(n112) );
  BUFX2 U165 ( .A(\pc<13> ), .Y(n113) );
  BUFX2 U166 ( .A(\pc<12> ), .Y(n114) );
  INVX1 U167 ( .A(\pc<10> ), .Y(n115) );
  INVX2 U168 ( .A(n115), .Y(n116) );
  INVX1 U169 ( .A(\pc<4> ), .Y(n117) );
  INVX4 U170 ( .A(n117), .Y(n118) );
  BUFX2 U171 ( .A(\pc<14> ), .Y(n119) );
  INVX1 U172 ( .A(\pc<8> ), .Y(n120) );
  INVX2 U173 ( .A(n120), .Y(n121) );
  BUFX2 U174 ( .A(\pc<15> ), .Y(n122) );
  INVX1 U175 ( .A(\pc<11> ), .Y(n123) );
  INVX2 U176 ( .A(n123), .Y(n124) );
  BUFX4 U177 ( .A(n11), .Y(n125) );
  NAND2X1 U178 ( .A(\epc<15> ), .B(n134), .Y(n135) );
  NAND3X1 U179 ( .A(n135), .B(n57), .C(n85), .Y(\actualNextPC<15> ) );
  NOR2X1 U180 ( .A(n125), .B(n176), .Y(n136) );
  AOI21X1 U181 ( .A(\NextPC<14> ), .B(n12), .C(n136), .Y(n137) );
  NOR2X1 U182 ( .A(n125), .B(n175), .Y(n138) );
  AOI21X1 U183 ( .A(\NextPC<13> ), .B(n12), .C(n138), .Y(n139) );
  NAND2X1 U184 ( .A(\epc<12> ), .B(n140), .Y(n141) );
  NAND3X1 U185 ( .A(n141), .B(n59), .C(n87), .Y(\actualNextPC<12> ) );
  NAND2X1 U186 ( .A(\epc<11> ), .B(n142), .Y(n143) );
  NAND3X1 U187 ( .A(n143), .B(n61), .C(n89), .Y(\actualNextPC<11> ) );
  NAND2X1 U188 ( .A(\epc<10> ), .B(n144), .Y(n145) );
  NAND3X1 U189 ( .A(n145), .B(n63), .C(n91), .Y(\actualNextPC<10> ) );
  NAND2X1 U190 ( .A(\epc<9> ), .B(n142), .Y(n146) );
  NAND3X1 U191 ( .A(n146), .B(n65), .C(n93), .Y(\actualNextPC<9> ) );
  NAND2X1 U192 ( .A(\epc<8> ), .B(n147), .Y(n148) );
  NAND3X1 U193 ( .A(n148), .B(n67), .C(n95), .Y(\actualNextPC<8> ) );
  NAND2X1 U194 ( .A(\epc<7> ), .B(n149), .Y(n150) );
  NAND3X1 U195 ( .A(n150), .B(n69), .C(n97), .Y(\actualNextPC<7> ) );
  NAND2X1 U196 ( .A(\epc<6> ), .B(n151), .Y(n152) );
  NAND3X1 U197 ( .A(n152), .B(n71), .C(n99), .Y(\actualNextPC<6> ) );
  NAND2X1 U198 ( .A(\epc<5> ), .B(n153), .Y(n154) );
  NAND3X1 U199 ( .A(n154), .B(n73), .C(n101), .Y(\actualNextPC<5> ) );
  NAND2X1 U200 ( .A(\epc<4> ), .B(n151), .Y(n155) );
  NAND3X1 U201 ( .A(n155), .B(n75), .C(n103), .Y(\actualNextPC<4> ) );
  NAND2X1 U202 ( .A(\epc<3> ), .B(n149), .Y(n156) );
  NAND3X1 U203 ( .A(n156), .B(n77), .C(n105), .Y(\actualNextPC<3> ) );
  NAND2X1 U204 ( .A(\epc<2> ), .B(n147), .Y(n157) );
  NAND3X1 U205 ( .A(n157), .B(n79), .C(n107), .Y(\actualNextPC<2> ) );
  NAND2X1 U206 ( .A(\epc<1> ), .B(n134), .Y(n159) );
  MUX2X1 U207 ( .B(Exception), .A(\IncPC<1> ), .S(n126), .Y(n158) );
  NAND3X1 U208 ( .A(n159), .B(n81), .C(n158), .Y(\actualNextPC<1> ) );
  NAND2X1 U209 ( .A(\epc<0> ), .B(n140), .Y(n160) );
  NAND3X1 U210 ( .A(n160), .B(n83), .C(n109), .Y(\actualNextPC<0> ) );
endmodule


module decode ( clk, rst, .Instr({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , 
        \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , 
        \Instr<1> , \Instr<0> }), .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .IncPC({\IncPC<15> , \IncPC<14> , 
        \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , 
        \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , 
        \IncPC<2> , \IncPC<1> , \IncPC<0> }), .ALUOp1({\ALUOp1<15> , 
        \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , 
        \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , 
        \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), 
    .ALUOp2({\ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , 
        \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , 
        \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , 
        \ALUOp2<1> , \ALUOp2<0> }), ALUSrc, .Immediate({\Immediate<15> , 
        \Immediate<14> , \Immediate<13> , \Immediate<12> , \Immediate<11> , 
        \Immediate<10> , \Immediate<9> , \Immediate<8> , \Immediate<7> , 
        \Immediate<6> , \Immediate<5> , \Immediate<4> , \Immediate<3> , 
        \Immediate<2> , \Immediate<1> , \Immediate<0> }), Branch, Jump, 
        JumpReg, Set, Btr, InvA, InvB, Cin, .ALUOpcode({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .Func({\Func<1> , \Func<0> }), 
        MemWrite, MemRead, MemToReg, Halt, Exception, Err, Rti );
  input clk, rst, \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> ,
         \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> ,
         \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> ,
         \Instr<1> , \Instr<0> , \WriteData<15> , \WriteData<14> ,
         \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> ,
         \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> ,
         \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> ,
         \WriteData<1> , \WriteData<0> , \IncPC<15> , \IncPC<14> , \IncPC<13> ,
         \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> ,
         \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> ,
         \IncPC<2> , \IncPC<1> , \IncPC<0> ;
  output \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> ,
         \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> ,
         \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> ,
         \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , ALUSrc, \Immediate<15> , \Immediate<14> ,
         \Immediate<13> , \Immediate<12> , \Immediate<11> , \Immediate<10> ,
         \Immediate<9> , \Immediate<8> , \Immediate<7> , \Immediate<6> ,
         \Immediate<5> , \Immediate<4> , \Immediate<3> , \Immediate<2> ,
         \Immediate<1> , \Immediate<0> , Branch, Jump, JumpReg, Set, Btr, InvA,
         InvB, Cin, \ALUOpcode<2> , \ALUOpcode<1> , \ALUOpcode<0> , \Func<1> ,
         \Func<0> , MemWrite, MemRead, MemToReg, Halt, Exception, Err, Rti;
  wire   Instr_15, Instr_14, Instr_13, n182, n183, n184, \write_reg<2> ,
         \write_reg<1> , \write_reg<0> , rf_wr_en, \rs_out<15> , \rs_out<14> ,
         \rs_out<13> , \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> ,
         \rs_out<8> , \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> ,
         \rs_out<3> , \rs_out<2> , \rs_out<1> , \rs_out<0> , link, If2, If1,
         Rf, stu, N32, N33, N35, slbi, lbi, ZeroExt, N73, N74, N75, N76, N77,
         N83, N84, n60, n64, n69, n70, n71, n77, n79, n1, n2, n4, n6, n7, n8,
         n10, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n44, n45, n46, n47, n48, n49, n50, n51, n52, n54, n55, n56, n57,
         n58, n59, n61, n62, n63, n65, n66, n67, n68, n72, n73, n74, n75, n76,
         n78, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181;
  assign Instr_15 = \Instr<15> ;
  assign Instr_14 = \Instr<14> ;
  assign Instr_13 = \Instr<13> ;
  assign Err = 1'b0;

  LATCH \write_reg_reg<2>  ( .CLK(n58), .D(N35), .Q(\write_reg<2> ) );
  LATCH \write_reg_reg<1>  ( .CLK(n58), .D(N33), .Q(\write_reg<1> ) );
  LATCH \write_reg_reg<0>  ( .CLK(n58), .D(N32), .Q(\write_reg<0> ) );
  LATCH \ImmReg_reg<15>  ( .CLK(N83), .D(N84), .Q(\Immediate<15> ) );
  LATCH \ImmReg_reg<14>  ( .CLK(N83), .D(N84), .Q(\Immediate<14> ) );
  LATCH \ImmReg_reg<13>  ( .CLK(N83), .D(N84), .Q(\Immediate<13> ) );
  LATCH \ImmReg_reg<12>  ( .CLK(N83), .D(N84), .Q(\Immediate<12> ) );
  LATCH \ImmReg_reg<11>  ( .CLK(N83), .D(N84), .Q(\Immediate<11> ) );
  LATCH \ImmReg_reg<10>  ( .CLK(N83), .D(N84), .Q(\Immediate<10> ) );
  LATCH \ImmReg_reg<9>  ( .CLK(N83), .D(N77), .Q(\Immediate<9> ) );
  LATCH \ImmReg_reg<8>  ( .CLK(N83), .D(N76), .Q(\Immediate<8> ) );
  LATCH \ImmReg_reg<7>  ( .CLK(N83), .D(N75), .Q(\Immediate<7> ) );
  LATCH \ImmReg_reg<6>  ( .CLK(N83), .D(N74), .Q(\Immediate<6> ) );
  LATCH \ImmReg_reg<5>  ( .CLK(N83), .D(N73), .Q(\Immediate<5> ) );
  LATCH \ImmReg_reg<4>  ( .CLK(N83), .D(\Instr<4> ), .Q(\Immediate<4> ) );
  LATCH \ImmReg_reg<3>  ( .CLK(N83), .D(\Instr<3> ), .Q(\Immediate<3> ) );
  LATCH \ImmReg_reg<2>  ( .CLK(N83), .D(\Instr<2> ), .Q(\Immediate<2> ) );
  LATCH \ImmReg_reg<1>  ( .CLK(N83), .D(n40), .Q(\Immediate<1> ) );
  LATCH \ImmReg_reg<0>  ( .CLK(N83), .D(n39), .Q(\Immediate<0> ) );
  OAI21X1 U67 ( .A(Jump), .B(n86), .C(n172), .Y(N83) );
  OAI21X1 U68 ( .A(n61), .B(n177), .C(n171), .Y(N84) );
  OAI21X1 U69 ( .A(n61), .B(n178), .C(n171), .Y(N77) );
  OAI21X1 U70 ( .A(n61), .B(n179), .C(n171), .Y(N76) );
  OAI21X1 U71 ( .A(n94), .B(n181), .C(n56), .Y(n60) );
  OAI21X1 U72 ( .A(n172), .B(n181), .C(n56), .Y(N75) );
  OAI21X1 U73 ( .A(n172), .B(n180), .C(n56), .Y(N74) );
  OAI21X1 U74 ( .A(n172), .B(n103), .C(n56), .Y(N73) );
  NAND3X1 U77 ( .A(n94), .B(n61), .C(n82), .Y(n64) );
  NAND3X1 U82 ( .A(n74), .B(n154), .C(n80), .Y(N35) );
  AOI22X1 U83 ( .A(\Instr<10> ), .B(n70), .C(n71), .D(\Instr<4> ), .Y(n69) );
  NAND3X1 U87 ( .A(n72), .B(n154), .C(n78), .Y(N33) );
  AOI22X1 U88 ( .A(n108), .B(n70), .C(\Instr<3> ), .D(n71), .Y(n77) );
  NAND3X1 U90 ( .A(n67), .B(n154), .C(n76), .Y(N32) );
  AOI22X1 U91 ( .A(n105), .B(n70), .C(\Instr<2> ), .D(n71), .Y(n79) );
  NOR3X1 U92 ( .A(If1), .B(If2), .C(n175), .Y(n71) );
  OAI21X1 U93 ( .A(n91), .B(n176), .C(n84), .Y(n70) );
  rf regfile ( .read1data({\rs_out<15> , \rs_out<14> , \rs_out<13> , 
        \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> , \rs_out<8> , 
        \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> , \rs_out<3> , 
        \rs_out<2> , \rs_out<1> , \rs_out<0> }), .read2data({\ALUOp2<15> , 
        \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , 
        \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , 
        \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), 
        .err(), .clk(clk), .rst(rst), .read1regsel({\Instr<10> , \Instr<9> , 
        \Instr<8> }), .read2regsel({n46, n45, n118}), .writeregsel({
        \write_reg<2> , \write_reg<1> , \write_reg<0> }), .writedata({n170, 
        n169, n168, n167, n166, n165, n164, n163, n162, n161, n160, n159, n158, 
        n157, n156, n155}), .write(rf_wr_en) );
  control_unit cu ( .opcode({Instr_15, Instr_14, Instr_13, \Instr<12> , 
        \Instr<11> }), .func({n40, n39}), .aluop({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .alusrc(ALUSrc), .branch(Branch), 
        .jump(Jump), .i1(If1), .i2(If2), .r(Rf), .jumpreg(n182), .set(Set), 
        .btr(n183), .regwrite(rf_wr_en), .memwrite(MemWrite), .memread(MemRead), .memtoreg(MemToReg), .invA(InvA), .invB(InvB), .cin(Cin), .excp(Exception), 
        .zeroext(ZeroExt), .halt(n184), .slbi(slbi), .link(link), .lbi(lbi), 
        .stu(stu), .rti(Rti) );
  BUFX2 U3 ( .A(\rs_out<7> ), .Y(n1) );
  INVX1 U4 ( .A(\IncPC<1> ), .Y(n148) );
  INVX1 U5 ( .A(\IncPC<8> ), .Y(n134) );
  INVX1 U6 ( .A(\IncPC<9> ), .Y(n132) );
  INVX1 U7 ( .A(\IncPC<0> ), .Y(n150) );
  INVX1 U8 ( .A(\IncPC<7> ), .Y(n136) );
  INVX1 U9 ( .A(\IncPC<4> ), .Y(n142) );
  INVX1 U10 ( .A(\IncPC<5> ), .Y(n140) );
  INVX1 U11 ( .A(\IncPC<10> ), .Y(n130) );
  INVX1 U12 ( .A(\IncPC<14> ), .Y(n122) );
  INVX1 U13 ( .A(\IncPC<11> ), .Y(n128) );
  INVX1 U14 ( .A(\IncPC<12> ), .Y(n126) );
  INVX1 U15 ( .A(\IncPC<15> ), .Y(n120) );
  INVX1 U16 ( .A(\IncPC<6> ), .Y(n138) );
  INVX1 U17 ( .A(\IncPC<2> ), .Y(n146) );
  INVX1 U18 ( .A(\IncPC<3> ), .Y(n144) );
  INVX1 U19 ( .A(\IncPC<13> ), .Y(n124) );
  INVX1 U20 ( .A(If2), .Y(n173) );
  INVX1 U21 ( .A(ZeroExt), .Y(n174) );
  INVX1 U22 ( .A(Rf), .Y(n175) );
  INVX1 U23 ( .A(n60), .Y(n171) );
  OR2X1 U24 ( .A(n91), .B(stu), .Y(n89) );
  INVX1 U25 ( .A(stu), .Y(n176) );
  AND2X1 U26 ( .A(n90), .B(n49), .Y(n73) );
  INVX1 U27 ( .A(n117), .Y(n154) );
  INVX1 U28 ( .A(\Instr<10> ), .Y(n177) );
  AND2X1 U29 ( .A(n88), .B(n174), .Y(n93) );
  INVX4 U30 ( .A(n110), .Y(\ALUOp1<9> ) );
  AND2X2 U31 ( .A(n33), .B(n23), .Y(n2) );
  INVX1 U32 ( .A(n2), .Y(\ALUOp1<11> ) );
  AND2X2 U33 ( .A(n29), .B(n7), .Y(n4) );
  INVX1 U34 ( .A(n4), .Y(\ALUOp1<8> ) );
  AND2X2 U35 ( .A(\rs_out<8> ), .B(n52), .Y(n6) );
  INVX1 U36 ( .A(n6), .Y(n7) );
  AND2X2 U37 ( .A(n31), .B(n21), .Y(n8) );
  INVX1 U38 ( .A(n8), .Y(\ALUOp1<10> ) );
  AND2X2 U39 ( .A(n35), .B(n25), .Y(n10) );
  INVX1 U40 ( .A(n10), .Y(\ALUOp1<12> ) );
  AND2X2 U41 ( .A(n37), .B(n27), .Y(n12) );
  INVX1 U42 ( .A(n12), .Y(\ALUOp1<13> ) );
  AND2X2 U43 ( .A(\rs_out<14> ), .B(n52), .Y(n14) );
  INVX1 U44 ( .A(n14), .Y(n15) );
  AND2X2 U45 ( .A(n38), .B(\rs_out<1> ), .Y(n16) );
  INVX1 U46 ( .A(n16), .Y(n17) );
  AND2X2 U47 ( .A(\rs_out<9> ), .B(n52), .Y(n18) );
  INVX1 U48 ( .A(n18), .Y(n19) );
  AND2X2 U49 ( .A(n100), .B(n38), .Y(n20) );
  INVX1 U50 ( .A(n20), .Y(n21) );
  AND2X2 U51 ( .A(n102), .B(n38), .Y(n22) );
  INVX1 U52 ( .A(n22), .Y(n23) );
  AND2X2 U53 ( .A(\rs_out<4> ), .B(n38), .Y(n24) );
  INVX1 U54 ( .A(n24), .Y(n25) );
  AND2X2 U55 ( .A(\rs_out<5> ), .B(n38), .Y(n26) );
  INVX1 U56 ( .A(n26), .Y(n27) );
  AND2X2 U57 ( .A(n54), .B(\rs_out<0> ), .Y(n28) );
  INVX1 U58 ( .A(n28), .Y(n29) );
  AND2X2 U59 ( .A(\rs_out<10> ), .B(n52), .Y(n30) );
  INVX1 U60 ( .A(n30), .Y(n31) );
  AND2X2 U61 ( .A(\rs_out<11> ), .B(n50), .Y(n32) );
  INVX1 U62 ( .A(n32), .Y(n33) );
  AND2X2 U63 ( .A(\rs_out<12> ), .B(n50), .Y(n34) );
  INVX1 U64 ( .A(n34), .Y(n35) );
  AND2X2 U65 ( .A(\rs_out<13> ), .B(n50), .Y(n36) );
  INVX1 U66 ( .A(n36), .Y(n37) );
  AND2X2 U75 ( .A(n152), .B(n112), .Y(n38) );
  BUFX2 U76 ( .A(\Instr<0> ), .Y(n39) );
  BUFX2 U78 ( .A(\Instr<1> ), .Y(n40) );
  BUFX2 U79 ( .A(n184), .Y(Halt) );
  BUFX2 U80 ( .A(n183), .Y(Btr) );
  BUFX2 U81 ( .A(n182), .Y(JumpReg) );
  BUFX2 U84 ( .A(n153), .Y(n44) );
  BUFX2 U85 ( .A(\Instr<6> ), .Y(n45) );
  BUFX2 U86 ( .A(\Instr<7> ), .Y(n46) );
  AND2X2 U89 ( .A(\rs_out<6> ), .B(n38), .Y(n47) );
  INVX1 U94 ( .A(n47), .Y(n48) );
  INVX4 U95 ( .A(n113), .Y(\Func<1> ) );
  BUFX2 U96 ( .A(n46), .Y(n49) );
  INVX1 U97 ( .A(lbi), .Y(n152) );
  AND2X2 U98 ( .A(n107), .B(n111), .Y(n50) );
  INVX1 U99 ( .A(n1), .Y(n51) );
  AND2X2 U100 ( .A(n107), .B(n111), .Y(n52) );
  BUFX2 U101 ( .A(\Instr<11> ), .Y(\Func<0> ) );
  INVX1 U102 ( .A(n104), .Y(n54) );
  OR2X1 U103 ( .A(n117), .B(n71), .Y(n55) );
  OR2X1 U104 ( .A(n97), .B(n57), .Y(n56) );
  OR2X1 U105 ( .A(n65), .B(n86), .Y(n57) );
  OR2X1 U106 ( .A(n92), .B(n59), .Y(n58) );
  OR2X1 U107 ( .A(n55), .B(n83), .Y(n59) );
  OR2X1 U108 ( .A(n93), .B(n62), .Y(n61) );
  OR2X1 U109 ( .A(n63), .B(n98), .Y(n62) );
  OR2X1 U110 ( .A(ZeroExt), .B(If1), .Y(n63) );
  OR2X2 U111 ( .A(ZeroExt), .B(Jump), .Y(n65) );
  AND2X1 U112 ( .A(n90), .B(n109), .Y(n66) );
  INVX1 U113 ( .A(n66), .Y(n67) );
  AND2X1 U114 ( .A(n90), .B(n115), .Y(n68) );
  INVX1 U115 ( .A(n68), .Y(n72) );
  INVX1 U116 ( .A(n73), .Y(n74) );
  BUFX2 U117 ( .A(n64), .Y(n75) );
  INVX1 U118 ( .A(n75), .Y(n172) );
  BUFX2 U119 ( .A(n79), .Y(n76) );
  BUFX2 U120 ( .A(n77), .Y(n78) );
  BUFX2 U121 ( .A(n69), .Y(n80) );
  AND2X1 U122 ( .A(n88), .B(n98), .Y(n81) );
  INVX1 U123 ( .A(n81), .Y(n82) );
  AND2X1 U124 ( .A(n88), .B(n175), .Y(n83) );
  INVX1 U125 ( .A(n83), .Y(n84) );
  AND2X1 U126 ( .A(If1), .B(n173), .Y(n85) );
  INVX1 U127 ( .A(n85), .Y(n86) );
  OR2X1 U128 ( .A(n173), .B(If1), .Y(n87) );
  INVX1 U129 ( .A(n87), .Y(n88) );
  INVX1 U130 ( .A(n89), .Y(n90) );
  INVX1 U131 ( .A(n92), .Y(n91) );
  AND2X1 U132 ( .A(n85), .B(n175), .Y(n92) );
  INVX1 U133 ( .A(n93), .Y(n94) );
  AND2X2 U134 ( .A(n15), .B(n48), .Y(n95) );
  INVX4 U135 ( .A(n95), .Y(\ALUOp1<14> ) );
  INVX1 U136 ( .A(\Instr<4> ), .Y(n97) );
  INVX1 U137 ( .A(Jump), .Y(n98) );
  INVX1 U138 ( .A(n49), .Y(n181) );
  INVX1 U139 ( .A(\Instr<12> ), .Y(n113) );
  INVX1 U140 ( .A(\rs_out<2> ), .Y(n99) );
  INVX1 U141 ( .A(n99), .Y(n100) );
  INVX1 U142 ( .A(\WriteData<13> ), .Y(n125) );
  INVX4 U143 ( .A(n44), .Y(\ALUOp1<15> ) );
  INVX1 U144 ( .A(\WriteData<10> ), .Y(n131) );
  INVX1 U145 ( .A(\rs_out<3> ), .Y(n101) );
  INVX1 U146 ( .A(n101), .Y(n102) );
  INVX1 U147 ( .A(n109), .Y(n103) );
  INVX1 U148 ( .A(\Instr<5> ), .Y(n119) );
  INVX1 U149 ( .A(\WriteData<11> ), .Y(n129) );
  INVX4 U150 ( .A(n119), .Y(n118) );
  INVX1 U151 ( .A(n38), .Y(n104) );
  INVX1 U152 ( .A(\WriteData<9> ), .Y(n133) );
  INVX1 U153 ( .A(\WriteData<8> ), .Y(n135) );
  INVX1 U154 ( .A(\WriteData<15> ), .Y(n121) );
  INVX1 U155 ( .A(lbi), .Y(n107) );
  BUFX2 U156 ( .A(\Instr<8> ), .Y(n105) );
  INVX1 U157 ( .A(n51), .Y(n106) );
  BUFX2 U158 ( .A(\Instr<9> ), .Y(n108) );
  INVX1 U159 ( .A(\WriteData<12> ), .Y(n127) );
  BUFX2 U160 ( .A(n118), .Y(n109) );
  AND2X2 U161 ( .A(n17), .B(n19), .Y(n110) );
  INVX1 U162 ( .A(slbi), .Y(n111) );
  INVX1 U163 ( .A(n111), .Y(n112) );
  INVX1 U164 ( .A(\WriteData<14> ), .Y(n123) );
  INVX1 U165 ( .A(n115), .Y(n180) );
  INVX1 U166 ( .A(n108), .Y(n178) );
  INVX1 U167 ( .A(n105), .Y(n179) );
  BUFX2 U168 ( .A(n45), .Y(n115) );
  INVX1 U169 ( .A(\WriteData<1> ), .Y(n149) );
  INVX1 U170 ( .A(\WriteData<2> ), .Y(n147) );
  INVX1 U171 ( .A(\WriteData<0> ), .Y(n151) );
  INVX1 U172 ( .A(\WriteData<4> ), .Y(n143) );
  INVX1 U173 ( .A(\WriteData<3> ), .Y(n145) );
  INVX1 U174 ( .A(\WriteData<6> ), .Y(n139) );
  INVX1 U175 ( .A(\WriteData<5> ), .Y(n141) );
  INVX1 U176 ( .A(\WriteData<7> ), .Y(n137) );
  BUFX4 U177 ( .A(link), .Y(n116) );
  BUFX4 U178 ( .A(link), .Y(n117) );
  MUX2X1 U179 ( .B(n121), .A(n120), .S(n116), .Y(n170) );
  MUX2X1 U180 ( .B(n123), .A(n122), .S(n116), .Y(n169) );
  MUX2X1 U181 ( .B(n125), .A(n124), .S(n116), .Y(n168) );
  MUX2X1 U182 ( .B(n127), .A(n126), .S(n116), .Y(n167) );
  MUX2X1 U183 ( .B(n129), .A(n128), .S(n116), .Y(n166) );
  MUX2X1 U184 ( .B(n131), .A(n130), .S(n116), .Y(n165) );
  MUX2X1 U185 ( .B(n133), .A(n132), .S(n116), .Y(n164) );
  MUX2X1 U186 ( .B(n135), .A(n134), .S(n116), .Y(n163) );
  MUX2X1 U187 ( .B(n137), .A(n136), .S(n116), .Y(n162) );
  MUX2X1 U188 ( .B(n139), .A(n138), .S(n117), .Y(n161) );
  MUX2X1 U189 ( .B(n141), .A(n140), .S(n117), .Y(n160) );
  MUX2X1 U190 ( .B(n143), .A(n142), .S(n117), .Y(n159) );
  MUX2X1 U191 ( .B(n145), .A(n144), .S(n117), .Y(n158) );
  MUX2X1 U192 ( .B(n147), .A(n146), .S(n117), .Y(n157) );
  MUX2X1 U193 ( .B(n149), .A(n148), .S(n117), .Y(n156) );
  MUX2X1 U194 ( .B(n151), .A(n150), .S(n117), .Y(n155) );
  AND2X2 U195 ( .A(n50), .B(\rs_out<0> ), .Y(\ALUOp1<0> ) );
  AND2X2 U196 ( .A(n50), .B(\rs_out<1> ), .Y(\ALUOp1<1> ) );
  AND2X2 U197 ( .A(n52), .B(\rs_out<2> ), .Y(\ALUOp1<2> ) );
  AND2X2 U198 ( .A(n50), .B(\rs_out<3> ), .Y(\ALUOp1<3> ) );
  AND2X2 U199 ( .A(n50), .B(\rs_out<4> ), .Y(\ALUOp1<4> ) );
  AND2X2 U200 ( .A(n50), .B(\rs_out<5> ), .Y(\ALUOp1<5> ) );
  AND2X2 U201 ( .A(n52), .B(\rs_out<6> ), .Y(\ALUOp1<6> ) );
  AND2X2 U202 ( .A(n52), .B(\rs_out<7> ), .Y(\ALUOp1<7> ) );
  AOI22X1 U203 ( .A(n106), .B(n38), .C(\rs_out<15> ), .D(n50), .Y(n153) );
endmodule


module execute ( .ALUOp1({\ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , 
        \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , 
        \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , 
        \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), .ALUOp2({\ALUOp2<15> , 
        \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , 
        \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , 
        \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), 
    .Opcode({\Opcode<2> , \Opcode<1> , \Opcode<0> }), .IncPC({\IncPC<15> , 
        \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , 
        \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , 
        \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> }), Jump, Branch, 
        JumpReg, Set, InvA, InvB, Cin, Btr, .Func({\Func<1> , \Func<0> }), 
    .Imm({\Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> , \Imm<11> , \Imm<10> , 
        \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> , \Imm<5> , \Imm<4> , \Imm<3> , 
        \Imm<2> , \Imm<1> , \Imm<0> }), ALUSrc, .Result({\Result<15> , 
        \Result<14> , \Result<13> , \Result<12> , \Result<11> , \Result<10> , 
        \Result<9> , \Result<8> , \Result<7> , \Result<6> , \Result<5> , 
        \Result<4> , \Result<3> , \Result<2> , \Result<1> , \Result<0> }), 
    .NextPC({\NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> , 
        \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> , 
        \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> , 
        \NextPC<1> , \NextPC<0> }) );
  input \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> ,
         \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> ,
         \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> ,
         \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , \Opcode<2> , \Opcode<1> , \Opcode<0> ,
         \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> ,
         \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> ,
         \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> ,
         \IncPC<0> , Jump, Branch, JumpReg, Set, InvA, InvB, Cin, Btr,
         \Func<1> , \Func<0> , \Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> ,
         \Imm<11> , \Imm<10> , \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> ,
         \Imm<5> , \Imm<4> , \Imm<3> , \Imm<2> , \Imm<1> , \Imm<0> , ALUSrc;
  output \Result<15> , \Result<14> , \Result<13> , \Result<12> , \Result<11> ,
         \Result<10> , \Result<9> , \Result<8> , \Result<7> , \Result<6> ,
         \Result<5> , \Result<4> , \Result<3> , \Result<2> , \Result<1> ,
         \Result<0> , \NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> ,
         \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> ,
         \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> ,
         \NextPC<1> , \NextPC<0> ;
  wire   n323, \_0_net_<15> , \aluResult<15> , \aluResult<14> ,
         \aluResult<13> , \aluResult<12> , \aluResult<11> , \aluResult<10> ,
         \aluResult<9> , \aluResult<8> , \aluResult<7> , \aluResult<6> ,
         \aluResult<5> , \aluResult<4> , \aluResult<3> , \aluResult<2> ,
         \aluResult<1> , \aluResult<0> , Zero, cout, \_3_net_<0> ,
         \setResult<15> , \setResult<14> , \setResult<13> , \setResult<12> ,
         \setResult<11> , \setResult<10> , \setResult<9> , \setResult<8> ,
         \setResult<7> , \setResult<6> , \setResult<5> , \setResult<4> ,
         \setResult<3> , \setResult<2> , \setResult<1> , \setResult<0> ,
         \offsetAddr<15> , \offsetAddr<14> , \offsetAddr<13> ,
         \offsetAddr<12> , \offsetAddr<11> , \offsetAddr<10> , \offsetAddr<9> ,
         \offsetAddr<8> , \offsetAddr<7> , \offsetAddr<6> , \offsetAddr<5> ,
         \offsetAddr<4> , \offsetAddr<3> , \offsetAddr<2> , \offsetAddr<1> ,
         \offsetAddr<0> , branch_en, _8_net_, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n21, n23, n25, n27,
         n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n125, n127, n130, n131, n132, n133,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322;

  alu primary_alu ( .A({\ALUOp1<15> , \ALUOp1<14> , n137, n140, n135, n218, 
        \ALUOp1<9> , n219, \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , 
        \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), .B({
        \_0_net_<15> , n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316, n317, n318, n319, n320}), .Cin(Cin), .Op({\Opcode<2> , 
        \Opcode<1> , \Opcode<0> }), .invA(InvA), .invB(InvB), .sign(1'b1), 
        .Out({\aluResult<15> , \aluResult<14> , \aluResult<13> , 
        \aluResult<12> , \aluResult<11> , \aluResult<10> , \aluResult<9> , 
        \aluResult<8> , \aluResult<7> , \aluResult<6> , \aluResult<5> , 
        \aluResult<4> , \aluResult<3> , \aluResult<2> , \aluResult<1> , 
        \aluResult<0> }), .Ofl(), .Z(Zero), .Cout(cout) );
  mux4to1_16_5 set_mux ( .InA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n230}), .InB({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \_3_net_<0> }), .InC({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n14}), .InD({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout}), .S({\Func<1> , \Func<0> }), .Out({\setResult<15> , 
        \setResult<14> , \setResult<13> , \setResult<12> , \setResult<11> , 
        \setResult<10> , \setResult<9> , \setResult<8> , \setResult<7> , 
        \setResult<6> , \setResult<5> , \setResult<4> , \setResult<3> , 
        \setResult<2> , \setResult<1> , \setResult<0> }) );
  cla16_1 addr_adder ( .A({\IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , 
        \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , 
        \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> , 
        \IncPC<0> }), .B({\Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> , 
        \Imm<11> , \Imm<10> , \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> , \Imm<5> , 
        \Imm<4> , \Imm<3> , \Imm<2> , \Imm<1> , \Imm<0> }), .Cin(1'b0), .S({
        \offsetAddr<15> , \offsetAddr<14> , \offsetAddr<13> , \offsetAddr<12> , 
        \offsetAddr<11> , \offsetAddr<10> , \offsetAddr<9> , \offsetAddr<8> , 
        \offsetAddr<7> , \offsetAddr<6> , \offsetAddr<5> , \offsetAddr<4> , 
        \offsetAddr<3> , \offsetAddr<2> , \offsetAddr<1> , \offsetAddr<0> }), 
        .Cout() );
  mux4to1 branchMux ( .InA(n321), .InB(n130), .InC(\ALUOp1<15> ), .InD(n322), 
        .S({\Func<1> , \Func<0> }), .Out(branch_en) );
  MUX2X1 U3 ( .B(n245), .A(n261), .S(n238), .Y(n310) );
  MUX2X1 U4 ( .B(n242), .A(n258), .S(ALUSrc), .Y(n313) );
  INVX2 U5 ( .A(n232), .Y(n318) );
  INVX1 U6 ( .A(Zero), .Y(n1) );
  AND2X1 U7 ( .A(n65), .B(n92), .Y(n187) );
  INVX1 U8 ( .A(Jump), .Y(n267) );
  INVX1 U9 ( .A(n10), .Y(\Result<7> ) );
  INVX1 U10 ( .A(n224), .Y(n7) );
  INVX1 U11 ( .A(\Imm<8> ), .Y(n259) );
  INVX1 U12 ( .A(\Imm<9> ), .Y(n260) );
  INVX1 U13 ( .A(\Imm<0> ), .Y(n256) );
  INVX1 U14 ( .A(\ALUOp1<15> ), .Y(n322) );
  INVX1 U15 ( .A(\Imm<11> ), .Y(n262) );
  INVX1 U16 ( .A(\Imm<15> ), .Y(n266) );
  AND2X1 U17 ( .A(n109), .B(n160), .Y(n43) );
  AND2X1 U18 ( .A(n180), .B(n161), .Y(n45) );
  INVX1 U19 ( .A(\Imm<4> ), .Y(n257) );
  INVX1 U20 ( .A(\Imm<7> ), .Y(n258) );
  INVX1 U21 ( .A(\Imm<10> ), .Y(n261) );
  INVX1 U22 ( .A(\Imm<12> ), .Y(n263) );
  INVX1 U23 ( .A(\Imm<13> ), .Y(n264) );
  AND2X1 U24 ( .A(n74), .B(n60), .Y(n144) );
  INVX1 U25 ( .A(n237), .Y(n238) );
  INVX1 U26 ( .A(\ALUOp2<15> ), .Y(n250) );
  BUFX2 U27 ( .A(\aluResult<5> ), .Y(n2) );
  MUX2X1 U28 ( .B(n264), .A(n248), .S(n214), .Y(n307) );
  NOR3X1 U29 ( .A(n200), .B(n195), .C(n123), .Y(n3) );
  INVX1 U30 ( .A(n3), .Y(\Result<10> ) );
  AND2X2 U31 ( .A(\aluResult<10> ), .B(n303), .Y(n123) );
  MUX2X1 U32 ( .B(n265), .A(n249), .S(n4), .Y(n306) );
  INVX8 U33 ( .A(n207), .Y(n4) );
  MUX2X1 U34 ( .B(n260), .A(n244), .S(n215), .Y(n311) );
  BUFX2 U35 ( .A(\aluResult<10> ), .Y(n5) );
  MUX2X1 U36 ( .B(\ALUOp2<3> ), .A(\Imm<3> ), .S(ALUSrc), .Y(n233) );
  INVX1 U37 ( .A(n6), .Y(n314) );
  INVX1 U38 ( .A(n231), .Y(n315) );
  MUX2X1 U39 ( .B(\Imm<2> ), .A(\ALUOp2<2> ), .S(n220), .Y(n232) );
  AND2X2 U40 ( .A(\aluResult<9> ), .B(n303), .Y(n121) );
  MUX2X1 U41 ( .B(\Imm<6> ), .A(\ALUOp2<6> ), .S(n217), .Y(n6) );
  INVX1 U42 ( .A(n233), .Y(n317) );
  MUX2X1 U43 ( .B(n246), .A(n262), .S(n7), .Y(n309) );
  INVX1 U44 ( .A(n9), .Y(n319) );
  NOR3X1 U45 ( .A(n199), .B(n194), .C(n121), .Y(n8) );
  INVX1 U46 ( .A(n8), .Y(\Result<9> ) );
  MUX2X1 U47 ( .B(\Imm<1> ), .A(\ALUOp2<1> ), .S(n220), .Y(n9) );
  MUX2X1 U48 ( .B(\Imm<5> ), .A(\ALUOp2<5> ), .S(n237), .Y(n231) );
  NOR3X1 U49 ( .A(n198), .B(n193), .C(n118), .Y(n10) );
  MUX2X1 U50 ( .B(n241), .A(n257), .S(n208), .Y(n316) );
  AND2X2 U51 ( .A(n303), .B(\aluResult<12> ), .Y(n63) );
  AND2X1 U52 ( .A(\aluResult<8> ), .B(n303), .Y(n87) );
  MUX2X1 U53 ( .B(n240), .A(n256), .S(n216), .Y(n320) );
  OR2X2 U54 ( .A(\ALUOp1<9> ), .B(\ALUOp1<8> ), .Y(n11) );
  INVX1 U55 ( .A(n11), .Y(n12) );
  AND2X2 U56 ( .A(n1), .B(n254), .Y(n13) );
  INVX1 U57 ( .A(n13), .Y(n14) );
  OR2X2 U58 ( .A(JumpReg), .B(Jump), .Y(n15) );
  INVX1 U59 ( .A(n15), .Y(n16) );
  AND2X2 U60 ( .A(n99), .B(n147), .Y(n17) );
  INVX1 U61 ( .A(n17), .Y(\NextPC<0> ) );
  AND2X2 U62 ( .A(n164), .B(n148), .Y(n19) );
  INVX1 U63 ( .A(n19), .Y(\NextPC<1> ) );
  AND2X2 U64 ( .A(n166), .B(n149), .Y(n21) );
  INVX1 U65 ( .A(n21), .Y(\NextPC<2> ) );
  AND2X2 U66 ( .A(n168), .B(n150), .Y(n23) );
  INVX1 U67 ( .A(n23), .Y(\NextPC<3> ) );
  AND2X2 U68 ( .A(n170), .B(n151), .Y(n25) );
  INVX1 U69 ( .A(n25), .Y(\NextPC<4> ) );
  AND2X2 U70 ( .A(n172), .B(n152), .Y(n27) );
  INVX1 U71 ( .A(n27), .Y(\NextPC<5> ) );
  AND2X2 U72 ( .A(n174), .B(n153), .Y(n29) );
  INVX1 U73 ( .A(n29), .Y(\NextPC<6> ) );
  AND2X2 U74 ( .A(n176), .B(n154), .Y(n31) );
  INVX1 U75 ( .A(n31), .Y(\NextPC<7> ) );
  AND2X2 U76 ( .A(n101), .B(n155), .Y(n33) );
  INVX1 U77 ( .A(n33), .Y(\NextPC<8> ) );
  AND2X2 U78 ( .A(n103), .B(n156), .Y(n35) );
  INVX1 U79 ( .A(n35), .Y(\NextPC<9> ) );
  AND2X2 U80 ( .A(n178), .B(n157), .Y(n37) );
  INVX1 U81 ( .A(n37), .Y(\NextPC<10> ) );
  AND2X2 U82 ( .A(n105), .B(n158), .Y(n39) );
  INVX1 U83 ( .A(n39), .Y(\NextPC<11> ) );
  AND2X2 U84 ( .A(n107), .B(n159), .Y(n41) );
  INVX1 U85 ( .A(n41), .Y(\NextPC<12> ) );
  INVX1 U86 ( .A(n43), .Y(\NextPC<13> ) );
  INVX1 U87 ( .A(n45), .Y(\NextPC<14> ) );
  AND2X2 U88 ( .A(n111), .B(n162), .Y(n47) );
  INVX1 U89 ( .A(n47), .Y(\NextPC<15> ) );
  OR2X2 U90 ( .A(n186), .B(n63), .Y(\Result<12> ) );
  OR2X2 U91 ( .A(n226), .B(n227), .Y(n50) );
  OR2X2 U92 ( .A(\ALUOp1<1> ), .B(\ALUOp1<0> ), .Y(n51) );
  INVX1 U93 ( .A(n51), .Y(n52) );
  OR2X2 U94 ( .A(n206), .B(\ALUOp1<7> ), .Y(n53) );
  INVX1 U95 ( .A(n53), .Y(n54) );
  AND2X2 U96 ( .A(n54), .B(n97), .Y(n55) );
  INVX1 U97 ( .A(n55), .Y(n56) );
  OR2X2 U98 ( .A(n113), .B(n56), .Y(n57) );
  INVX1 U99 ( .A(n57), .Y(n58) );
  AND2X2 U100 ( .A(Btr), .B(\ALUOp1<7> ), .Y(n59) );
  INVX1 U101 ( .A(n59), .Y(n60) );
  AND2X2 U102 ( .A(\setResult<11> ), .B(n304), .Y(n61) );
  INVX1 U103 ( .A(n61), .Y(n62) );
  AND2X2 U104 ( .A(\setResult<14> ), .B(n304), .Y(n64) );
  INVX1 U105 ( .A(n64), .Y(n65) );
  BUFX2 U106 ( .A(n302), .Y(n66) );
  OR2X2 U107 ( .A(\ALUOp1<15> ), .B(\ALUOp1<14> ), .Y(n67) );
  INVX1 U108 ( .A(n67), .Y(n68) );
  OR2X2 U109 ( .A(n142), .B(n223), .Y(n69) );
  INVX1 U110 ( .A(n69), .Y(n70) );
  OR2X2 U111 ( .A(n210), .B(\ALUOp1<2> ), .Y(n71) );
  INVX1 U112 ( .A(n71), .Y(n72) );
  AND2X2 U113 ( .A(\setResult<8> ), .B(n304), .Y(n73) );
  INVX1 U114 ( .A(n73), .Y(n74) );
  AND2X2 U115 ( .A(Btr), .B(n211), .Y(n75) );
  INVX1 U116 ( .A(n75), .Y(n76) );
  AND2X2 U117 ( .A(Btr), .B(n210), .Y(n77) );
  INVX1 U118 ( .A(n77), .Y(n78) );
  AND2X2 U119 ( .A(Btr), .B(\ALUOp1<2> ), .Y(n79) );
  INVX1 U120 ( .A(n79), .Y(n80) );
  OR2X2 U121 ( .A(n138), .B(n141), .Y(n81) );
  INVX1 U122 ( .A(n81), .Y(n82) );
  AND2X1 U123 ( .A(\aluResult<1> ), .B(n303), .Y(n83) );
  INVX1 U124 ( .A(n83), .Y(n84) );
  AND2X1 U125 ( .A(\aluResult<5> ), .B(n303), .Y(n85) );
  INVX1 U126 ( .A(n85), .Y(n86) );
  INVX1 U127 ( .A(n87), .Y(n88) );
  AND2X2 U128 ( .A(\setResult<13> ), .B(n304), .Y(n89) );
  INVX1 U129 ( .A(n89), .Y(n90) );
  AND2X2 U130 ( .A(\ALUOp1<1> ), .B(Btr), .Y(n91) );
  INVX1 U131 ( .A(n91), .Y(n92) );
  BUFX2 U132 ( .A(n292), .Y(n93) );
  BUFX2 U133 ( .A(n295), .Y(n94) );
  BUFX2 U134 ( .A(n298), .Y(n95) );
  OR2X2 U135 ( .A(n209), .B(n211), .Y(n96) );
  INVX1 U136 ( .A(n96), .Y(n97) );
  AND2X2 U137 ( .A(JumpReg), .B(\aluResult<0> ), .Y(n98) );
  INVX1 U138 ( .A(n98), .Y(n99) );
  AND2X2 U139 ( .A(n239), .B(\aluResult<8> ), .Y(n100) );
  INVX1 U140 ( .A(n100), .Y(n101) );
  AND2X2 U141 ( .A(n239), .B(n213), .Y(n102) );
  INVX1 U142 ( .A(n102), .Y(n103) );
  AND2X2 U143 ( .A(n239), .B(\aluResult<11> ), .Y(n104) );
  INVX1 U144 ( .A(n104), .Y(n105) );
  AND2X2 U145 ( .A(n239), .B(n212), .Y(n106) );
  INVX1 U146 ( .A(n106), .Y(n107) );
  AND2X2 U147 ( .A(n239), .B(\aluResult<13> ), .Y(n108) );
  INVX1 U148 ( .A(n108), .Y(n109) );
  AND2X2 U149 ( .A(JumpReg), .B(n229), .Y(n110) );
  INVX1 U150 ( .A(n110), .Y(n111) );
  AND2X2 U151 ( .A(n72), .B(n52), .Y(n112) );
  INVX1 U152 ( .A(n112), .Y(n113) );
  AND2X2 U153 ( .A(n182), .B(n84), .Y(n114) );
  INVX1 U154 ( .A(n114), .Y(n115) );
  AND2X2 U155 ( .A(n184), .B(n86), .Y(n116) );
  INVX1 U156 ( .A(n116), .Y(n117) );
  AND2X2 U157 ( .A(n303), .B(\aluResult<7> ), .Y(n118) );
  AND2X1 U158 ( .A(\aluResult<6> ), .B(n303), .Y(n119) );
  INVX1 U159 ( .A(n119), .Y(n120) );
  BUFX2 U160 ( .A(n290), .Y(n122) );
  BUFX2 U161 ( .A(n305), .Y(\Result<0> ) );
  AND2X2 U162 ( .A(n66), .B(n143), .Y(n125) );
  INVX1 U163 ( .A(n125), .Y(\Result<11> ) );
  AND2X2 U164 ( .A(n144), .B(n88), .Y(n127) );
  INVX1 U165 ( .A(n127), .Y(\Result<8> ) );
  BUFX2 U166 ( .A(n323), .Y(\Result<6> ) );
  BUFX2 U167 ( .A(_8_net_), .Y(n130) );
  AND2X2 U168 ( .A(Branch), .B(branch_en), .Y(n131) );
  INVX1 U169 ( .A(n131), .Y(n132) );
  INVX1 U170 ( .A(n131), .Y(n133) );
  OR2X2 U171 ( .A(n50), .B(n225), .Y(\Result<15> ) );
  BUFX2 U172 ( .A(\ALUOp1<11> ), .Y(n135) );
  INVX2 U173 ( .A(n122), .Y(\Result<1> ) );
  INVX1 U174 ( .A(\ALUOp1<13> ), .Y(n136) );
  INVX1 U175 ( .A(n136), .Y(n137) );
  INVX1 U176 ( .A(n136), .Y(n138) );
  INVX1 U177 ( .A(\ALUOp1<12> ), .Y(n139) );
  INVX1 U178 ( .A(n139), .Y(n140) );
  INVX1 U179 ( .A(n139), .Y(n141) );
  BUFX2 U180 ( .A(n135), .Y(n142) );
  INVX1 U181 ( .A(n138), .Y(n293) );
  INVX1 U182 ( .A(n141), .Y(n296) );
  AND2X2 U183 ( .A(n76), .B(n62), .Y(n143) );
  AND2X2 U184 ( .A(\setResult<12> ), .B(n304), .Y(n145) );
  INVX1 U185 ( .A(n145), .Y(n146) );
  INVX8 U186 ( .A(n289), .Y(n304) );
  BUFX2 U187 ( .A(n268), .Y(n147) );
  BUFX2 U188 ( .A(n269), .Y(n148) );
  BUFX2 U189 ( .A(n270), .Y(n149) );
  BUFX2 U190 ( .A(n271), .Y(n150) );
  BUFX2 U191 ( .A(n272), .Y(n151) );
  BUFX2 U192 ( .A(n273), .Y(n152) );
  BUFX2 U193 ( .A(n274), .Y(n153) );
  BUFX2 U194 ( .A(n275), .Y(n154) );
  BUFX2 U195 ( .A(n276), .Y(n155) );
  BUFX2 U196 ( .A(n277), .Y(n156) );
  BUFX2 U197 ( .A(n278), .Y(n157) );
  BUFX2 U198 ( .A(n279), .Y(n158) );
  BUFX2 U199 ( .A(n280), .Y(n159) );
  BUFX2 U200 ( .A(n281), .Y(n160) );
  BUFX2 U201 ( .A(n282), .Y(n161) );
  BUFX2 U202 ( .A(n285), .Y(n162) );
  AND2X2 U203 ( .A(\aluResult<1> ), .B(JumpReg), .Y(n163) );
  INVX1 U204 ( .A(n163), .Y(n164) );
  AND2X2 U205 ( .A(\aluResult<2> ), .B(JumpReg), .Y(n165) );
  INVX1 U206 ( .A(n165), .Y(n166) );
  AND2X2 U207 ( .A(\aluResult<3> ), .B(JumpReg), .Y(n167) );
  INVX1 U208 ( .A(n167), .Y(n168) );
  AND2X2 U209 ( .A(\aluResult<4> ), .B(JumpReg), .Y(n169) );
  INVX1 U210 ( .A(n169), .Y(n170) );
  AND2X2 U211 ( .A(n2), .B(JumpReg), .Y(n171) );
  INVX1 U212 ( .A(n171), .Y(n172) );
  AND2X2 U213 ( .A(\aluResult<6> ), .B(n239), .Y(n173) );
  INVX1 U214 ( .A(n173), .Y(n174) );
  AND2X2 U215 ( .A(\aluResult<7> ), .B(n239), .Y(n175) );
  INVX1 U216 ( .A(n175), .Y(n176) );
  AND2X2 U217 ( .A(n5), .B(n239), .Y(n177) );
  INVX1 U218 ( .A(n177), .Y(n178) );
  AND2X2 U219 ( .A(\aluResult<14> ), .B(n239), .Y(n179) );
  INVX1 U220 ( .A(n179), .Y(n180) );
  AND2X2 U221 ( .A(\setResult<1> ), .B(n304), .Y(n181) );
  INVX1 U222 ( .A(n181), .Y(n182) );
  AND2X2 U223 ( .A(\setResult<5> ), .B(n304), .Y(n183) );
  INVX1 U224 ( .A(n183), .Y(n184) );
  AND2X2 U225 ( .A(n78), .B(n146), .Y(n185) );
  INVX1 U226 ( .A(n185), .Y(n186) );
  INVX1 U227 ( .A(n187), .Y(n188) );
  AND2X2 U228 ( .A(n80), .B(n90), .Y(n189) );
  INVX1 U229 ( .A(n189), .Y(n190) );
  AND2X2 U230 ( .A(\setResult<6> ), .B(n304), .Y(n191) );
  INVX1 U231 ( .A(n191), .Y(n192) );
  AND2X2 U232 ( .A(\setResult<7> ), .B(n304), .Y(n193) );
  AND2X2 U233 ( .A(\setResult<9> ), .B(n304), .Y(n194) );
  AND2X2 U234 ( .A(\setResult<10> ), .B(n304), .Y(n195) );
  AND2X2 U235 ( .A(Btr), .B(\ALUOp1<9> ), .Y(n196) );
  INVX1 U236 ( .A(n196), .Y(n197) );
  AND2X2 U237 ( .A(Btr), .B(\ALUOp1<8> ), .Y(n198) );
  AND2X2 U238 ( .A(Btr), .B(\ALUOp1<6> ), .Y(n199) );
  AND2X2 U239 ( .A(Btr), .B(n209), .Y(n200) );
  INVX1 U240 ( .A(n130), .Y(n321) );
  BUFX2 U241 ( .A(n288), .Y(n201) );
  BUFX2 U242 ( .A(JumpReg), .Y(n239) );
  BUFX2 U243 ( .A(n283), .Y(n236) );
  AOI21X1 U244 ( .A(\aluResult<14> ), .B(n303), .C(n188), .Y(n202) );
  INVX1 U245 ( .A(n202), .Y(\Result<14> ) );
  INVX1 U246 ( .A(n286), .Y(n303) );
  NAND3X1 U247 ( .A(n299), .B(n203), .C(\aluResult<11> ), .Y(n302) );
  INVX1 U248 ( .A(Set), .Y(n203) );
  AOI21X1 U249 ( .A(\aluResult<13> ), .B(n303), .C(n190), .Y(n204) );
  INVX1 U250 ( .A(n204), .Y(\Result<13> ) );
  INVX1 U251 ( .A(\ALUOp1<6> ), .Y(n205) );
  INVX1 U252 ( .A(n205), .Y(n206) );
  INVX1 U253 ( .A(n215), .Y(n207) );
  INVX1 U254 ( .A(n237), .Y(n208) );
  BUFX2 U255 ( .A(\ALUOp1<5> ), .Y(n209) );
  BUFX2 U256 ( .A(\ALUOp1<3> ), .Y(n210) );
  BUFX2 U257 ( .A(\ALUOp1<4> ), .Y(n211) );
  BUFX2 U258 ( .A(\aluResult<12> ), .Y(n212) );
  BUFX2 U259 ( .A(\aluResult<9> ), .Y(n213) );
  INVX1 U260 ( .A(\ALUOp1<8> ), .Y(n221) );
  INVX2 U261 ( .A(ALUSrc), .Y(n237) );
  INVX1 U262 ( .A(n216), .Y(n214) );
  MUX2X1 U263 ( .B(n259), .A(n243), .S(n214), .Y(n312) );
  INVX1 U264 ( .A(n208), .Y(n224) );
  INVX1 U265 ( .A(n142), .Y(n300) );
  INVX1 U266 ( .A(ALUSrc), .Y(n215) );
  INVX1 U267 ( .A(n237), .Y(n216) );
  INVX1 U268 ( .A(ALUSrc), .Y(n220) );
  INVX1 U269 ( .A(n208), .Y(n217) );
  INVX1 U270 ( .A(\ALUOp2<9> ), .Y(n244) );
  INVX1 U271 ( .A(n222), .Y(n218) );
  INVX1 U272 ( .A(n221), .Y(n219) );
  INVX1 U273 ( .A(\ALUOp2<10> ), .Y(n245) );
  INVX1 U274 ( .A(\ALUOp2<12> ), .Y(n247) );
  INVX1 U275 ( .A(\ALUOp2<8> ), .Y(n243) );
  INVX1 U276 ( .A(\ALUOp2<14> ), .Y(n249) );
  INVX1 U277 ( .A(\ALUOp1<10> ), .Y(n222) );
  INVX1 U278 ( .A(n222), .Y(n223) );
  AND2X2 U279 ( .A(\aluResult<15> ), .B(n303), .Y(n225) );
  AND2X2 U280 ( .A(\setResult<15> ), .B(n304), .Y(n226) );
  AND2X2 U281 ( .A(Btr), .B(\ALUOp1<0> ), .Y(n227) );
  INVX1 U282 ( .A(\ALUOp2<13> ), .Y(n248) );
  INVX1 U283 ( .A(\aluResult<15> ), .Y(n228) );
  INVX1 U284 ( .A(n228), .Y(n229) );
  INVX1 U285 ( .A(n301), .Y(\Result<5> ) );
  INVX1 U286 ( .A(n254), .Y(\_3_net_<0> ) );
  INVX1 U287 ( .A(n255), .Y(n230) );
  INVX1 U288 ( .A(Zero), .Y(n255) );
  INVX1 U289 ( .A(\ALUOp2<11> ), .Y(n246) );
  INVX1 U290 ( .A(\ALUOp2<4> ), .Y(n241) );
  INVX1 U291 ( .A(\ALUOp2<0> ), .Y(n240) );
  INVX1 U292 ( .A(\ALUOp2<7> ), .Y(n242) );
  INVX1 U293 ( .A(\setResult<0> ), .Y(n287) );
  BUFX4 U294 ( .A(n284), .Y(n234) );
  BUFX4 U295 ( .A(n284), .Y(n235) );
  AND2X2 U296 ( .A(n68), .B(n82), .Y(n252) );
  AND2X2 U297 ( .A(n70), .B(n12), .Y(n251) );
  NAND3X1 U298 ( .A(n252), .B(n251), .C(n58), .Y(_8_net_) );
  XOR2X1 U299 ( .A(\ALUOp2<15> ), .B(\ALUOp1<15> ), .Y(n253) );
  MUX2X1 U300 ( .B(\aluResult<15> ), .A(\ALUOp1<15> ), .S(n253), .Y(n254) );
  MUX2X1 U301 ( .B(n247), .A(n263), .S(n238), .Y(n308) );
  INVX2 U302 ( .A(\Imm<14> ), .Y(n265) );
  MUX2X1 U303 ( .B(n250), .A(n266), .S(n238), .Y(\_0_net_<15> ) );
  AND2X2 U304 ( .A(n133), .B(n16), .Y(n284) );
  AOI21X1 U305 ( .A(n267), .B(n132), .C(JumpReg), .Y(n283) );
  AOI22X1 U306 ( .A(\IncPC<0> ), .B(n234), .C(\offsetAddr<0> ), .D(n236), .Y(
        n268) );
  AOI22X1 U307 ( .A(\IncPC<1> ), .B(n234), .C(\offsetAddr<1> ), .D(n236), .Y(
        n269) );
  AOI22X1 U308 ( .A(\IncPC<2> ), .B(n234), .C(\offsetAddr<2> ), .D(n236), .Y(
        n270) );
  AOI22X1 U309 ( .A(\IncPC<3> ), .B(n234), .C(\offsetAddr<3> ), .D(n236), .Y(
        n271) );
  AOI22X1 U310 ( .A(\IncPC<4> ), .B(n234), .C(\offsetAddr<4> ), .D(n236), .Y(
        n272) );
  AOI22X1 U311 ( .A(\IncPC<5> ), .B(n234), .C(\offsetAddr<5> ), .D(n236), .Y(
        n273) );
  AOI22X1 U312 ( .A(\IncPC<6> ), .B(n234), .C(\offsetAddr<6> ), .D(n236), .Y(
        n274) );
  AOI22X1 U313 ( .A(\IncPC<7> ), .B(n234), .C(\offsetAddr<7> ), .D(n236), .Y(
        n275) );
  AOI22X1 U314 ( .A(\IncPC<8> ), .B(n235), .C(\offsetAddr<8> ), .D(n236), .Y(
        n276) );
  AOI22X1 U315 ( .A(\IncPC<9> ), .B(n235), .C(\offsetAddr<9> ), .D(n236), .Y(
        n277) );
  AOI22X1 U316 ( .A(\IncPC<10> ), .B(n235), .C(\offsetAddr<10> ), .D(n236), 
        .Y(n278) );
  AOI22X1 U317 ( .A(\IncPC<11> ), .B(n235), .C(\offsetAddr<11> ), .D(n236), 
        .Y(n279) );
  AOI22X1 U318 ( .A(\IncPC<12> ), .B(n235), .C(\offsetAddr<12> ), .D(n236), 
        .Y(n280) );
  AOI22X1 U319 ( .A(\IncPC<13> ), .B(n235), .C(\offsetAddr<13> ), .D(n236), 
        .Y(n281) );
  AOI22X1 U320 ( .A(\IncPC<14> ), .B(n235), .C(\offsetAddr<14> ), .D(n236), 
        .Y(n282) );
  AOI22X1 U321 ( .A(\IncPC<15> ), .B(n235), .C(\offsetAddr<15> ), .D(n236), 
        .Y(n285) );
  OR2X2 U322 ( .A(Btr), .B(Set), .Y(n286) );
  AOI22X1 U323 ( .A(Btr), .B(\ALUOp1<15> ), .C(\aluResult<0> ), .D(n303), .Y(
        n288) );
  OR2X2 U324 ( .A(Btr), .B(n203), .Y(n289) );
  AOI22X1 U325 ( .A(n201), .B(n289), .C(n201), .D(n287), .Y(n305) );
  AOI21X1 U326 ( .A(Btr), .B(\ALUOp1<14> ), .C(n115), .Y(n290) );
  INVX2 U327 ( .A(Btr), .Y(n299) );
  AND2X2 U328 ( .A(\setResult<2> ), .B(n304), .Y(n291) );
  AOI21X1 U329 ( .A(\aluResult<2> ), .B(n303), .C(n291), .Y(n292) );
  OAI21X1 U330 ( .A(n293), .B(n299), .C(n93), .Y(\Result<2> ) );
  AND2X2 U331 ( .A(\setResult<3> ), .B(n304), .Y(n294) );
  AOI21X1 U332 ( .A(\aluResult<3> ), .B(n303), .C(n294), .Y(n295) );
  OAI21X1 U333 ( .A(n296), .B(n299), .C(n94), .Y(\Result<3> ) );
  AND2X2 U334 ( .A(\setResult<4> ), .B(n304), .Y(n297) );
  AOI21X1 U335 ( .A(\aluResult<4> ), .B(n303), .C(n297), .Y(n298) );
  OAI21X1 U336 ( .A(n300), .B(n299), .C(n95), .Y(\Result<4> ) );
  AOI21X1 U337 ( .A(Btr), .B(n223), .C(n117), .Y(n301) );
  NAND3X1 U338 ( .A(n120), .B(n192), .C(n197), .Y(n323) );
endmodule


module memory ( MemRead, MemWrite, halt, clk, rst, .Address({\Address<15> , 
        \Address<14> , \Address<13> , \Address<12> , \Address<11> , 
        \Address<10> , \Address<9> , \Address<8> , \Address<7> , \Address<6> , 
        \Address<5> , \Address<4> , \Address<3> , \Address<2> , \Address<1> , 
        \Address<0> }), .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .ReadData({\ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }) );
  input MemRead, MemWrite, halt, clk, rst, \Address<15> , \Address<14> ,
         \Address<13> , \Address<12> , \Address<11> , \Address<10> ,
         \Address<9> , \Address<8> , \Address<7> , \Address<6> , \Address<5> ,
         \Address<4> , \Address<3> , \Address<2> , \Address<1> , \Address<0> ,
         \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ;
  output \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> ,
         \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> ,
         \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> ,
         \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  memory2c_0 data_mem ( .data_out({\ReadData<15> , \ReadData<14> , 
        \ReadData<13> , \ReadData<12> , \ReadData<11> , \ReadData<10> , 
        \ReadData<9> , \ReadData<8> , \ReadData<7> , \ReadData<6> , 
        \ReadData<5> , \ReadData<4> , \ReadData<3> , \ReadData<2> , 
        \ReadData<1> , \ReadData<0> }), .data_in({n17, n15, n13, n11, n9, n7, 
        n5, n3, \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> , 
        \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> }), 
        .addr({\Address<15> , \Address<14> , \Address<13> , \Address<12> , 
        \Address<11> , \Address<10> , \Address<9> , \Address<8> , \Address<7> , 
        \Address<6> , \Address<5> , \Address<4> , \Address<3> , n1, 
        \Address<1> , \Address<0> }), .enable(n19), .wr(MemWrite), 
        .createdump(halt), .clk(clk), .rst(rst) );
  INVX2 U1 ( .A(n4), .Y(n3) );
  INVX2 U2 ( .A(n8), .Y(n7) );
  INVX1 U3 ( .A(\WriteData<8> ), .Y(n4) );
  INVX1 U4 ( .A(n6), .Y(n5) );
  INVX1 U5 ( .A(n10), .Y(n9) );
  INVX1 U6 ( .A(n16), .Y(n15) );
  INVX4 U7 ( .A(n2), .Y(n1) );
  INVX2 U8 ( .A(n12), .Y(n11) );
  INVX2 U9 ( .A(n14), .Y(n13) );
  INVX1 U10 ( .A(\WriteData<13> ), .Y(n14) );
  INVX1 U11 ( .A(\WriteData<14> ), .Y(n16) );
  INVX1 U12 ( .A(\WriteData<12> ), .Y(n12) );
  INVX1 U13 ( .A(halt), .Y(n19) );
  INVX2 U14 ( .A(\Address<2> ), .Y(n2) );
  INVX1 U15 ( .A(\WriteData<9> ), .Y(n6) );
  INVX1 U16 ( .A(\WriteData<11> ), .Y(n10) );
  INVX1 U17 ( .A(\WriteData<10> ), .Y(n8) );
  INVX8 U18 ( .A(n18), .Y(n17) );
  INVX8 U19 ( .A(\WriteData<15> ), .Y(n18) );
endmodule


module writeback ( .ExecuteOut({\ExecuteOut<15> , \ExecuteOut<14> , 
        \ExecuteOut<13> , \ExecuteOut<12> , \ExecuteOut<11> , \ExecuteOut<10> , 
        \ExecuteOut<9> , \ExecuteOut<8> , \ExecuteOut<7> , \ExecuteOut<6> , 
        \ExecuteOut<5> , \ExecuteOut<4> , \ExecuteOut<3> , \ExecuteOut<2> , 
        \ExecuteOut<1> , \ExecuteOut<0> }), .MemOut({\MemOut<15> , 
        \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> , \MemOut<10> , 
        \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> , \MemOut<5> , 
        \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> , \MemOut<0> }), 
        MemToReg, .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }) );
  input \ExecuteOut<15> , \ExecuteOut<14> , \ExecuteOut<13> , \ExecuteOut<12> ,
         \ExecuteOut<11> , \ExecuteOut<10> , \ExecuteOut<9> , \ExecuteOut<8> ,
         \ExecuteOut<7> , \ExecuteOut<6> , \ExecuteOut<5> , \ExecuteOut<4> ,
         \ExecuteOut<3> , \ExecuteOut<2> , \ExecuteOut<1> , \ExecuteOut<0> ,
         \MemOut<15> , \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> ,
         \MemOut<10> , \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> ,
         \MemOut<5> , \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> ,
         \MemOut<0> , MemToReg;
  output \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53;

  MUX2X1 U1 ( .B(n38), .A(n39), .S(n3), .Y(\WriteData<8> ) );
  INVX1 U2 ( .A(n22), .Y(n24) );
  INVX1 U3 ( .A(n22), .Y(n23) );
  INVX1 U4 ( .A(n23), .Y(n1) );
  INVX1 U5 ( .A(n23), .Y(n4) );
  INVX1 U6 ( .A(MemToReg), .Y(n22) );
  INVX1 U7 ( .A(\ExecuteOut<9> ), .Y(n41) );
  INVX1 U8 ( .A(n23), .Y(n3) );
  INVX1 U9 ( .A(n23), .Y(n2) );
  INVX1 U10 ( .A(n24), .Y(n28) );
  MUX2X1 U11 ( .B(n46), .A(n47), .S(n1), .Y(\WriteData<12> ) );
  MUX2X1 U12 ( .B(n44), .A(n45), .S(n2), .Y(\WriteData<11> ) );
  MUX2X1 U13 ( .B(n40), .A(n41), .S(n3), .Y(\WriteData<9> ) );
  MUX2X1 U14 ( .B(n42), .A(n43), .S(n2), .Y(\WriteData<10> ) );
  MUX2X1 U15 ( .B(n52), .A(n53), .S(n35), .Y(\WriteData<15> ) );
  MUX2X1 U16 ( .B(n50), .A(n51), .S(n1), .Y(\WriteData<14> ) );
  MUX2X1 U17 ( .B(n48), .A(n49), .S(n4), .Y(\WriteData<13> ) );
  BUFX2 U18 ( .A(\ExecuteOut<6> ), .Y(n5) );
  AND2X2 U19 ( .A(\ExecuteOut<0> ), .B(n36), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(n7) );
  AND2X2 U21 ( .A(\ExecuteOut<5> ), .B(n36), .Y(n8) );
  INVX1 U22 ( .A(n8), .Y(n9) );
  AND2X2 U23 ( .A(n5), .B(n36), .Y(n10) );
  INVX1 U24 ( .A(n10), .Y(n11) );
  INVX1 U25 ( .A(\MemOut<11> ), .Y(n44) );
  INVX1 U26 ( .A(\MemOut<12> ), .Y(n46) );
  INVX1 U27 ( .A(\MemOut<14> ), .Y(n50) );
  INVX1 U28 ( .A(\MemOut<15> ), .Y(n52) );
  INVX1 U29 ( .A(\MemOut<9> ), .Y(n40) );
  INVX1 U30 ( .A(\MemOut<13> ), .Y(n48) );
  INVX1 U31 ( .A(\MemOut<10> ), .Y(n42) );
  AND2X2 U32 ( .A(\ExecuteOut<1> ), .B(n36), .Y(n12) );
  INVX1 U33 ( .A(n12), .Y(n13) );
  AND2X2 U34 ( .A(\ExecuteOut<2> ), .B(n36), .Y(n14) );
  INVX1 U35 ( .A(n14), .Y(n15) );
  AND2X2 U36 ( .A(\ExecuteOut<3> ), .B(n36), .Y(n16) );
  INVX1 U37 ( .A(n16), .Y(n17) );
  AND2X2 U38 ( .A(\ExecuteOut<4> ), .B(n36), .Y(n18) );
  INVX1 U39 ( .A(n18), .Y(n19) );
  AND2X2 U40 ( .A(\ExecuteOut<7> ), .B(n36), .Y(n20) );
  INVX1 U41 ( .A(n20), .Y(n21) );
  OAI21X1 U42 ( .A(n25), .B(n26), .C(n7), .Y(\WriteData<0> ) );
  INVX1 U43 ( .A(n24), .Y(n26) );
  OAI21X1 U44 ( .A(n34), .B(n35), .C(n11), .Y(\WriteData<6> ) );
  INVX1 U45 ( .A(n24), .Y(n35) );
  OAI21X1 U46 ( .A(n32), .B(n33), .C(n9), .Y(\WriteData<5> ) );
  INVX1 U47 ( .A(n24), .Y(n33) );
  INVX1 U48 ( .A(\MemOut<8> ), .Y(n38) );
  INVX1 U49 ( .A(\MemOut<1> ), .Y(n27) );
  INVX1 U50 ( .A(\ExecuteOut<15> ), .Y(n53) );
  INVX1 U51 ( .A(\ExecuteOut<11> ), .Y(n45) );
  INVX1 U52 ( .A(\ExecuteOut<8> ), .Y(n39) );
  INVX1 U53 ( .A(\ExecuteOut<12> ), .Y(n47) );
  INVX1 U54 ( .A(\MemOut<0> ), .Y(n25) );
  INVX1 U55 ( .A(\MemOut<6> ), .Y(n34) );
  INVX1 U56 ( .A(\MemOut<5> ), .Y(n32) );
  INVX1 U57 ( .A(\MemOut<3> ), .Y(n30) );
  INVX1 U58 ( .A(\MemOut<4> ), .Y(n31) );
  INVX1 U59 ( .A(\ExecuteOut<10> ), .Y(n43) );
  INVX1 U60 ( .A(\MemOut<2> ), .Y(n29) );
  INVX1 U61 ( .A(\ExecuteOut<14> ), .Y(n51) );
  INVX1 U62 ( .A(\MemOut<7> ), .Y(n37) );
  INVX1 U63 ( .A(\ExecuteOut<13> ), .Y(n49) );
  INVX2 U64 ( .A(n24), .Y(n36) );
  AOI22X1 U65 ( .A(n13), .B(n28), .C(n13), .D(n27), .Y(\WriteData<1> ) );
  AOI22X1 U66 ( .A(n15), .B(n26), .C(n15), .D(n29), .Y(\WriteData<2> ) );
  AOI22X1 U67 ( .A(n17), .B(n28), .C(n17), .D(n30), .Y(\WriteData<3> ) );
  AOI22X1 U68 ( .A(n19), .B(n26), .C(n19), .D(n31), .Y(\WriteData<4> ) );
  AOI22X1 U69 ( .A(n21), .B(n33), .C(n21), .D(n37), .Y(\WriteData<7> ) );
endmodule


module proc ( err, clk, rst );
  input clk, rst;
  output err;
  wire   n31, \nextPC<15> , \nextPC<14> , \nextPC<13> , \nextPC<12> ,
         \nextPC<11> , \nextPC<10> , \nextPC<9> , \nextPC<8> , \nextPC<7> ,
         \nextPC<6> , \nextPC<5> , \nextPC<4> , \nextPC<3> , \nextPC<2> ,
         \nextPC<1> , \nextPC<0> , halt, exception, rti, \instr<15> ,
         \instr<14> , \instr<13> , \instr<12> , \instr<11> , \instr<10> ,
         \instr<9> , \instr<8> , \instr<7> , \instr<6> , \instr<5> ,
         \instr<4> , \instr<3> , \instr<2> , \instr<1> , \instr<0> ,
         \incPC<15> , \incPC<14> , \incPC<13> , \incPC<12> , \incPC<11> ,
         \incPC<10> , \incPC<9> , \incPC<8> , \incPC<7> , \incPC<6> ,
         \incPC<5> , \incPC<4> , \incPC<3> , \incPC<2> , \incPC<1> ,
         \incPC<0> , \decode_wr_data<15> , \decode_wr_data<14> ,
         \decode_wr_data<13> , \decode_wr_data<12> , \decode_wr_data<11> ,
         \decode_wr_data<10> , \decode_wr_data<9> , \decode_wr_data<8> ,
         \decode_wr_data<7> , \decode_wr_data<6> , \decode_wr_data<5> ,
         \decode_wr_data<4> , \decode_wr_data<3> , \decode_wr_data<2> ,
         \decode_wr_data<1> , \decode_wr_data<0> , \aluop1<15> , \aluop1<14> ,
         \aluop1<13> , \aluop1<12> , \aluop1<11> , \aluop1<10> , \aluop1<9> ,
         \aluop1<8> , \aluop1<7> , \aluop1<6> , \aluop1<5> , \aluop1<4> ,
         \aluop1<3> , \aluop1<2> , \aluop1<1> , \aluop1<0> , \aluop2<15> ,
         \aluop2<14> , \aluop2<13> , \aluop2<12> , \aluop2<11> , \aluop2<10> ,
         \aluop2<9> , \aluop2<8> , \aluop2<7> , \aluop2<6> , \aluop2<5> ,
         \aluop2<4> , \aluop2<3> , \aluop2<2> , \aluop2<1> , \aluop2<0> ,
         alusrc, branch, jump, jumpreg, set, btr, \aluopcode<2> ,
         \aluopcode<1> , \aluopcode<0> , \func<1> , \func<0> , memwrite,
         memread, memtoreg, \imm<15> , \imm<14> , \imm<13> , \imm<12> ,
         \imm<11> , \imm<10> , \imm<9> , \imm<8> , \imm<7> , \imm<6> ,
         \imm<5> , \imm<4> , \imm<3> , \imm<2> , \imm<1> , \imm<0> , invA,
         invB, cin, \exec_out<15> , \exec_out<14> , \exec_out<13> ,
         \exec_out<12> , \exec_out<11> , \exec_out<10> , \exec_out<9> ,
         \exec_out<8> , \exec_out<7> , \exec_out<6> , \exec_out<5> ,
         \exec_out<4> , \exec_out<3> , \exec_out<2> , \exec_out<1> ,
         \exec_out<0> , \mem_read_data<15> , \mem_read_data<14> ,
         \mem_read_data<13> , \mem_read_data<12> , \mem_read_data<11> ,
         \mem_read_data<10> , \mem_read_data<9> , \mem_read_data<8> ,
         \mem_read_data<7> , \mem_read_data<6> , \mem_read_data<5> ,
         \mem_read_data<4> , \mem_read_data<3> , \mem_read_data<2> ,
         \mem_read_data<1> , \mem_read_data<0> , n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30;
  assign err = 1'b0;

  fetch f ( .NextPC({\nextPC<15> , \nextPC<14> , \nextPC<13> , \nextPC<12> , 
        \nextPC<11> , \nextPC<10> , \nextPC<9> , \nextPC<8> , \nextPC<7> , 
        \nextPC<6> , \nextPC<5> , \nextPC<4> , \nextPC<3> , \nextPC<2> , 
        \nextPC<1> , \nextPC<0> }), .clk(clk), .rst(n29), .Halt(halt), .Rti(
        rti), .Exception(exception), .Instr({\instr<15> , \instr<14> , 
        \instr<13> , \instr<12> , \instr<11> , \instr<10> , \instr<9> , 
        \instr<8> , \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , 
        \instr<2> , \instr<1> , \instr<0> }), .IncPC({\incPC<15> , \incPC<14> , 
        \incPC<13> , \incPC<12> , \incPC<11> , \incPC<10> , \incPC<9> , 
        \incPC<8> , \incPC<7> , \incPC<6> , \incPC<5> , \incPC<4> , \incPC<3> , 
        \incPC<2> , \incPC<1> , \incPC<0> }) );
  decode d ( .clk(clk), .rst(n29), .Instr({\instr<15> , \instr<14> , 
        \instr<13> , \instr<12> , \instr<11> , \instr<10> , \instr<9> , 
        \instr<8> , \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , 
        \instr<2> , \instr<1> , \instr<0> }), .WriteData({\decode_wr_data<15> , 
        \decode_wr_data<14> , \decode_wr_data<13> , \decode_wr_data<12> , 
        \decode_wr_data<11> , \decode_wr_data<10> , \decode_wr_data<9> , 
        \decode_wr_data<8> , \decode_wr_data<7> , \decode_wr_data<6> , 
        \decode_wr_data<5> , \decode_wr_data<4> , \decode_wr_data<3> , 
        \decode_wr_data<2> , \decode_wr_data<1> , \decode_wr_data<0> }), 
        .IncPC({\incPC<15> , \incPC<14> , \incPC<13> , \incPC<12> , 
        \incPC<11> , \incPC<10> , \incPC<9> , \incPC<8> , \incPC<7> , 
        \incPC<6> , \incPC<5> , \incPC<4> , \incPC<3> , \incPC<2> , \incPC<1> , 
        \incPC<0> }), .ALUOp1({\aluop1<15> , \aluop1<14> , \aluop1<13> , 
        \aluop1<12> , \aluop1<11> , \aluop1<10> , \aluop1<9> , \aluop1<8> , 
        \aluop1<7> , \aluop1<6> , \aluop1<5> , \aluop1<4> , \aluop1<3> , 
        \aluop1<2> , \aluop1<1> , \aluop1<0> }), .ALUOp2({\aluop2<15> , 
        \aluop2<14> , \aluop2<13> , \aluop2<12> , \aluop2<11> , \aluop2<10> , 
        \aluop2<9> , \aluop2<8> , \aluop2<7> , \aluop2<6> , \aluop2<5> , 
        \aluop2<4> , \aluop2<3> , \aluop2<2> , \aluop2<1> , \aluop2<0> }), 
        .ALUSrc(alusrc), .Immediate({\imm<15> , \imm<14> , \imm<13> , 
        \imm<12> , \imm<11> , \imm<10> , \imm<9> , \imm<8> , \imm<7> , 
        \imm<6> , \imm<5> , \imm<4> , \imm<3> , \imm<2> , \imm<1> , \imm<0> }), 
        .Branch(branch), .Jump(jump), .JumpReg(jumpreg), .Set(set), .Btr(btr), 
        .InvA(invA), .InvB(invB), .Cin(cin), .ALUOpcode({\aluopcode<2> , 
        \aluopcode<1> , \aluopcode<0> }), .Func({\func<1> , \func<0> }), 
        .MemWrite(memwrite), .MemRead(memread), .MemToReg(memtoreg), .Halt(
        halt), .Exception(exception), .Err(n31), .Rti(rti) );
  execute e ( .ALUOp1({\aluop1<15> , \aluop1<14> , \aluop1<13> , \aluop1<12> , 
        \aluop1<11> , \aluop1<10> , \aluop1<9> , \aluop1<8> , \aluop1<7> , 
        \aluop1<6> , \aluop1<5> , \aluop1<4> , \aluop1<3> , \aluop1<2> , 
        \aluop1<1> , \aluop1<0> }), .ALUOp2({\aluop2<15> , \aluop2<14> , 
        \aluop2<13> , \aluop2<12> , \aluop2<11> , \aluop2<10> , \aluop2<9> , 
        \aluop2<8> , \aluop2<7> , \aluop2<6> , \aluop2<5> , \aluop2<4> , 
        \aluop2<3> , \aluop2<2> , \aluop2<1> , \aluop2<0> }), .Opcode({
        \aluopcode<2> , \aluopcode<1> , \aluopcode<0> }), .IncPC({\incPC<15> , 
        \incPC<14> , \incPC<13> , \incPC<12> , \incPC<11> , \incPC<10> , 
        \incPC<9> , \incPC<8> , \incPC<7> , \incPC<6> , \incPC<5> , \incPC<4> , 
        \incPC<3> , \incPC<2> , \incPC<1> , \incPC<0> }), .Jump(jump), 
        .Branch(branch), .JumpReg(jumpreg), .Set(set), .InvA(invA), .InvB(invB), .Cin(cin), .Btr(btr), .Func({\func<1> , \func<0> }), .Imm({\imm<15> , 
        \imm<14> , \imm<13> , \imm<12> , \imm<11> , \imm<10> , \imm<9> , 
        \imm<8> , \imm<7> , \imm<6> , \imm<5> , \imm<4> , \imm<3> , \imm<2> , 
        \imm<1> , \imm<0> }), .ALUSrc(alusrc), .Result({\exec_out<15> , 
        \exec_out<14> , \exec_out<13> , \exec_out<12> , \exec_out<11> , 
        \exec_out<10> , \exec_out<9> , \exec_out<8> , \exec_out<7> , 
        \exec_out<6> , \exec_out<5> , \exec_out<4> , \exec_out<3> , 
        \exec_out<2> , \exec_out<1> , \exec_out<0> }), .NextPC({\nextPC<15> , 
        \nextPC<14> , \nextPC<13> , \nextPC<12> , \nextPC<11> , \nextPC<10> , 
        \nextPC<9> , \nextPC<8> , \nextPC<7> , \nextPC<6> , \nextPC<5> , 
        \nextPC<4> , \nextPC<3> , \nextPC<2> , \nextPC<1> , \nextPC<0> }) );
  memory m ( .MemRead(memread), .MemWrite(memwrite), .halt(halt), .clk(clk), 
        .rst(n29), .Address({\exec_out<15> , \exec_out<14> , \exec_out<13> , 
        \exec_out<12> , \exec_out<11> , \exec_out<10> , \exec_out<9> , 
        \exec_out<8> , \exec_out<7> , \exec_out<6> , \exec_out<5> , 
        \exec_out<4> , \exec_out<3> , \exec_out<2> , \exec_out<1> , 
        \exec_out<0> }), .WriteData({\aluop2<15> , \aluop2<14> , \aluop2<13> , 
        \aluop2<12> , \aluop2<11> , n7, n9, n8, n22, n2, n4, n3, n13, n19, n1, 
        n5}), .ReadData({\mem_read_data<15> , \mem_read_data<14> , 
        \mem_read_data<13> , \mem_read_data<12> , \mem_read_data<11> , 
        \mem_read_data<10> , \mem_read_data<9> , \mem_read_data<8> , 
        \mem_read_data<7> , \mem_read_data<6> , \mem_read_data<5> , 
        \mem_read_data<4> , \mem_read_data<3> , \mem_read_data<2> , 
        \mem_read_data<1> , \mem_read_data<0> }) );
  writeback w ( .ExecuteOut({n18, n16, n28, n15, \exec_out<11> , n12, n27, n25, 
        n24, \exec_out<6> , n23, n14, n11, \exec_out<2> , \exec_out<1> , n6}), 
        .MemOut({\mem_read_data<15> , \mem_read_data<14> , \mem_read_data<13> , 
        \mem_read_data<12> , \mem_read_data<11> , \mem_read_data<10> , 
        \mem_read_data<9> , \mem_read_data<8> , \mem_read_data<7> , 
        \mem_read_data<6> , \mem_read_data<5> , \mem_read_data<4> , 
        \mem_read_data<3> , \mem_read_data<2> , \mem_read_data<1> , 
        \mem_read_data<0> }), .MemToReg(memtoreg), .WriteData({
        \decode_wr_data<15> , \decode_wr_data<14> , \decode_wr_data<13> , 
        \decode_wr_data<12> , \decode_wr_data<11> , \decode_wr_data<10> , 
        \decode_wr_data<9> , \decode_wr_data<8> , \decode_wr_data<7> , 
        \decode_wr_data<6> , \decode_wr_data<5> , \decode_wr_data<4> , 
        \decode_wr_data<3> , \decode_wr_data<2> , \decode_wr_data<1> , 
        \decode_wr_data<0> }) );
  INVX1 U1 ( .A(n30), .Y(n29) );
  INVX1 U2 ( .A(rst), .Y(n30) );
  BUFX2 U3 ( .A(\aluop2<1> ), .Y(n1) );
  BUFX2 U4 ( .A(\aluop2<6> ), .Y(n2) );
  BUFX2 U5 ( .A(\aluop2<4> ), .Y(n3) );
  BUFX2 U6 ( .A(\aluop2<5> ), .Y(n4) );
  BUFX2 U7 ( .A(\aluop2<0> ), .Y(n5) );
  BUFX2 U8 ( .A(\exec_out<0> ), .Y(n6) );
  BUFX2 U9 ( .A(\aluop2<10> ), .Y(n7) );
  BUFX2 U10 ( .A(\aluop2<8> ), .Y(n8) );
  BUFX2 U11 ( .A(\aluop2<9> ), .Y(n9) );
  INVX1 U12 ( .A(\exec_out<3> ), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(n11) );
  BUFX2 U14 ( .A(\exec_out<10> ), .Y(n12) );
  BUFX2 U15 ( .A(\aluop2<3> ), .Y(n13) );
  BUFX2 U16 ( .A(\exec_out<4> ), .Y(n14) );
  BUFX2 U17 ( .A(\exec_out<12> ), .Y(n15) );
  BUFX2 U18 ( .A(\exec_out<14> ), .Y(n16) );
  INVX1 U19 ( .A(\exec_out<15> ), .Y(n17) );
  INVX1 U20 ( .A(n17), .Y(n18) );
  BUFX2 U21 ( .A(\aluop2<2> ), .Y(n19) );
  INVX1 U23 ( .A(\aluop2<7> ), .Y(n21) );
  INVX2 U24 ( .A(n21), .Y(n22) );
  BUFX2 U25 ( .A(\exec_out<5> ), .Y(n23) );
  BUFX2 U26 ( .A(\exec_out<7> ), .Y(n24) );
  BUFX2 U27 ( .A(\exec_out<8> ), .Y(n25) );
  INVX1 U28 ( .A(\exec_out<9> ), .Y(n26) );
  INVX1 U29 ( .A(n26), .Y(n27) );
  BUFX2 U30 ( .A(\exec_out<13> ), .Y(n28) );
endmodule

