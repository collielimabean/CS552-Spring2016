
module fulladder1_15 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3, n4, n5;

  INVX1 U1 ( .A(Cin), .Y(n5) );
  XOR2X1 U2 ( .A(n4), .B(A), .Y(P) );
  BUFX2 U3 ( .A(P), .Y(n2) );
  INVX1 U4 ( .A(B), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  AND2X2 U6 ( .A(B), .B(A), .Y(G) );
  XNOR2X1 U7 ( .A(n2), .B(n5), .Y(S) );
endmodule


module fulladder1_14 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n4;

  BUFX2 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(A), .Y(n2) );
  XNOR2X1 U3 ( .A(n2), .B(B), .Y(P) );
  BUFX2 U4 ( .A(P), .Y(n4) );
  AND2X2 U5 ( .A(n1), .B(A), .Y(G) );
  XOR2X1 U6 ( .A(Cin), .B(n4), .Y(S) );
endmodule


module fulladder1_13 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  BUFX2 U1 ( .A(B), .Y(n1) );
  AND2X2 U2 ( .A(B), .B(A), .Y(G) );
  XOR2X1 U3 ( .A(B), .B(A), .Y(P) );
  FAX1 U4 ( .A(A), .B(n1), .C(Cin), .YC(), .YS(S) );
endmodule


module fulladder1_12 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(A), .Y(n1) );
  XNOR2X1 U2 ( .A(B), .B(n1), .Y(P) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(B), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  BUFX2 U6 ( .A(n4), .Y(n5) );
  AND2X2 U7 ( .A(n2), .B(n4), .Y(G) );
  XOR2X1 U8 ( .A(n2), .B(n5), .Y(n6) );
  XOR2X1 U9 ( .A(Cin), .B(n6), .Y(S) );
endmodule


module fulladder1_11 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  BUFX2 U1 ( .A(P), .Y(n1) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module fulladder1_10 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  BUFX2 U2 ( .A(P), .Y(n2) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module fulladder1_9 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3, n4;

  BUFX2 U1 ( .A(P), .Y(n1) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  INVX1 U3 ( .A(A), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  AND2X2 U5 ( .A(n4), .B(B), .Y(G) );
  XOR2X1 U6 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module fulladder1_8 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  XOR2X1 U1 ( .A(B), .B(A), .Y(P) );
  BUFX2 U2 ( .A(B), .Y(n1) );
  BUFX2 U3 ( .A(P), .Y(n2) );
  AND2X2 U4 ( .A(A), .B(n1), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module fulladder1_7 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3;

  INVX1 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U3 ( .A(B), .B(A), .Y(G) );
  XNOR2X1 U4 ( .A(n2), .B(A), .Y(n3) );
  INVX2 U5 ( .A(n3), .Y(P) );
  XOR2X1 U6 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_6 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n6, n7;

  XNOR2X1 U1 ( .A(n3), .B(n6), .Y(n1) );
  INVX1 U2 ( .A(n7), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  INVX2 U4 ( .A(A), .Y(n7) );
  XNOR2X1 U5 ( .A(n4), .B(n1), .Y(S) );
  INVX1 U6 ( .A(Cin), .Y(n4) );
  INVX1 U7 ( .A(B), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  XNOR2X1 U9 ( .A(n7), .B(B), .Y(P) );
  AND2X2 U10 ( .A(B), .B(A), .Y(G) );
endmodule


module fulladder1_5 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n3;

  BUFX2 U1 ( .A(P), .Y(n1) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  BUFX2 U3 ( .A(Cin), .Y(n3) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(n3), .B(n1), .Y(S) );
endmodule


module fulladder1_4 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3, n4;

  INVX1 U1 ( .A(P), .Y(n3) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  BUFX2 U3 ( .A(Cin), .Y(n2) );
  XNOR2X1 U4 ( .A(n2), .B(n3), .Y(S) );
  BUFX2 U5 ( .A(B), .Y(n4) );
  AND2X2 U6 ( .A(A), .B(n4), .Y(G) );
endmodule


module fulladder1_3 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10;

  INVX1 U1 ( .A(Cin), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U3 ( .A(n8), .B(n6), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(S) );
  AND2X2 U5 ( .A(n2), .B(n10), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  AND2X2 U7 ( .A(n9), .B(P), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(n8) );
  XNOR2X1 U9 ( .A(A), .B(B), .Y(n10) );
  INVX1 U10 ( .A(Cin), .Y(n9) );
  AND2X2 U11 ( .A(A), .B(B), .Y(G) );
  INVX2 U12 ( .A(n10), .Y(P) );
endmodule


module fulladder1_2 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3, n4, n6, n7, n8, n9, n10;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  AND2X2 U2 ( .A(n8), .B(n10), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  AND2X2 U4 ( .A(n3), .B(n7), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(S) );
  AND2X2 U6 ( .A(n9), .B(P), .Y(n6) );
  INVX1 U7 ( .A(n6), .Y(n7) );
  BUFX2 U8 ( .A(Cin), .Y(n8) );
  INVX1 U9 ( .A(n8), .Y(n9) );
  INVX1 U10 ( .A(P), .Y(n10) );
  AND2X2 U11 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_1 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  INVX1 U2 ( .A(P), .Y(n2) );
  XNOR2X1 U3 ( .A(Cin), .B(n2), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_0 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  INVX1 U2 ( .A(P), .Y(n3) );
  BUFX2 U3 ( .A(Cin), .Y(n2) );
  XNOR2X1 U4 ( .A(n2), .B(n3), .Y(S) );
  AND2X2 U5 ( .A(A), .B(B), .Y(G) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module mux4to1_16_3 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module mux4to1_16_2 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module mux4to1_16_1 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module mux4to1_16_0 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module demux1to8_0 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_1 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_2 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_3 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_4 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_5 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  NOR3X1 U4 ( .A(n7), .B(n4), .C(n6), .Y(Out7) );
  NOR3X1 U5 ( .A(n7), .B(n5), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n6), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(n5), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n6), .C(n7), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(n5), .C(n7), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n6), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out0) );
  INVX1 U1 ( .A(n6), .Y(n5) );
  INVX1 U2 ( .A(n9), .Y(n8) );
  INVX1 U3 ( .A(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(\S<0> ), .Y(n6) );
  INVX1 U13 ( .A(\S<2> ), .Y(n9) );
  AND2X1 U14 ( .A(In), .B(n9), .Y(n1) );
  INVX1 U15 ( .A(n1), .Y(n2) );
  AND2X1 U16 ( .A(n8), .B(In), .Y(n3) );
  INVX1 U17 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_6 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  NOR3X1 U4 ( .A(n7), .B(n4), .C(n6), .Y(Out7) );
  NOR3X1 U5 ( .A(n7), .B(n5), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n6), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(n5), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n6), .C(n7), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(n5), .C(n7), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n6), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out0) );
  INVX1 U1 ( .A(n6), .Y(n5) );
  INVX1 U2 ( .A(n9), .Y(n8) );
  INVX1 U3 ( .A(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(\S<0> ), .Y(n6) );
  INVX1 U13 ( .A(\S<2> ), .Y(n9) );
  AND2X1 U14 ( .A(In), .B(n9), .Y(n1) );
  INVX1 U15 ( .A(n1), .Y(n2) );
  AND2X1 U16 ( .A(n8), .B(In), .Y(n3) );
  INVX1 U17 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_7 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_8 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_9 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_10 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_11 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_12 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_13 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_14 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_15 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to4_17 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n6;

  INVX2 U1 ( .A(\S<0> ), .Y(n3) );
  INVX1 U2 ( .A(\S<1> ), .Y(n4) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n6) );
  INVX1 U6 ( .A(In), .Y(n5) );
  NOR3X1 U7 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U8 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U9 ( .A(n3), .B(n6), .C(\S<1> ), .Y(Out1) );
  AND2X2 U10 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_18 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4;

  INVX1 U1 ( .A(In), .Y(n4) );
  INVX1 U2 ( .A(\S<1> ), .Y(n2) );
  INVX1 U3 ( .A(\S<0> ), .Y(n1) );
  INVX1 U4 ( .A(In), .Y(n3) );
  NOR3X1 U5 ( .A(n2), .B(n1), .C(n3), .Y(Out3) );
  NOR3X1 U6 ( .A(n2), .B(n3), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U7 ( .A(n1), .B(n4), .C(\S<1> ), .Y(Out1) );
  NOR3X1 U8 ( .A(\S<1> ), .B(\S<0> ), .C(n4), .Y(Out0) );
endmodule


module demux1to4_19 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4;

  INVX1 U1 ( .A(\S<0> ), .Y(n1) );
  INVX1 U2 ( .A(\S<1> ), .Y(n2) );
  INVX1 U3 ( .A(In), .Y(n3) );
  INVX1 U4 ( .A(In), .Y(n4) );
  NOR3X1 U5 ( .A(n2), .B(n1), .C(n3), .Y(Out3) );
  NOR3X1 U6 ( .A(n2), .B(n3), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U7 ( .A(n1), .B(n3), .C(\S<1> ), .Y(Out1) );
  NOR3X1 U8 ( .A(\S<1> ), .B(\S<0> ), .C(n4), .Y(Out0) );
endmodule


module demux1to4_20 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<1> ), .Y(n4) );
  INVX1 U2 ( .A(\S<0> ), .Y(n3) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_21 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  INVX1 U2 ( .A(In), .Y(n9) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X1 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(Out0) );
  INVX8 U10 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_22 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<1> ), .Y(n4) );
  INVX1 U2 ( .A(\S<0> ), .Y(n3) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_23 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<0> ), .Y(n3) );
  INVX1 U2 ( .A(\S<1> ), .Y(n4) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_24 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10;

  INVX1 U1 ( .A(\S<1> ), .Y(n9) );
  OR2X1 U2 ( .A(\S<0> ), .B(n8), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n9), .Y(n8) );
  AND2X1 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n9), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  INVX1 U9 ( .A(In), .Y(n10) );
  INVX1 U10 ( .A(\S<0> ), .Y(n7) );
  AND2X2 U11 ( .A(n2), .B(In), .Y(Out0) );
  NOR3X1 U12 ( .A(n9), .B(n7), .C(n10), .Y(Out3) );
  NOR3X1 U13 ( .A(n7), .B(n10), .C(n8), .Y(Out1) );
endmodule


module demux1to4_25 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  AND2X2 U1 ( .A(n7), .B(In), .Y(n3) );
  OR2X1 U2 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  OR2X2 U5 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out2) );
  AND2X2 U7 ( .A(In), .B(n2), .Y(Out0) );
  INVX1 U8 ( .A(\S<0> ), .Y(n7) );
  INVX1 U9 ( .A(\S<1> ), .Y(n8) );
  INVX1 U10 ( .A(In), .Y(n9) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_26 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4;

  INVX1 U1 ( .A(\S<1> ), .Y(n3) );
  INVX1 U2 ( .A(\S<0> ), .Y(n2) );
  INVX1 U3 ( .A(In), .Y(n1) );
  INVX1 U4 ( .A(In), .Y(n4) );
  NOR3X1 U5 ( .A(n3), .B(n2), .C(n4), .Y(Out3) );
  NOR3X1 U6 ( .A(n3), .B(n4), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U7 ( .A(n2), .B(n4), .C(\S<1> ), .Y(Out1) );
  NOR3X1 U8 ( .A(\S<1> ), .B(\S<0> ), .C(n1), .Y(Out0) );
endmodule


module demux1to4_27 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13;

  OR2X1 U1 ( .A(n6), .B(n12), .Y(n7) );
  INVX1 U2 ( .A(n12), .Y(n11) );
  OR2X2 U3 ( .A(n4), .B(n11), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(Out0) );
  AND2X2 U5 ( .A(n10), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  AND2X1 U7 ( .A(n10), .B(n9), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  INVX1 U9 ( .A(n7), .Y(Out2) );
  BUFX2 U10 ( .A(In), .Y(n9) );
  INVX1 U11 ( .A(\S<0> ), .Y(n10) );
  INVX1 U12 ( .A(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(n9), .Y(n13) );
  NOR3X1 U14 ( .A(n12), .B(n10), .C(n13), .Y(Out3) );
  NOR3X1 U15 ( .A(n10), .B(n13), .C(n11), .Y(Out1) );
endmodule


module demux1to4_28 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<0> ), .Y(n7) );
  INVX1 U2 ( .A(\S<1> ), .Y(n8) );
  OR2X2 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X1 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(Out0) );
  INVX1 U10 ( .A(In), .Y(n9) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_29 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n6, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  INVX1 U2 ( .A(In), .Y(n9) );
  AND2X2 U3 ( .A(n7), .B(In), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  OR2X1 U5 ( .A(n2), .B(n8), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(Out2) );
  INVX2 U7 ( .A(n6), .Y(Out0) );
  OR2X2 U8 ( .A(n2), .B(\S<1> ), .Y(n6) );
  INVX8 U9 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U10 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U11 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_30 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n8, n9, n10;

  OR2X1 U1 ( .A(n5), .B(n9), .Y(n6) );
  INVX1 U2 ( .A(In), .Y(n10) );
  INVX1 U3 ( .A(\S<1> ), .Y(n9) );
  OR2X2 U4 ( .A(n3), .B(\S<1> ), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(Out0) );
  INVX1 U6 ( .A(n4), .Y(n3) );
  AND2X2 U7 ( .A(n8), .B(In), .Y(n4) );
  INVX1 U8 ( .A(n4), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(Out2) );
  INVX8 U10 ( .A(\S<0> ), .Y(n8) );
  NOR3X1 U11 ( .A(n9), .B(n8), .C(n10), .Y(Out3) );
  NOR3X1 U12 ( .A(n8), .B(n10), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_31 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n6, n8, n9, n10, n11;

  OR2X1 U1 ( .A(n3), .B(n10), .Y(n4) );
  INVX1 U2 ( .A(n10), .Y(n9) );
  INVX1 U3 ( .A(In), .Y(n11) );
  INVX1 U4 ( .A(n2), .Y(n1) );
  AND2X2 U5 ( .A(n8), .B(In), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(n3) );
  INVX1 U7 ( .A(n4), .Y(Out2) );
  OR2X2 U8 ( .A(n1), .B(n9), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(Out0) );
  INVX1 U10 ( .A(\S<0> ), .Y(n8) );
  INVX1 U11 ( .A(\S<1> ), .Y(n10) );
  NOR3X1 U12 ( .A(n10), .B(n8), .C(n11), .Y(Out3) );
  NOR3X1 U13 ( .A(n8), .B(n11), .C(n9), .Y(Out1) );
endmodule


module demux1to4_32 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<0> ), .Y(n7) );
  INVX1 U2 ( .A(\S<1> ), .Y(n8) );
  INVX1 U3 ( .A(In), .Y(n9) );
  OR2X1 U4 ( .A(n4), .B(n8), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(Out2) );
  AND2X1 U6 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(n4) );
  OR2X2 U8 ( .A(n4), .B(\S<1> ), .Y(n5) );
  INVX1 U9 ( .A(n5), .Y(Out0) );
  NOR3X1 U10 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U11 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_15 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13, n14;

  INVX1 U1 ( .A(\S<0> ), .Y(n14) );
  OR2X2 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  OR2X1 U4 ( .A(n12), .B(n14), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out3) );
  AND2X1 U6 ( .A(\S<0> ), .B(n13), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(n13), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  BUFX2 U14 ( .A(In), .Y(n13) );
  AND2X2 U15 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_14 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13, n14;

  INVX1 U1 ( .A(\S<0> ), .Y(n14) );
  OR2X2 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  OR2X1 U4 ( .A(n12), .B(n14), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out3) );
  AND2X1 U6 ( .A(\S<0> ), .B(n13), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(n13), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  BUFX2 U14 ( .A(In), .Y(n13) );
  AND2X2 U15 ( .A(n2), .B(In), .Y(Out0) );
endmodule


module demux1to4_13 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15;

  INVX1 U1 ( .A(\S<1> ), .Y(n11) );
  OR2X1 U2 ( .A(n10), .B(n14), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  AND2X1 U4 ( .A(n13), .B(n12), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  OR2X2 U6 ( .A(n4), .B(\S<1> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out1) );
  OR2X1 U8 ( .A(n10), .B(n13), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out2) );
  AND2X1 U10 ( .A(n12), .B(\S<1> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(n10) );
  AND2X2 U12 ( .A(n11), .B(n14), .Y(n15) );
  BUFX2 U13 ( .A(In), .Y(n12) );
  INVX1 U14 ( .A(n14), .Y(n13) );
  INVX1 U15 ( .A(\S<0> ), .Y(n14) );
  AND2X2 U16 ( .A(n15), .B(In), .Y(Out0) );
endmodule


module demux1to4_12 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13, n14, n15;

  INVX1 U1 ( .A(\S<0> ), .Y(n15) );
  INVX1 U2 ( .A(n15), .Y(n14) );
  OR2X2 U3 ( .A(\S<1> ), .B(n14), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  OR2X1 U5 ( .A(n12), .B(n15), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(Out3) );
  AND2X1 U7 ( .A(n14), .B(n13), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  OR2X2 U9 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(Out1) );
  OR2X1 U11 ( .A(n12), .B(n14), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Out2) );
  AND2X1 U13 ( .A(n13), .B(\S<1> ), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(n12) );
  BUFX2 U15 ( .A(In), .Y(n13) );
  AND2X2 U16 ( .A(n2), .B(In), .Y(Out0) );
endmodule


module demux1to4_11 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  AND2X2 U2 ( .A(In), .B(\S<1> ), .Y(n11) );
  AND2X2 U3 ( .A(\S<0> ), .B(In), .Y(n5) );
  OR2X1 U4 ( .A(n12), .B(n13), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(Out3) );
  OR2X1 U6 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(n4) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  OR2X2 U9 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(Out1) );
  OR2X1 U11 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Out2) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_10 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9, n10;

  INVX1 U1 ( .A(\S<0> ), .Y(n9) );
  OR2X1 U2 ( .A(n8), .B(n9), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X1 U4 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  OR2X1 U6 ( .A(n8), .B(\S<0> ), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out2) );
  AND2X2 U8 ( .A(In), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(n8) );
  INVX1 U10 ( .A(In), .Y(n10) );
  NOR3X1 U11 ( .A(n9), .B(\S<1> ), .C(n10), .Y(Out1) );
  AND2X2 U12 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_9 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  AND2X2 U2 ( .A(\S<0> ), .B(In), .Y(n5) );
  AND2X2 U3 ( .A(In), .B(\S<1> ), .Y(n11) );
  OR2X2 U4 ( .A(\S<1> ), .B(\S<0> ), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  OR2X1 U6 ( .A(n12), .B(n13), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(Out3) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  OR2X2 U9 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(Out1) );
  OR2X1 U11 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Out2) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_8 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13;

  AND2X2 U1 ( .A(In), .B(\S<1> ), .Y(n11) );
  AND2X2 U2 ( .A(\S<0> ), .B(In), .Y(n5) );
  OR2X2 U3 ( .A(\S<1> ), .B(\S<0> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  OR2X1 U5 ( .A(n12), .B(n13), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(Out3) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  INVX1 U13 ( .A(\S<0> ), .Y(n13) );
  AND2X2 U14 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_7 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n5, n6, n7, n8, n10, n12, n13, n14;

  INVX1 U1 ( .A(\S<0> ), .Y(n14) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(n1), .B(\S<1> ), .Y(n12) );
  AND2X2 U4 ( .A(\S<0> ), .B(n1), .Y(n6) );
  OR2X1 U5 ( .A(n13), .B(n14), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(Out3) );
  OR2X1 U7 ( .A(\S<1> ), .B(\S<0> ), .Y(n4) );
  INVX1 U8 ( .A(n4), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(n7) );
  OR2X2 U10 ( .A(n7), .B(\S<1> ), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(Out1) );
  OR2X1 U12 ( .A(n13), .B(\S<0> ), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(Out2) );
  INVX1 U14 ( .A(n12), .Y(n13) );
  AND2X2 U15 ( .A(In), .B(n5), .Y(Out0) );
endmodule


module demux1to4_6 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n6, n7, n8, n10, n12, n13, n14;

  INVX1 U1 ( .A(\S<0> ), .Y(n14) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(n1), .B(\S<0> ), .Y(n6) );
  AND2X2 U4 ( .A(n1), .B(\S<1> ), .Y(n12) );
  OR2X2 U5 ( .A(\S<1> ), .B(\S<0> ), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(n3) );
  OR2X1 U7 ( .A(n13), .B(n14), .Y(n4) );
  INVX1 U8 ( .A(n4), .Y(Out3) );
  INVX1 U9 ( .A(n6), .Y(n7) );
  OR2X2 U10 ( .A(n7), .B(\S<1> ), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(Out1) );
  OR2X1 U12 ( .A(n13), .B(\S<0> ), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(Out2) );
  INVX1 U14 ( .A(n12), .Y(n13) );
  AND2X2 U15 ( .A(In), .B(n3), .Y(Out0) );
endmodule


module demux1to4_5 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(\S<0> ), .Y(n4) );
  INVX1 U2 ( .A(\S<1> ), .Y(n5) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  BUFX2 U5 ( .A(In), .Y(n3) );
  INVX2 U6 ( .A(n3), .Y(n6) );
  NOR3X1 U7 ( .A(n5), .B(n4), .C(n6), .Y(Out3) );
  NOR3X1 U8 ( .A(n5), .B(n6), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U9 ( .A(n4), .B(n6), .C(\S<1> ), .Y(Out1) );
  AND2X2 U10 ( .A(n2), .B(In), .Y(Out0) );
endmodule


module demux1to4_4 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<0> ), .Y(n3) );
  INVX1 U2 ( .A(\S<1> ), .Y(n4) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_3 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  INVX1 U2 ( .A(In), .Y(n9) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X1 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(Out0) );
  INVX1 U10 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_2 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  OR2X1 U2 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  AND2X1 U4 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  OR2X2 U6 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out2) );
  INVX1 U8 ( .A(In), .Y(n9) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(Out0) );
  INVX1 U10 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_1 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  OR2X1 U2 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  OR2X1 U4 ( .A(n12), .B(n13), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(Out3) );
  AND2X1 U6 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_0 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13, n15;

  OR2X2 U1 ( .A(n12), .B(n15), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out3) );
  AND2X2 U3 ( .A(n15), .B(In), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  AND2X2 U5 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  OR2X2 U7 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(Out1) );
  OR2X1 U9 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(Out2) );
  AND2X1 U11 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  OR2X2 U13 ( .A(n4), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out0) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
endmodule


module cla4_3 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \C<1> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;

  fulladder1_15 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n79), .G(n75) );
  fulladder1_14 \fa[1]  ( .A(n57), .B(\B<1> ), .Cin(\C<1> ), .S(\S<1> ), .P(
        n80), .G(n76) );
  fulladder1_13 \fa[2]  ( .A(n58), .B(\B<2> ), .Cin(n5), .S(\S<2> ), .P(n81), 
        .G(n77) );
  fulladder1_12 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n73), .S(\S<3> ), .P(
        n82), .G(n78) );
  INVX1 U1 ( .A(n15), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(\B<2> ), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  INVX4 U5 ( .A(n61), .Y(n5) );
  INVX2 U6 ( .A(n74), .Y(n61) );
  XNOR2X1 U7 ( .A(\B<1> ), .B(\A<1> ), .Y(n6) );
  INVX1 U8 ( .A(n51), .Y(n10) );
  BUFX2 U9 ( .A(\B<1> ), .Y(n7) );
  BUFX2 U10 ( .A(n40), .Y(n8) );
  INVX1 U11 ( .A(n6), .Y(n9) );
  XNOR2X1 U12 ( .A(n49), .B(n10), .Y(n15) );
  INVX1 U13 ( .A(\A<3> ), .Y(n12) );
  BUFX2 U14 ( .A(n33), .Y(n11) );
  XNOR2X1 U15 ( .A(\B<3> ), .B(n12), .Y(n16) );
  AND2X2 U16 ( .A(n31), .B(n14), .Y(n13) );
  INVX1 U17 ( .A(n69), .Y(n14) );
  OR2X2 U18 ( .A(n56), .B(n22), .Y(n17) );
  INVX1 U19 ( .A(n17), .Y(PG) );
  AND2X2 U20 ( .A(n16), .B(n82), .Y(n19) );
  INVX1 U21 ( .A(n19), .Y(n20) );
  AND2X2 U22 ( .A(n79), .B(n29), .Y(n21) );
  INVX1 U23 ( .A(n21), .Y(n22) );
  BUFX2 U24 ( .A(n66), .Y(n23) );
  BUFX2 U25 ( .A(n68), .Y(n24) );
  OR2X2 U26 ( .A(n40), .B(n6), .Y(n25) );
  INVX1 U27 ( .A(n25), .Y(n26) );
  AND2X2 U28 ( .A(n30), .B(n34), .Y(n27) );
  INVX1 U29 ( .A(n27), .Y(n28) );
  AND2X2 U30 ( .A(n81), .B(n60), .Y(n29) );
  INVX1 U31 ( .A(n29), .Y(n30) );
  AND2X2 U32 ( .A(n9), .B(n80), .Y(n31) );
  INVX1 U33 ( .A(n31), .Y(n32) );
  INVX1 U34 ( .A(n41), .Y(n33) );
  INVX1 U35 ( .A(n33), .Y(n34) );
  INVX1 U36 ( .A(n11), .Y(n35) );
  BUFX2 U37 ( .A(n35), .Y(n36) );
  INVX1 U38 ( .A(n63), .Y(n37) );
  INVX1 U39 ( .A(n64), .Y(n38) );
  INVX1 U40 ( .A(n38), .Y(n39) );
  BUFX2 U41 ( .A(n62), .Y(n40) );
  NAND3X1 U42 ( .A(n54), .B(n4), .C(n77), .Y(n41) );
  INVX1 U43 ( .A(n37), .Y(n65) );
  INVX1 U44 ( .A(n80), .Y(n42) );
  INVX1 U45 ( .A(n42), .Y(n43) );
  BUFX2 U46 ( .A(\B<3> ), .Y(n44) );
  BUFX2 U47 ( .A(\A<3> ), .Y(n45) );
  INVX1 U48 ( .A(n57), .Y(n46) );
  INVX1 U49 ( .A(n46), .Y(n47) );
  INVX1 U50 ( .A(n29), .Y(n48) );
  INVX1 U51 ( .A(n70), .Y(n63) );
  INVX1 U52 ( .A(\B<0> ), .Y(n49) );
  INVX1 U53 ( .A(n49), .Y(n50) );
  INVX1 U54 ( .A(\A<0> ), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(n52) );
  INVX1 U56 ( .A(n58), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(n54) );
  AND2X2 U58 ( .A(n8), .B(n59), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\C<1> ) );
  INVX1 U60 ( .A(n73), .Y(n71) );
  INVX1 U61 ( .A(n13), .Y(n56) );
  BUFX4 U62 ( .A(\A<1> ), .Y(n57) );
  BUFX4 U63 ( .A(\A<2> ), .Y(n58) );
  NAND3X1 U64 ( .A(n2), .B(Cin), .C(n79), .Y(n59) );
  NAND3X1 U65 ( .A(n52), .B(n50), .C(n75), .Y(n62) );
  NAND3X1 U66 ( .A(n47), .B(n7), .C(n76), .Y(n64) );
  OAI21X1 U67 ( .A(n32), .B(n55), .C(n39), .Y(n74) );
  XOR2X1 U68 ( .A(\B<2> ), .B(n58), .Y(n60) );
  OAI21X1 U69 ( .A(n48), .B(n61), .C(n36), .Y(n73) );
  NAND3X1 U70 ( .A(n45), .B(n44), .C(n78), .Y(n70) );
  AOI21X1 U71 ( .A(n43), .B(n26), .C(n63), .Y(n68) );
  AND2X2 U72 ( .A(n35), .B(n39), .Y(n67) );
  AOI21X1 U73 ( .A(n28), .B(n19), .C(n65), .Y(n66) );
  AOI21X1 U74 ( .A(n24), .B(n67), .C(n23), .Y(GG) );
  NAND3X1 U75 ( .A(n15), .B(n16), .C(n82), .Y(n69) );
  OAI21X1 U76 ( .A(n20), .B(n71), .C(n37), .Y(Cout) );
endmodule


module cla4_2 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88;

  fulladder1_11 \fa[0]  ( .A(n62), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(n85), 
        .G(n81) );
  fulladder1_10 \fa[1]  ( .A(\A<1> ), .B(n63), .Cin(n11), .S(\S<1> ), .P(n86), 
        .G(n82) );
  fulladder1_9 \fa[2]  ( .A(\A<2> ), .B(n5), .Cin(n12), .S(\S<2> ), .P(n87), 
        .G(n83) );
  fulladder1_8 \fa[3]  ( .A(n67), .B(\B<3> ), .Cin(n37), .S(\S<3> ), .P(n88), 
        .G(n84) );
  BUFX2 U1 ( .A(Cin), .Y(n1) );
  AND2X1 U2 ( .A(n2), .B(n44), .Y(n22) );
  AND2X1 U3 ( .A(n56), .B(n57), .Y(n24) );
  INVX1 U4 ( .A(n52), .Y(n2) );
  INVX1 U5 ( .A(n8), .Y(n68) );
  INVX1 U6 ( .A(n9), .Y(n3) );
  INVX1 U7 ( .A(n39), .Y(n9) );
  XOR2X1 U8 ( .A(n6), .B(n55), .Y(n10) );
  INVX2 U9 ( .A(\B<0> ), .Y(n6) );
  INVX1 U10 ( .A(n53), .Y(n4) );
  INVX1 U11 ( .A(n60), .Y(n5) );
  INVX1 U12 ( .A(\B<2> ), .Y(n60) );
  INVX1 U13 ( .A(n6), .Y(n7) );
  NOR3X1 U14 ( .A(n9), .B(n34), .C(n31), .Y(n8) );
  AND2X2 U15 ( .A(n10), .B(n85), .Y(n40) );
  AND2X2 U16 ( .A(n64), .B(\B<1> ), .Y(n41) );
  INVX1 U17 ( .A(n31), .Y(n11) );
  AND2X2 U18 ( .A(n47), .B(n23), .Y(n12) );
  AND2X2 U19 ( .A(n61), .B(\A<1> ), .Y(n13) );
  INVX1 U20 ( .A(n13), .Y(n14) );
  AND2X2 U21 ( .A(n10), .B(n66), .Y(n15) );
  INVX1 U22 ( .A(n15), .Y(n16) );
  OR2X2 U23 ( .A(n28), .B(n16), .Y(n17) );
  AND2X2 U24 ( .A(n27), .B(n25), .Y(n18) );
  INVX1 U25 ( .A(n18), .Y(n19) );
  AND2X2 U26 ( .A(n42), .B(n14), .Y(n20) );
  INVX1 U27 ( .A(n20), .Y(n21) );
  INVX1 U28 ( .A(n22), .Y(n23) );
  INVX1 U29 ( .A(n24), .Y(n25) );
  AND2X2 U30 ( .A(n60), .B(\A<2> ), .Y(n26) );
  INVX1 U31 ( .A(n26), .Y(n27) );
  BUFX2 U32 ( .A(n77), .Y(n28) );
  AND2X2 U33 ( .A(n54), .B(n35), .Y(n29) );
  INVX1 U34 ( .A(n29), .Y(n30) );
  AND2X2 U35 ( .A(n49), .B(n2), .Y(n31) );
  BUFX2 U36 ( .A(n76), .Y(n32) );
  AND2X2 U37 ( .A(n21), .B(n86), .Y(n33) );
  INVX1 U38 ( .A(n33), .Y(n34) );
  BUFX2 U39 ( .A(n71), .Y(n35) );
  AND2X2 U40 ( .A(n45), .B(n68), .Y(n36) );
  INVX1 U41 ( .A(n36), .Y(n37) );
  INVX1 U42 ( .A(n36), .Y(n38) );
  AND2X2 U43 ( .A(n87), .B(n19), .Y(n39) );
  INVX1 U44 ( .A(n41), .Y(n42) );
  OR2X1 U45 ( .A(n53), .B(n48), .Y(n43) );
  INVX1 U46 ( .A(n43), .Y(n44) );
  BUFX2 U47 ( .A(n69), .Y(n45) );
  AND2X1 U48 ( .A(n4), .B(n34), .Y(n46) );
  INVX1 U49 ( .A(n46), .Y(n47) );
  INVX1 U50 ( .A(n70), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n49) );
  BUFX2 U52 ( .A(n78), .Y(n50) );
  INVX1 U53 ( .A(n17), .Y(PG) );
  INVX1 U54 ( .A(n35), .Y(n74) );
  AND2X2 U55 ( .A(n1), .B(n40), .Y(n52) );
  INVX1 U56 ( .A(n72), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(n54) );
  INVX1 U58 ( .A(n62), .Y(n55) );
  INVX1 U59 ( .A(n60), .Y(n56) );
  INVX1 U60 ( .A(\A<2> ), .Y(n57) );
  BUFX2 U61 ( .A(\B<3> ), .Y(n58) );
  BUFX2 U62 ( .A(\A<2> ), .Y(n59) );
  INVX1 U63 ( .A(\B<1> ), .Y(n61) );
  BUFX4 U64 ( .A(\A<0> ), .Y(n62) );
  BUFX2 U65 ( .A(\B<1> ), .Y(n63) );
  INVX1 U66 ( .A(\A<1> ), .Y(n64) );
  INVX1 U67 ( .A(n64), .Y(n65) );
  AND2X2 U68 ( .A(n73), .B(n88), .Y(n66) );
  INVX1 U69 ( .A(n66), .Y(n80) );
  BUFX4 U70 ( .A(\A<3> ), .Y(n67) );
  INVX1 U71 ( .A(n38), .Y(n79) );
  NAND3X1 U72 ( .A(n62), .B(n7), .C(n81), .Y(n70) );
  NAND3X1 U73 ( .A(n65), .B(n63), .C(n82), .Y(n72) );
  NAND3X1 U74 ( .A(n59), .B(n5), .C(n83), .Y(n71) );
  AOI21X1 U75 ( .A(n3), .B(n53), .C(n74), .Y(n69) );
  AOI21X1 U76 ( .A(n48), .B(n33), .C(n30), .Y(n76) );
  XOR2X1 U77 ( .A(\B<3> ), .B(n67), .Y(n73) );
  OAI21X1 U78 ( .A(n74), .B(n39), .C(n66), .Y(n75) );
  NAND3X1 U79 ( .A(n67), .B(n58), .C(n84), .Y(n78) );
  OAI21X1 U80 ( .A(n32), .B(n75), .C(n50), .Y(GG) );
  NAND3X1 U81 ( .A(n85), .B(n39), .C(n33), .Y(n77) );
  OAI21X1 U82 ( .A(n80), .B(n79), .C(n50), .Y(Cout) );
endmodule


module cla4_1 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;

  fulladder1_7 \fa[0]  ( .A(n65), .B(\B<0> ), .Cin(n5), .S(\S<0> ), .P(n97), 
        .G(n93) );
  fulladder1_6 \fa[1]  ( .A(n71), .B(n61), .Cin(n90), .S(\S<1> ), .P(n98), .G(
        n94) );
  fulladder1_5 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n91), .S(\S<2> ), .P(n99), .G(n95) );
  fulladder1_4 \fa[3]  ( .A(n68), .B(\B<3> ), .Cin(n92), .S(\S<3> ), .P(n100), 
        .G(n96) );
  INVX1 U1 ( .A(n51), .Y(n82) );
  XOR2X1 U2 ( .A(n59), .B(n6), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(n4), .Y(n3) );
  INVX1 U5 ( .A(Cin), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(n5) );
  BUFX2 U7 ( .A(\A<0> ), .Y(n6) );
  BUFX2 U8 ( .A(\A<0> ), .Y(n65) );
  BUFX2 U9 ( .A(\B<2> ), .Y(n7) );
  INVX1 U10 ( .A(n58), .Y(n8) );
  XOR2X1 U11 ( .A(\A<2> ), .B(\B<2> ), .Y(n9) );
  INVX1 U12 ( .A(n3), .Y(n75) );
  XOR2X1 U13 ( .A(n61), .B(n71), .Y(n10) );
  INVX1 U14 ( .A(\B<1> ), .Y(n12) );
  INVX1 U15 ( .A(n94), .Y(n13) );
  NOR3X1 U16 ( .A(n66), .B(n12), .C(n13), .Y(n11) );
  BUFX2 U17 ( .A(n35), .Y(n14) );
  BUFX4 U18 ( .A(\B<1> ), .Y(n61) );
  AND2X2 U19 ( .A(n29), .B(n47), .Y(n15) );
  INVX1 U20 ( .A(n15), .Y(GG) );
  OR2X2 U21 ( .A(n30), .B(n32), .Y(n17) );
  INVX1 U22 ( .A(n17), .Y(PG) );
  AND2X2 U23 ( .A(n54), .B(n25), .Y(n19) );
  AND2X2 U24 ( .A(n27), .B(n19), .Y(n20) );
  INVX1 U25 ( .A(n20), .Y(n21) );
  OR2X2 U26 ( .A(n37), .B(n35), .Y(n22) );
  INVX1 U27 ( .A(n22), .Y(n23) );
  BUFX2 U28 ( .A(n72), .Y(n24) );
  BUFX2 U29 ( .A(n79), .Y(n25) );
  AND2X2 U30 ( .A(n23), .B(n63), .Y(n26) );
  INVX1 U31 ( .A(n26), .Y(n27) );
  AND2X2 U32 ( .A(n60), .B(n21), .Y(n28) );
  INVX1 U33 ( .A(n28), .Y(n29) );
  BUFX2 U34 ( .A(n80), .Y(n30) );
  AND2X2 U35 ( .A(n1), .B(n67), .Y(n31) );
  INVX1 U36 ( .A(n31), .Y(n32) );
  OR2X2 U37 ( .A(Cin), .B(n81), .Y(n33) );
  INVX1 U38 ( .A(n33), .Y(n34) );
  BUFX2 U39 ( .A(n78), .Y(n35) );
  AND2X2 U40 ( .A(n10), .B(n98), .Y(n36) );
  INVX1 U41 ( .A(n36), .Y(n37) );
  INVX1 U42 ( .A(n36), .Y(n38) );
  AND2X2 U43 ( .A(n55), .B(n49), .Y(n39) );
  AND2X1 U44 ( .A(n52), .B(n38), .Y(n40) );
  INVX1 U45 ( .A(n40), .Y(n41) );
  BUFX2 U46 ( .A(n83), .Y(n42) );
  BUFX2 U47 ( .A(n89), .Y(n43) );
  AND2X1 U48 ( .A(n52), .B(n55), .Y(n44) );
  INVX1 U49 ( .A(n44), .Y(n45) );
  INVX1 U50 ( .A(n87), .Y(n46) );
  INVX1 U51 ( .A(n46), .Y(n47) );
  INVX1 U52 ( .A(n49), .Y(n48) );
  AND2X2 U53 ( .A(n14), .B(n52), .Y(n49) );
  AND2X1 U54 ( .A(n97), .B(n1), .Y(n50) );
  INVX1 U55 ( .A(n50), .Y(n51) );
  INVX1 U56 ( .A(n11), .Y(n52) );
  INVX1 U57 ( .A(n84), .Y(n53) );
  INVX1 U58 ( .A(n53), .Y(n54) );
  INVX1 U59 ( .A(n53), .Y(n55) );
  INVX1 U60 ( .A(\A<2> ), .Y(n56) );
  INVX1 U61 ( .A(n56), .Y(n57) );
  INVX1 U62 ( .A(\B<0> ), .Y(n58) );
  INVX1 U63 ( .A(n58), .Y(n59) );
  INVX1 U64 ( .A(n88), .Y(n60) );
  INVX1 U65 ( .A(n55), .Y(n85) );
  BUFX2 U66 ( .A(\B<3> ), .Y(n62) );
  AND2X2 U67 ( .A(n99), .B(n9), .Y(n63) );
  INVX1 U68 ( .A(n63), .Y(n77) );
  BUFX2 U69 ( .A(n14), .Y(n64) );
  INVX1 U70 ( .A(n71), .Y(n66) );
  AND2X2 U71 ( .A(n100), .B(n76), .Y(n67) );
  INVX1 U72 ( .A(n67), .Y(n88) );
  BUFX4 U73 ( .A(\A<3> ), .Y(n68) );
  INVX1 U74 ( .A(n75), .Y(n69) );
  INVX1 U75 ( .A(n64), .Y(n81) );
  AND2X2 U76 ( .A(n98), .B(n10), .Y(n70) );
  BUFX4 U77 ( .A(\A<1> ), .Y(n71) );
  NAND3X1 U78 ( .A(n6), .B(n8), .C(n93), .Y(n78) );
  NAND3X1 U79 ( .A(n57), .B(n7), .C(n95), .Y(n84) );
  AOI22X1 U80 ( .A(n55), .B(n77), .C(n39), .D(n51), .Y(n72) );
  OAI21X1 U81 ( .A(n70), .B(n45), .C(n24), .Y(n73) );
  AOI21X1 U82 ( .A(n2), .B(n39), .C(n73), .Y(n92) );
  OAI21X1 U83 ( .A(n82), .B(n48), .C(n41), .Y(n74) );
  AOI21X1 U84 ( .A(n75), .B(n49), .C(n74), .Y(n91) );
  AOI21X1 U85 ( .A(n64), .B(n51), .C(n34), .Y(n90) );
  NAND3X1 U86 ( .A(n68), .B(n62), .C(n96), .Y(n87) );
  XOR2X1 U87 ( .A(\B<3> ), .B(n68), .Y(n76) );
  NAND3X1 U88 ( .A(n11), .B(n9), .C(n99), .Y(n79) );
  NAND3X1 U89 ( .A(n63), .B(n97), .C(n70), .Y(n80) );
  AOI21X1 U90 ( .A(n69), .B(n82), .C(n81), .Y(n83) );
  OAI21X1 U91 ( .A(n42), .B(n38), .C(n52), .Y(n86) );
  AOI21X1 U92 ( .A(n63), .B(n86), .C(n85), .Y(n89) );
  OAI21X1 U93 ( .A(n43), .B(n88), .C(n47), .Y(Cout) );
endmodule


module cla4_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  fulladder1_3 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(n74), .G(n70) );
  fulladder1_2 \fa[1]  ( .A(\A<1> ), .B(n39), .Cin(n68), .S(\S<1> ), .P(n75), 
        .G(n71) );
  fulladder1_1 \fa[2]  ( .A(\A<2> ), .B(n43), .Cin(n3), .S(\S<2> ), .P(n76), 
        .G(n72) );
  fulladder1_0 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n69), .S(\S<3> ), .P(n77), .G(n73) );
  INVX1 U1 ( .A(n45), .Y(n1) );
  INVX1 U2 ( .A(n40), .Y(n39) );
  INVX1 U3 ( .A(n50), .Y(n63) );
  AND2X1 U4 ( .A(n45), .B(n10), .Y(n14) );
  AND2X2 U5 ( .A(n4), .B(n35), .Y(n2) );
  INVX1 U6 ( .A(n11), .Y(n3) );
  INVX1 U7 ( .A(Cin), .Y(n4) );
  OR2X2 U8 ( .A(n13), .B(n23), .Y(n5) );
  INVX1 U9 ( .A(n5), .Y(PG) );
  AND2X2 U10 ( .A(\A<2> ), .B(n47), .Y(n7) );
  AND2X2 U11 ( .A(n75), .B(n51), .Y(n8) );
  OR2X2 U12 ( .A(n57), .B(n36), .Y(n9) );
  INVX1 U13 ( .A(n9), .Y(n10) );
  AND2X2 U14 ( .A(n56), .B(n15), .Y(n11) );
  AND2X2 U15 ( .A(n63), .B(n28), .Y(n12) );
  INVX1 U16 ( .A(n12), .Y(n13) );
  INVX1 U17 ( .A(n14), .Y(n15) );
  AND2X2 U18 ( .A(n76), .B(n48), .Y(n16) );
  INVX1 U19 ( .A(n16), .Y(n17) );
  INVX1 U20 ( .A(n16), .Y(n18) );
  AND2X2 U21 ( .A(n52), .B(n35), .Y(n19) );
  INVX1 U22 ( .A(n19), .Y(n20) );
  AND2X1 U23 ( .A(n28), .B(n66), .Y(n21) );
  INVX1 U24 ( .A(n21), .Y(n22) );
  BUFX2 U25 ( .A(n65), .Y(n23) );
  INVX1 U26 ( .A(n55), .Y(n49) );
  BUFX2 U27 ( .A(n62), .Y(n24) );
  AND2X2 U28 ( .A(n7), .B(n72), .Y(n25) );
  INVX1 U29 ( .A(n25), .Y(n26) );
  BUFX2 U30 ( .A(n67), .Y(n27) );
  AND2X2 U31 ( .A(n77), .B(n61), .Y(n28) );
  INVX1 U32 ( .A(n28), .Y(n29) );
  INVX1 U33 ( .A(n3), .Y(n30) );
  AND2X2 U34 ( .A(n26), .B(n17), .Y(n31) );
  INVX1 U35 ( .A(n31), .Y(n32) );
  INVX1 U36 ( .A(n59), .Y(n33) );
  INVX1 U37 ( .A(n26), .Y(n59) );
  INVX1 U38 ( .A(n58), .Y(n34) );
  INVX1 U39 ( .A(n34), .Y(n35) );
  INVX1 U40 ( .A(n8), .Y(n36) );
  INVX1 U41 ( .A(n8), .Y(n37) );
  INVX1 U42 ( .A(n49), .Y(n38) );
  INVX1 U43 ( .A(n40), .Y(n41) );
  INVX1 U44 ( .A(\B<1> ), .Y(n40) );
  AND2X2 U45 ( .A(n74), .B(n63), .Y(n42) );
  INVX1 U46 ( .A(n42), .Y(n57) );
  INVX1 U47 ( .A(n44), .Y(n43) );
  INVX1 U48 ( .A(\B<2> ), .Y(n44) );
  INVX1 U49 ( .A(n46), .Y(n47) );
  INVX1 U50 ( .A(n4), .Y(n45) );
  INVX1 U51 ( .A(\B<2> ), .Y(n46) );
  INVX1 U52 ( .A(n18), .Y(n64) );
  NAND3X1 U53 ( .A(\A<1> ), .B(n41), .C(n71), .Y(n55) );
  XOR2X1 U54 ( .A(n47), .B(\A<2> ), .Y(n48) );
  OAI21X1 U55 ( .A(n49), .B(n59), .C(n32), .Y(n52) );
  NAND3X1 U56 ( .A(\A<0> ), .B(\B<0> ), .C(n70), .Y(n58) );
  XNOR2X1 U57 ( .A(\A<0> ), .B(\B<0> ), .Y(n50) );
  XOR2X1 U58 ( .A(n41), .B(\A<1> ), .Y(n51) );
  OAI21X1 U59 ( .A(n36), .B(n31), .C(n52), .Y(n53) );
  OAI21X1 U60 ( .A(n20), .B(n42), .C(n53), .Y(n54) );
  AOI21X1 U61 ( .A(n19), .B(n1), .C(n54), .Y(n69) );
  OAI21X1 U62 ( .A(n35), .B(n37), .C(n38), .Y(n60) );
  INVX2 U63 ( .A(n60), .Y(n56) );
  AOI21X1 U64 ( .A(n35), .B(n57), .C(n2), .Y(n68) );
  AOI21X1 U65 ( .A(n64), .B(n60), .C(n59), .Y(n62) );
  XOR2X1 U66 ( .A(\B<3> ), .B(\A<3> ), .Y(n61) );
  NAND3X1 U67 ( .A(\A<3> ), .B(\B<3> ), .C(n73), .Y(n67) );
  OAI21X1 U68 ( .A(n29), .B(n24), .C(n27), .Y(GG) );
  NAND3X1 U69 ( .A(n74), .B(n8), .C(n64), .Y(n65) );
  OAI21X1 U70 ( .A(n18), .B(n30), .C(n33), .Y(n66) );
  NAND2X1 U71 ( .A(n27), .B(n22), .Y(Cout) );
endmodule


module fulladder1_44 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_45 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_46 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_47 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_43 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_42 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_41 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_40 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_39 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_38 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_37 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_36 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_35 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_34 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_33 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_32 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module register16_0 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n35;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n19) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n20) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n21) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n22) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n23) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n24) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n25) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n26) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n27) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n28) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n29) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n30) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n31) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n32) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n33) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n34) );
  dff_15 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_14 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_13 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_12 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_11 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_10 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_9 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_8 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_7 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_6 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_5 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_4 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_3 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_2 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_1 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_0 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n34), .Y(n18) );
  INVX1 U5 ( .A(n33), .Y(n12) );
  INVX1 U6 ( .A(n32), .Y(n13) );
  INVX1 U7 ( .A(n31), .Y(n14) );
  INVX1 U8 ( .A(n30), .Y(n15) );
  INVX1 U9 ( .A(n29), .Y(n16) );
  INVX1 U10 ( .A(n28), .Y(n17) );
  INVX1 U11 ( .A(n27), .Y(n3) );
  INVX1 U12 ( .A(n26), .Y(n4) );
  INVX1 U13 ( .A(n25), .Y(n5) );
  INVX1 U14 ( .A(n24), .Y(n6) );
  INVX1 U15 ( .A(n23), .Y(n7) );
  INVX1 U16 ( .A(n22), .Y(n8) );
  INVX1 U17 ( .A(n21), .Y(n9) );
  INVX1 U34 ( .A(n20), .Y(n10) );
  INVX1 U35 ( .A(n19), .Y(n11) );
endmodule


module register16_1 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_31 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_30 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_29 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_28 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_27 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_26 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_25 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_24 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_23 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_22 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_21 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_20 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_19 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_18 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_17 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_16 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_2 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_47 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_46 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_45 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_44 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_43 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_42 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_41 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_40 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_39 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_38 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_37 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_36 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_35 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_34 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_33 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_32 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_3 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_63 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_62 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_61 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_60 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_59 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_58 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_57 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_56 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_55 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_54 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_53 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_52 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_51 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_50 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_49 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_48 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_4 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_79 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_78 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_77 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_76 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_75 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_74 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_73 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_72 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_71 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_70 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_69 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_68 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_67 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_66 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_65 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_64 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_5 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_95 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_94 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_93 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_92 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_91 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_90 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_89 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_88 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_87 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_86 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_85 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_84 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_83 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_82 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_81 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_80 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_6 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_111 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_110 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_109 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_108 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_107 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_106 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_105 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_104 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_103 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_102 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_101 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_100 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_99 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_98 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_97 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_96 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_7 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_112 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_113 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_114 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_115 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_116 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_117 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_118 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_119 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_120 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_121 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_122 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_123 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_124 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_125 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_126 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_127 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module decoder3to8 ( .In({\In<2> , \In<1> , \In<0> }), .Out({\Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<2> , \In<1> , \In<0> ;
  output \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> ,
         \Out<0> ;
  wire   n1, n2, n3;

  NOR3X1 U4 ( .A(n3), .B(n1), .C(n2), .Y(\Out<7> ) );
  NOR3X1 U5 ( .A(n3), .B(\In<0> ), .C(n2), .Y(\Out<6> ) );
  NOR3X1 U6 ( .A(n3), .B(\In<1> ), .C(n1), .Y(\Out<5> ) );
  NOR3X1 U7 ( .A(n3), .B(\In<1> ), .C(\In<0> ), .Y(\Out<4> ) );
  NOR3X1 U8 ( .A(n2), .B(\In<2> ), .C(n1), .Y(\Out<3> ) );
  NOR3X1 U9 ( .A(n2), .B(\In<2> ), .C(\In<0> ), .Y(\Out<2> ) );
  NOR3X1 U10 ( .A(n1), .B(\In<2> ), .C(\In<1> ), .Y(\Out<1> ) );
  NOR3X1 U11 ( .A(\In<0> ), .B(\In<2> ), .C(\In<1> ), .Y(\Out<0> ) );
  INVX1 U1 ( .A(\In<0> ), .Y(n1) );
  INVX1 U2 ( .A(\In<1> ), .Y(n2) );
  INVX1 U3 ( .A(\In<2> ), .Y(n3) );
endmodule


module mux8to1_16_1 ( .In({\In<127> , \In<126> , \In<125> , \In<124> , 
        \In<123> , \In<122> , \In<121> , \In<120> , \In<119> , \In<118> , 
        \In<117> , \In<116> , \In<115> , \In<114> , \In<113> , \In<112> , 
        \In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , 
        \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , 
        \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , 
        \In<78> , \In<77> , \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , 
        \In<71> , \In<70> , \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , 
        \In<64> , \In<63> , \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , 
        \In<57> , \In<56> , \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , 
        \In<50> , \In<49> , \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , 
        \In<43> , \In<42> , \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , 
        \In<36> , \In<35> , \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , 
        \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , 
        \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , 
        \In<0> }), .Sel({\Sel<2> , \Sel<1> , \Sel<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<127> , \In<126> , \In<125> , \In<124> , \In<123> , \In<122> ,
         \In<121> , \In<120> , \In<119> , \In<118> , \In<117> , \In<116> ,
         \In<115> , \In<114> , \In<113> , \In<112> , \In<111> , \In<110> ,
         \In<109> , \In<108> , \In<107> , \In<106> , \In<105> , \In<104> ,
         \In<103> , \In<102> , \In<101> , \In<100> , \In<99> , \In<98> ,
         \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , \In<92> , \In<91> ,
         \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , \In<85> , \In<84> ,
         \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , \In<78> , \In<77> ,
         \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , \In<71> , \In<70> ,
         \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , \In<64> , \In<63> ,
         \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , \In<57> , \In<56> ,
         \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , \In<50> , \In<49> ,
         \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> ,
         \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> ,
         \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , \In<29> , \In<28> ,
         \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , \In<22> , \In<21> ,
         \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , \In<15> , \In<14> ,
         \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , \In<8> , \In<7> ,
         \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , \In<0> ,
         \Sel<2> , \Sel<1> , \Sel<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \mux0_out<15> , \mux0_out<14> , \mux0_out<13> , \mux0_out<12> ,
         \mux0_out<11> , \mux0_out<10> , \mux0_out<9> , \mux0_out<8> ,
         \mux0_out<7> , \mux0_out<6> , \mux0_out<5> , \mux0_out<4> ,
         \mux0_out<3> , \mux0_out<2> , \mux0_out<1> , \mux0_out<0> ,
         \mux1_out<15> , \mux1_out<14> , \mux1_out<13> , \mux1_out<12> ,
         \mux1_out<11> , \mux1_out<10> , \mux1_out<9> , \mux1_out<8> ,
         \mux1_out<7> , \mux1_out<6> , \mux1_out<5> , \mux1_out<4> ,
         \mux1_out<3> , \mux1_out<2> , \mux1_out<1> , \mux1_out<0> , n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  AOI22X1 U18 ( .A(\mux0_out<9> ), .B(n18), .C(\mux1_out<9> ), .D(n17), .Y(n19) );
  AOI22X1 U19 ( .A(\mux0_out<8> ), .B(n18), .C(\mux1_out<8> ), .D(n17), .Y(n20) );
  AOI22X1 U20 ( .A(\mux0_out<7> ), .B(n18), .C(\mux1_out<7> ), .D(n17), .Y(n21) );
  AOI22X1 U21 ( .A(\mux0_out<6> ), .B(n18), .C(\mux1_out<6> ), .D(n17), .Y(n22) );
  AOI22X1 U22 ( .A(\mux0_out<5> ), .B(n18), .C(\mux1_out<5> ), .D(n17), .Y(n23) );
  AOI22X1 U23 ( .A(\mux0_out<4> ), .B(n18), .C(\mux1_out<4> ), .D(n17), .Y(n24) );
  AOI22X1 U24 ( .A(\mux0_out<3> ), .B(n18), .C(\mux1_out<3> ), .D(n17), .Y(n25) );
  AOI22X1 U25 ( .A(\mux0_out<2> ), .B(n18), .C(\mux1_out<2> ), .D(n17), .Y(n26) );
  AOI22X1 U26 ( .A(\mux0_out<1> ), .B(n18), .C(\mux1_out<1> ), .D(n17), .Y(n27) );
  AOI22X1 U27 ( .A(\mux0_out<15> ), .B(n18), .C(\mux1_out<15> ), .D(n17), .Y(
        n28) );
  AOI22X1 U28 ( .A(\mux0_out<14> ), .B(n18), .C(\mux1_out<14> ), .D(n17), .Y(
        n29) );
  AOI22X1 U29 ( .A(\mux0_out<13> ), .B(n18), .C(\mux1_out<13> ), .D(n17), .Y(
        n30) );
  AOI22X1 U30 ( .A(\mux0_out<12> ), .B(n18), .C(\mux1_out<12> ), .D(n17), .Y(
        n31) );
  AOI22X1 U31 ( .A(\mux0_out<11> ), .B(n18), .C(\mux1_out<11> ), .D(n17), .Y(
        n32) );
  AOI22X1 U32 ( .A(\mux0_out<10> ), .B(n18), .C(\mux1_out<10> ), .D(n17), .Y(
        n33) );
  AOI22X1 U33 ( .A(\mux0_out<0> ), .B(n18), .C(\mux1_out<0> ), .D(n17), .Y(n34) );
  mux4to1_16_3 mux0 ( .InA({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .InB({\In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> }), 
        .InC({\In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> , 
        \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> , 
        \In<34> , \In<33> , \In<32> }), .InD({\In<63> , \In<62> , \In<61> , 
        \In<60> , \In<59> , \In<58> , \In<57> , \In<56> , \In<55> , \In<54> , 
        \In<53> , \In<52> , \In<51> , \In<50> , \In<49> , \In<48> }), .S({
        \Sel<1> , \Sel<0> }), .Out({\mux0_out<15> , \mux0_out<14> , 
        \mux0_out<13> , \mux0_out<12> , \mux0_out<11> , \mux0_out<10> , 
        \mux0_out<9> , \mux0_out<8> , \mux0_out<7> , \mux0_out<6> , 
        \mux0_out<5> , \mux0_out<4> , \mux0_out<3> , \mux0_out<2> , 
        \mux0_out<1> , \mux0_out<0> }) );
  mux4to1_16_2 mux1 ( .InA({\In<79> , \In<78> , \In<77> , \In<76> , \In<75> , 
        \In<74> , \In<73> , \In<72> , \In<71> , \In<70> , \In<69> , \In<68> , 
        \In<67> , \In<66> , \In<65> , \In<64> }), .InB({\In<95> , \In<94> , 
        \In<93> , \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , 
        \In<86> , \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> }), 
        .InC({\In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> }), .InD({\In<127> , \In<126> , 
        \In<125> , \In<124> , \In<123> , \In<122> , \In<121> , \In<120> , 
        \In<119> , \In<118> , \In<117> , \In<116> , \In<115> , \In<114> , 
        \In<113> , \In<112> }), .S({\Sel<1> , \Sel<0> }), .Out({\mux1_out<15> , 
        \mux1_out<14> , \mux1_out<13> , \mux1_out<12> , \mux1_out<11> , 
        \mux1_out<10> , \mux1_out<9> , \mux1_out<8> , \mux1_out<7> , 
        \mux1_out<6> , \mux1_out<5> , \mux1_out<4> , \mux1_out<3> , 
        \mux1_out<2> , \mux1_out<1> , \mux1_out<0> }) );
  INVX1 U1 ( .A(n18), .Y(n17) );
  INVX1 U2 ( .A(\Sel<2> ), .Y(n18) );
  BUFX2 U3 ( .A(n34), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(\Out<0> ) );
  BUFX2 U5 ( .A(n33), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(\Out<10> ) );
  BUFX2 U7 ( .A(n32), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(\Out<11> ) );
  BUFX2 U9 ( .A(n31), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(\Out<12> ) );
  BUFX2 U11 ( .A(n30), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(\Out<13> ) );
  BUFX2 U13 ( .A(n29), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(\Out<14> ) );
  BUFX2 U15 ( .A(n28), .Y(n7) );
  INVX1 U16 ( .A(n7), .Y(\Out<15> ) );
  BUFX2 U17 ( .A(n27), .Y(n8) );
  INVX1 U34 ( .A(n8), .Y(\Out<1> ) );
  BUFX2 U35 ( .A(n26), .Y(n9) );
  INVX1 U36 ( .A(n9), .Y(\Out<2> ) );
  BUFX2 U37 ( .A(n25), .Y(n10) );
  INVX1 U38 ( .A(n10), .Y(\Out<3> ) );
  BUFX2 U39 ( .A(n24), .Y(n11) );
  INVX1 U40 ( .A(n11), .Y(\Out<4> ) );
  BUFX2 U41 ( .A(n23), .Y(n12) );
  INVX1 U42 ( .A(n12), .Y(\Out<5> ) );
  BUFX2 U43 ( .A(n22), .Y(n13) );
  INVX1 U44 ( .A(n13), .Y(\Out<6> ) );
  BUFX2 U45 ( .A(n21), .Y(n14) );
  INVX1 U46 ( .A(n14), .Y(\Out<7> ) );
  BUFX2 U47 ( .A(n20), .Y(n15) );
  INVX1 U48 ( .A(n15), .Y(\Out<8> ) );
  BUFX2 U49 ( .A(n19), .Y(n16) );
  INVX1 U50 ( .A(n16), .Y(\Out<9> ) );
endmodule


module mux8to1_16_0 ( .In({\In<127> , \In<126> , \In<125> , \In<124> , 
        \In<123> , \In<122> , \In<121> , \In<120> , \In<119> , \In<118> , 
        \In<117> , \In<116> , \In<115> , \In<114> , \In<113> , \In<112> , 
        \In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , 
        \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , 
        \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , 
        \In<78> , \In<77> , \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , 
        \In<71> , \In<70> , \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , 
        \In<64> , \In<63> , \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , 
        \In<57> , \In<56> , \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , 
        \In<50> , \In<49> , \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , 
        \In<43> , \In<42> , \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , 
        \In<36> , \In<35> , \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , 
        \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , 
        \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , 
        \In<0> }), .Sel({\Sel<2> , \Sel<1> , \Sel<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<127> , \In<126> , \In<125> , \In<124> , \In<123> , \In<122> ,
         \In<121> , \In<120> , \In<119> , \In<118> , \In<117> , \In<116> ,
         \In<115> , \In<114> , \In<113> , \In<112> , \In<111> , \In<110> ,
         \In<109> , \In<108> , \In<107> , \In<106> , \In<105> , \In<104> ,
         \In<103> , \In<102> , \In<101> , \In<100> , \In<99> , \In<98> ,
         \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , \In<92> , \In<91> ,
         \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , \In<85> , \In<84> ,
         \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , \In<78> , \In<77> ,
         \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , \In<71> , \In<70> ,
         \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , \In<64> , \In<63> ,
         \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , \In<57> , \In<56> ,
         \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , \In<50> , \In<49> ,
         \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> ,
         \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> ,
         \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , \In<29> , \In<28> ,
         \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , \In<22> , \In<21> ,
         \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , \In<15> , \In<14> ,
         \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , \In<8> , \In<7> ,
         \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , \In<0> ,
         \Sel<2> , \Sel<1> , \Sel<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \mux0_out<15> , \mux0_out<14> , \mux0_out<13> , \mux0_out<12> ,
         \mux0_out<11> , \mux0_out<10> , \mux0_out<9> , \mux0_out<8> ,
         \mux0_out<7> , \mux0_out<6> , \mux0_out<5> , \mux0_out<4> ,
         \mux0_out<3> , \mux0_out<2> , \mux0_out<1> , \mux0_out<0> ,
         \mux1_out<15> , \mux1_out<14> , \mux1_out<13> , \mux1_out<12> ,
         \mux1_out<11> , \mux1_out<10> , \mux1_out<9> , \mux1_out<8> ,
         \mux1_out<7> , \mux1_out<6> , \mux1_out<5> , \mux1_out<4> ,
         \mux1_out<3> , \mux1_out<2> , \mux1_out<1> , \mux1_out<0> , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66;

  AOI22X1 U18 ( .A(\mux0_out<9> ), .B(n18), .C(\mux1_out<9> ), .D(n17), .Y(n66) );
  AOI22X1 U19 ( .A(\mux0_out<8> ), .B(n18), .C(\mux1_out<8> ), .D(n17), .Y(n65) );
  AOI22X1 U20 ( .A(\mux0_out<7> ), .B(n18), .C(\mux1_out<7> ), .D(n17), .Y(n64) );
  AOI22X1 U21 ( .A(\mux0_out<6> ), .B(n18), .C(\mux1_out<6> ), .D(n17), .Y(n63) );
  AOI22X1 U22 ( .A(\mux0_out<5> ), .B(n18), .C(\mux1_out<5> ), .D(n17), .Y(n62) );
  AOI22X1 U23 ( .A(\mux0_out<4> ), .B(n18), .C(\mux1_out<4> ), .D(n17), .Y(n61) );
  AOI22X1 U24 ( .A(\mux0_out<3> ), .B(n18), .C(\mux1_out<3> ), .D(n17), .Y(n60) );
  AOI22X1 U25 ( .A(\mux0_out<2> ), .B(n18), .C(\mux1_out<2> ), .D(n17), .Y(n59) );
  AOI22X1 U26 ( .A(\mux0_out<1> ), .B(n18), .C(\mux1_out<1> ), .D(n17), .Y(n58) );
  AOI22X1 U27 ( .A(\mux0_out<15> ), .B(n18), .C(\mux1_out<15> ), .D(n17), .Y(
        n57) );
  AOI22X1 U28 ( .A(\mux0_out<14> ), .B(n18), .C(\mux1_out<14> ), .D(n17), .Y(
        n56) );
  AOI22X1 U29 ( .A(\mux0_out<13> ), .B(n18), .C(\mux1_out<13> ), .D(n17), .Y(
        n55) );
  AOI22X1 U30 ( .A(\mux0_out<12> ), .B(n18), .C(\mux1_out<12> ), .D(n17), .Y(
        n54) );
  AOI22X1 U31 ( .A(\mux0_out<11> ), .B(n18), .C(\mux1_out<11> ), .D(n17), .Y(
        n53) );
  AOI22X1 U32 ( .A(\mux0_out<10> ), .B(n18), .C(\mux1_out<10> ), .D(n17), .Y(
        n52) );
  AOI22X1 U33 ( .A(\mux0_out<0> ), .B(n18), .C(\mux1_out<0> ), .D(n17), .Y(n51) );
  mux4to1_16_1 mux0 ( .InA({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .InB({\In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> }), 
        .InC({\In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> , 
        \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> , 
        \In<34> , \In<33> , \In<32> }), .InD({\In<63> , \In<62> , \In<61> , 
        \In<60> , \In<59> , \In<58> , \In<57> , \In<56> , \In<55> , \In<54> , 
        \In<53> , \In<52> , \In<51> , \In<50> , \In<49> , \In<48> }), .S({
        \Sel<1> , \Sel<0> }), .Out({\mux0_out<15> , \mux0_out<14> , 
        \mux0_out<13> , \mux0_out<12> , \mux0_out<11> , \mux0_out<10> , 
        \mux0_out<9> , \mux0_out<8> , \mux0_out<7> , \mux0_out<6> , 
        \mux0_out<5> , \mux0_out<4> , \mux0_out<3> , \mux0_out<2> , 
        \mux0_out<1> , \mux0_out<0> }) );
  mux4to1_16_0 mux1 ( .InA({\In<79> , \In<78> , \In<77> , \In<76> , \In<75> , 
        \In<74> , \In<73> , \In<72> , \In<71> , \In<70> , \In<69> , \In<68> , 
        \In<67> , \In<66> , \In<65> , \In<64> }), .InB({\In<95> , \In<94> , 
        \In<93> , \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , 
        \In<86> , \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> }), 
        .InC({\In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> }), .InD({\In<127> , \In<126> , 
        \In<125> , \In<124> , \In<123> , \In<122> , \In<121> , \In<120> , 
        \In<119> , \In<118> , \In<117> , \In<116> , \In<115> , \In<114> , 
        \In<113> , \In<112> }), .S({\Sel<1> , \Sel<0> }), .Out({\mux1_out<15> , 
        \mux1_out<14> , \mux1_out<13> , \mux1_out<12> , \mux1_out<11> , 
        \mux1_out<10> , \mux1_out<9> , \mux1_out<8> , \mux1_out<7> , 
        \mux1_out<6> , \mux1_out<5> , \mux1_out<4> , \mux1_out<3> , 
        \mux1_out<2> , \mux1_out<1> , \mux1_out<0> }) );
  INVX1 U1 ( .A(n18), .Y(n17) );
  INVX1 U2 ( .A(\Sel<2> ), .Y(n18) );
  BUFX2 U3 ( .A(n51), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(\Out<0> ) );
  BUFX2 U5 ( .A(n52), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(\Out<10> ) );
  BUFX2 U7 ( .A(n53), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(\Out<11> ) );
  BUFX2 U9 ( .A(n54), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(\Out<12> ) );
  BUFX2 U11 ( .A(n55), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(\Out<13> ) );
  BUFX2 U13 ( .A(n56), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(\Out<14> ) );
  BUFX2 U15 ( .A(n57), .Y(n7) );
  INVX1 U16 ( .A(n7), .Y(\Out<15> ) );
  BUFX2 U17 ( .A(n58), .Y(n8) );
  INVX1 U34 ( .A(n8), .Y(\Out<1> ) );
  BUFX2 U35 ( .A(n59), .Y(n9) );
  INVX1 U36 ( .A(n9), .Y(\Out<2> ) );
  BUFX2 U37 ( .A(n60), .Y(n10) );
  INVX1 U38 ( .A(n10), .Y(\Out<3> ) );
  BUFX2 U39 ( .A(n61), .Y(n11) );
  INVX1 U40 ( .A(n11), .Y(\Out<4> ) );
  BUFX2 U41 ( .A(n62), .Y(n12) );
  INVX1 U42 ( .A(n12), .Y(\Out<5> ) );
  BUFX2 U43 ( .A(n63), .Y(n13) );
  INVX1 U44 ( .A(n13), .Y(\Out<6> ) );
  BUFX2 U45 ( .A(n64), .Y(n14) );
  INVX1 U46 ( .A(n14), .Y(\Out<7> ) );
  BUFX2 U47 ( .A(n65), .Y(n15) );
  INVX1 U48 ( .A(n15), .Y(\Out<8> ) );
  BUFX2 U49 ( .A(n66), .Y(n16) );
  INVX1 U50 ( .A(n16), .Y(\Out<9> ) );
endmodule


module demux1to8_16 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<2> , \S<1> , \S<0> }), 
    .Out0({\Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , 
        \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , 
        \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({
        \Out1<15> , \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , 
        \Out1<9> , \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , 
        \Out1<3> , \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , 
        \Out2<14> , \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , 
        \Out2<8> , \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , 
        \Out2<2> , \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , 
        \Out3<13> , \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , 
        \Out3<7> , \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , 
        \Out3<1> , \Out3<0> }), .Out4({\Out4<15> , \Out4<14> , \Out4<13> , 
        \Out4<12> , \Out4<11> , \Out4<10> , \Out4<9> , \Out4<8> , \Out4<7> , 
        \Out4<6> , \Out4<5> , \Out4<4> , \Out4<3> , \Out4<2> , \Out4<1> , 
        \Out4<0> }), .Out5({\Out5<15> , \Out5<14> , \Out5<13> , \Out5<12> , 
        \Out5<11> , \Out5<10> , \Out5<9> , \Out5<8> , \Out5<7> , \Out5<6> , 
        \Out5<5> , \Out5<4> , \Out5<3> , \Out5<2> , \Out5<1> , \Out5<0> }), 
    .Out6({\Out6<15> , \Out6<14> , \Out6<13> , \Out6<12> , \Out6<11> , 
        \Out6<10> , \Out6<9> , \Out6<8> , \Out6<7> , \Out6<6> , \Out6<5> , 
        \Out6<4> , \Out6<3> , \Out6<2> , \Out6<1> , \Out6<0> }), .Out7({
        \Out7<15> , \Out7<14> , \Out7<13> , \Out7<12> , \Out7<11> , \Out7<10> , 
        \Out7<9> , \Out7<8> , \Out7<7> , \Out7<6> , \Out7<5> , \Out7<4> , 
        \Out7<3> , \Out7<2> , \Out7<1> , \Out7<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<2> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> , \Out4<15> ,
         \Out4<14> , \Out4<13> , \Out4<12> , \Out4<11> , \Out4<10> , \Out4<9> ,
         \Out4<8> , \Out4<7> , \Out4<6> , \Out4<5> , \Out4<4> , \Out4<3> ,
         \Out4<2> , \Out4<1> , \Out4<0> , \Out5<15> , \Out5<14> , \Out5<13> ,
         \Out5<12> , \Out5<11> , \Out5<10> , \Out5<9> , \Out5<8> , \Out5<7> ,
         \Out5<6> , \Out5<5> , \Out5<4> , \Out5<3> , \Out5<2> , \Out5<1> ,
         \Out5<0> , \Out6<15> , \Out6<14> , \Out6<13> , \Out6<12> , \Out6<11> ,
         \Out6<10> , \Out6<9> , \Out6<8> , \Out6<7> , \Out6<6> , \Out6<5> ,
         \Out6<4> , \Out6<3> , \Out6<2> , \Out6<1> , \Out6<0> , \Out7<15> ,
         \Out7<14> , \Out7<13> , \Out7<12> , \Out7<11> , \Out7<10> , \Out7<9> ,
         \Out7<8> , \Out7<7> , \Out7<6> , \Out7<5> , \Out7<4> , \Out7<3> ,
         \Out7<2> , \Out7<1> , \Out7<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  demux1to8_0 \demux[0]  ( .In(\In<0> ), .S({n8, n3, \S<0> }), .Out0(\Out0<0> ), .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ), .Out4(\Out4<0> ), 
        .Out5(\Out5<0> ), .Out6(\Out6<0> ), .Out7(\Out7<0> ) );
  demux1to8_1 \demux[1]  ( .In(\In<1> ), .S({n9, n6, n4}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ), .Out4(\Out4<1> ), 
        .Out5(\Out5<1> ), .Out6(\Out6<1> ), .Out7(\Out7<1> ) );
  demux1to8_2 \demux[2]  ( .In(\In<2> ), .S({n9, n6, n4}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ), .Out4(\Out4<2> ), 
        .Out5(\Out5<2> ), .Out6(\Out6<2> ), .Out7(\Out7<2> ) );
  demux1to8_3 \demux[3]  ( .In(\In<3> ), .S({n9, n6, n4}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ), .Out4(\Out4<3> ), 
        .Out5(\Out5<3> ), .Out6(\Out6<3> ), .Out7(\Out7<3> ) );
  demux1to8_4 \demux[4]  ( .In(\In<4> ), .S({n9, n6, n4}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ), .Out4(\Out4<4> ), 
        .Out5(\Out5<4> ), .Out6(\Out6<4> ), .Out7(\Out7<4> ) );
  demux1to8_5 \demux[5]  ( .In(\In<5> ), .S({n8, n1, \S<0> }), .Out0(\Out0<5> ), .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ), .Out4(\Out4<5> ), 
        .Out5(\Out5<5> ), .Out6(\Out6<5> ), .Out7(\Out7<5> ) );
  demux1to8_6 \demux[6]  ( .In(\In<6> ), .S({n8, n2, \S<0> }), .Out0(\Out0<6> ), .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ), .Out4(\Out4<6> ), 
        .Out5(\Out5<6> ), .Out6(\Out6<6> ), .Out7(\Out7<6> ) );
  demux1to8_7 \demux[7]  ( .In(\In<7> ), .S({n8, n3, \S<0> }), .Out0(\Out0<7> ), .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ), .Out4(\Out4<7> ), 
        .Out5(\Out5<7> ), .Out6(\Out6<7> ), .Out7(\Out7<7> ) );
  demux1to8_8 \demux[8]  ( .In(\In<8> ), .S({n8, n1, \S<0> }), .Out0(\Out0<8> ), .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ), .Out4(\Out4<8> ), 
        .Out5(\Out5<8> ), .Out6(\Out6<8> ), .Out7(\Out7<8> ) );
  demux1to8_9 \demux[9]  ( .In(\In<9> ), .S({n8, n2, \S<0> }), .Out0(\Out0<9> ), .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ), .Out4(\Out4<9> ), 
        .Out5(\Out5<9> ), .Out6(\Out6<9> ), .Out7(\Out7<9> ) );
  demux1to8_10 \demux[10]  ( .In(\In<10> ), .S({n8, n3, \S<0> }), .Out0(
        \Out0<10> ), .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ), 
        .Out4(\Out4<10> ), .Out5(\Out5<10> ), .Out6(\Out6<10> ), .Out7(
        \Out7<10> ) );
  demux1to8_11 \demux[11]  ( .In(\In<11> ), .S({n8, n1, \S<0> }), .Out0(
        \Out0<11> ), .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ), 
        .Out4(\Out4<11> ), .Out5(\Out5<11> ), .Out6(\Out6<11> ), .Out7(
        \Out7<11> ) );
  demux1to8_12 \demux[12]  ( .In(\In<12> ), .S({n8, n2, \S<0> }), .Out0(
        \Out0<12> ), .Out1(\Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ), 
        .Out4(\Out4<12> ), .Out5(\Out5<12> ), .Out6(\Out6<12> ), .Out7(
        \Out7<12> ) );
  demux1to8_13 \demux[13]  ( .In(\In<13> ), .S({n8, n3, \S<0> }), .Out0(
        \Out0<13> ), .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ), 
        .Out4(\Out4<13> ), .Out5(\Out5<13> ), .Out6(\Out6<13> ), .Out7(
        \Out7<13> ) );
  demux1to8_14 \demux[14]  ( .In(\In<14> ), .S({n8, n1, \S<0> }), .Out0(
        \Out0<14> ), .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ), 
        .Out4(\Out4<14> ), .Out5(\Out5<14> ), .Out6(\Out6<14> ), .Out7(
        \Out7<14> ) );
  demux1to8_15 \demux[15]  ( .In(\In<15> ), .S({n8, n2, \S<0> }), .Out0(
        \Out0<15> ), .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ), 
        .Out4(\Out4<15> ), .Out5(\Out5<15> ), .Out6(\Out6<15> ), .Out7(
        \Out7<15> ) );
  INVX1 U1 ( .A(n7), .Y(n6) );
  INVX1 U2 ( .A(n7), .Y(n3) );
  INVX1 U3 ( .A(n7), .Y(n1) );
  INVX1 U4 ( .A(n7), .Y(n2) );
  INVX1 U5 ( .A(n5), .Y(n4) );
  INVX1 U6 ( .A(\S<2> ), .Y(n10) );
  INVX1 U7 ( .A(n10), .Y(n9) );
  INVX1 U8 ( .A(n10), .Y(n8) );
  INVX1 U9 ( .A(\S<0> ), .Y(n5) );
  INVX1 U10 ( .A(\S<1> ), .Y(n7) );
endmodule


module demux1to2_17 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_18 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_19 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_20 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  AND2X1 U1 ( .A(In), .B(S), .Y(Out1) );
  INVX1 U2 ( .A(S), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_21 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_22 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_23 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_24 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_25 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(S), .Y(n2) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_26 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_27 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_28 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(S), .Y(n2) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_29 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_30 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_31 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_32 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_15 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_14 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_13 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_12 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_11 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_10 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_9 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_8 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_7 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_6 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_5 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  INVX1 U1 ( .A(n1), .Y(n2) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  BUFX2 U4 ( .A(In), .Y(n1) );
endmodule


module demux1to2_4 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_3 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_2 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_1 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_0 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to4_16_1 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<1> , \S<0> }), .Out0({
        \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , 
        \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , 
        \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , 
        \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , 
        \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , 
        \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , \Out2<14> , 
        \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , 
        \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , 
        \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , \Out3<13> , 
        \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , 
        \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , 
        \Out3<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> ;
  wire   n10, n2, n3, n4, n5, n6, n7, n8, n9;

  demux1to4_17 \demux[0]  ( .In(\In<0> ), .S({n5, n2}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ) );
  demux1to4_18 \demux[1]  ( .In(\In<1> ), .S({n7, n4}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ) );
  demux1to4_19 \demux[2]  ( .In(\In<2> ), .S({n7, n4}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ) );
  demux1to4_20 \demux[3]  ( .In(\In<3> ), .S({n5, n2}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ) );
  demux1to4_21 \demux[4]  ( .In(\In<4> ), .S({n6, n3}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ) );
  demux1to4_22 \demux[5]  ( .In(\In<5> ), .S({n5, n2}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ) );
  demux1to4_23 \demux[6]  ( .In(\In<6> ), .S({n5, n2}), .Out0(\Out0<6> ), 
        .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ) );
  demux1to4_24 \demux[7]  ( .In(\In<7> ), .S({n7, n4}), .Out0(\Out0<7> ), 
        .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ) );
  demux1to4_25 \demux[8]  ( .In(\In<8> ), .S({n7, n4}), .Out0(\Out0<8> ), 
        .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ) );
  demux1to4_26 \demux[9]  ( .In(\In<9> ), .S({n6, n3}), .Out0(\Out0<9> ), 
        .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ) );
  demux1to4_27 \demux[10]  ( .In(\In<10> ), .S({n7, n4}), .Out0(n10), .Out1(
        \Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ) );
  demux1to4_28 \demux[11]  ( .In(\In<11> ), .S({n6, n3}), .Out0(\Out0<11> ), 
        .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ) );
  demux1to4_29 \demux[12]  ( .In(\In<12> ), .S({n6, n3}), .Out0(\Out0<12> ), 
        .Out1(\Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ) );
  demux1to4_30 \demux[13]  ( .In(\In<13> ), .S({n6, n3}), .Out0(\Out0<13> ), 
        .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ) );
  demux1to4_31 \demux[14]  ( .In(\In<14> ), .S({n7, n4}), .Out0(\Out0<14> ), 
        .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ) );
  demux1to4_32 \demux[15]  ( .In(\In<15> ), .S({n6, n3}), .Out0(\Out0<15> ), 
        .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ) );
  INVX4 U1 ( .A(\S<0> ), .Y(n8) );
  BUFX2 U2 ( .A(n10), .Y(\Out0<10> ) );
  INVX4 U3 ( .A(\S<1> ), .Y(n9) );
  INVX8 U4 ( .A(n8), .Y(n2) );
  INVX8 U5 ( .A(n8), .Y(n3) );
  INVX8 U6 ( .A(n8), .Y(n4) );
  INVX8 U7 ( .A(n9), .Y(n5) );
  INVX8 U8 ( .A(n9), .Y(n6) );
  INVX8 U9 ( .A(n9), .Y(n7) );
endmodule


module demux1to4_16_0 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<1> , \S<0> }), .Out0({
        \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , 
        \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , 
        \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , 
        \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , 
        \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , 
        \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , \Out2<14> , 
        \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , 
        \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , 
        \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , \Out3<13> , 
        \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , 
        \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , 
        \Out3<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> ;
  wire   n8, n1, n3, n4, n5, n6, n7;

  demux1to4_15 \demux[0]  ( .In(\In<0> ), .S({n6, n4}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ) );
  demux1to4_14 \demux[1]  ( .In(\In<1> ), .S({n6, n4}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ) );
  demux1to4_13 \demux[2]  ( .In(\In<2> ), .S({n6, n3}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ) );
  demux1to4_12 \demux[3]  ( .In(\In<3> ), .S({n6, n4}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ) );
  demux1to4_11 \demux[4]  ( .In(\In<4> ), .S({n6, n3}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ) );
  demux1to4_10 \demux[5]  ( .In(\In<5> ), .S({n6, n3}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ) );
  demux1to4_9 \demux[6]  ( .In(\In<6> ), .S({n6, n3}), .Out0(\Out0<6> ), 
        .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ) );
  demux1to4_8 \demux[7]  ( .In(\In<7> ), .S({n6, n4}), .Out0(\Out0<7> ), 
        .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ) );
  demux1to4_7 \demux[8]  ( .In(\In<8> ), .S({n6, n3}), .Out0(\Out0<8> ), 
        .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ) );
  demux1to4_6 \demux[9]  ( .In(\In<9> ), .S({n6, n4}), .Out0(\Out0<9> ), 
        .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ) );
  demux1to4_5 \demux[10]  ( .In(\In<10> ), .S({n6, n3}), .Out0(\Out0<10> ), 
        .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ) );
  demux1to4_4 \demux[11]  ( .In(\In<11> ), .S({n6, n4}), .Out0(\Out0<11> ), 
        .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ) );
  demux1to4_3 \demux[12]  ( .In(\In<12> ), .S({n6, n3}), .Out0(n8), .Out1(
        \Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ) );
  demux1to4_2 \demux[13]  ( .In(\In<13> ), .S({n6, n3}), .Out0(\Out0<13> ), 
        .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ) );
  demux1to4_1 \demux[14]  ( .In(\In<14> ), .S({n6, n4}), .Out0(\Out0<14> ), 
        .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ) );
  demux1to4_0 \demux[15]  ( .In(\In<15> ), .S({n6, n4}), .Out0(\Out0<15> ), 
        .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ) );
  INVX2 U1 ( .A(\S<0> ), .Y(n5) );
  INVX2 U2 ( .A(n1), .Y(\Out0<12> ) );
  INVX1 U3 ( .A(\S<1> ), .Y(n7) );
  INVX4 U4 ( .A(n5), .Y(n3) );
  INVX1 U5 ( .A(n8), .Y(n1) );
  INVX8 U6 ( .A(n5), .Y(n4) );
  INVX8 U7 ( .A(n7), .Y(n6) );
endmodule


module cla16_0 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  cla4_3 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_2 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n8), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_1 ca2 ( .A({\A<11> , n22, \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n10), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_0 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n3), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  INVX1 U1 ( .A(n17), .Y(n8) );
  AND2X2 U2 ( .A(n16), .B(\P<1> ), .Y(n13) );
  INVX1 U3 ( .A(\G<3> ), .Y(n28) );
  INVX1 U4 ( .A(\P<0> ), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  OR2X2 U6 ( .A(n4), .B(n5), .Y(n3) );
  INVX1 U7 ( .A(n24), .Y(n4) );
  INVX1 U8 ( .A(n23), .Y(n5) );
  INVX1 U9 ( .A(n26), .Y(n6) );
  INVX1 U10 ( .A(n6), .Y(n7) );
  AND2X2 U11 ( .A(n14), .B(n27), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(n10) );
  AND2X2 U13 ( .A(n28), .B(n20), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(Cout) );
  INVX1 U15 ( .A(n13), .Y(n14) );
  AND2X2 U16 ( .A(n21), .B(n7), .Y(n15) );
  INVX1 U17 ( .A(n15), .Y(n16) );
  AND2X2 U18 ( .A(n25), .B(n26), .Y(n17) );
  INVX1 U19 ( .A(n17), .Y(n18) );
  AND2X2 U20 ( .A(\P<3> ), .B(n3), .Y(n19) );
  INVX1 U21 ( .A(n19), .Y(n20) );
  NAND2X1 U22 ( .A(Cin), .B(n2), .Y(n21) );
  INVX1 U23 ( .A(\G<1> ), .Y(n27) );
  BUFX4 U24 ( .A(\A<10> ), .Y(n22) );
  INVX1 U25 ( .A(\G<0> ), .Y(n26) );
  AOI21X1 U26 ( .A(\G<1> ), .B(\P<2> ), .C(\G<2> ), .Y(n24) );
  NAND2X1 U27 ( .A(Cin), .B(\P<0> ), .Y(n25) );
  NAND3X1 U28 ( .A(\P<1> ), .B(\P<2> ), .C(n18), .Y(n23) );
endmodule


module mux4to1_16_4 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n3, n5, n6, n8, n10, n12, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n103, n104, n105, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148;

  NOR3X1 U1 ( .A(n2), .B(n41), .C(n98), .Y(n1) );
  INVX1 U2 ( .A(n123), .Y(n2) );
  AND2X1 U3 ( .A(\InA<6> ), .B(n136), .Y(n41) );
  AND2X2 U4 ( .A(\InB<6> ), .B(n99), .Y(n98) );
  INVX1 U5 ( .A(\InD<10> ), .Y(n128) );
  OR2X1 U6 ( .A(\InA<11> ), .B(n133), .Y(n37) );
  AND2X2 U7 ( .A(\InA<1> ), .B(n136), .Y(n17) );
  AND2X2 U8 ( .A(n136), .B(\InA<8> ), .Y(n27) );
  AND2X2 U9 ( .A(n136), .B(\InA<4> ), .Y(n22) );
  AND2X2 U10 ( .A(n19), .B(n47), .Y(n3) );
  INVX1 U11 ( .A(n3), .Y(\Out<2> ) );
  AND2X2 U12 ( .A(n23), .B(n48), .Y(n5) );
  AND2X2 U13 ( .A(n34), .B(n50), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(\Out<7> ) );
  OR2X2 U15 ( .A(n38), .B(n86), .Y(n8) );
  INVX1 U16 ( .A(n8), .Y(\Out<11> ) );
  AND2X2 U17 ( .A(n78), .B(n12), .Y(n10) );
  INVX1 U18 ( .A(n10), .Y(\Out<3> ) );
  AND2X2 U19 ( .A(n72), .B(n21), .Y(n12) );
  AND2X2 U20 ( .A(n74), .B(n32), .Y(\Out<13> ) );
  OR2X2 U21 ( .A(n104), .B(n46), .Y(\Out<0> ) );
  OR2X2 U22 ( .A(n105), .B(n16), .Y(\Out<1> ) );
  OR2X2 U23 ( .A(n53), .B(n17), .Y(n16) );
  AND2X2 U24 ( .A(\InA<2> ), .B(n136), .Y(n18) );
  INVX1 U25 ( .A(n18), .Y(n19) );
  AND2X2 U26 ( .A(\InA<3> ), .B(n136), .Y(n20) );
  INVX1 U27 ( .A(n20), .Y(n21) );
  INVX1 U28 ( .A(n22), .Y(n23) );
  AND2X2 U29 ( .A(n36), .B(n71), .Y(n24) );
  INVX1 U30 ( .A(n24), .Y(\Out<10> ) );
  OR2X2 U31 ( .A(n40), .B(n88), .Y(n26) );
  INVX1 U32 ( .A(n27), .Y(n28) );
  AND2X1 U33 ( .A(\InB<15> ), .B(n99), .Y(n29) );
  INVX1 U34 ( .A(n29), .Y(n30) );
  AND2X2 U35 ( .A(n141), .B(n142), .Y(n31) );
  INVX1 U36 ( .A(n31), .Y(n32) );
  AND2X2 U37 ( .A(\InA<7> ), .B(n136), .Y(n33) );
  INVX1 U38 ( .A(n33), .Y(n34) );
  AND2X2 U39 ( .A(\InA<10> ), .B(n136), .Y(n35) );
  INVX1 U40 ( .A(n35), .Y(n36) );
  INVX1 U41 ( .A(n37), .Y(n38) );
  OR2X2 U42 ( .A(\InA<12> ), .B(n137), .Y(n39) );
  INVX1 U43 ( .A(n39), .Y(n40) );
  AND2X2 U44 ( .A(\InA<5> ), .B(n136), .Y(n42) );
  INVX1 U45 ( .A(n42), .Y(n43) );
  AND2X1 U46 ( .A(\InD<15> ), .B(n111), .Y(n44) );
  INVX1 U47 ( .A(n44), .Y(n45) );
  OR2X1 U48 ( .A(n52), .B(n51), .Y(n46) );
  AND2X1 U49 ( .A(n76), .B(n67), .Y(n47) );
  AND2X1 U50 ( .A(n80), .B(n68), .Y(n48) );
  AND2X1 U51 ( .A(n84), .B(n70), .Y(n49) );
  AND2X1 U52 ( .A(n82), .B(n69), .Y(n50) );
  AND2X1 U53 ( .A(\InA<0> ), .B(n136), .Y(n51) );
  AND2X1 U54 ( .A(\InB<0> ), .B(n99), .Y(n52) );
  AND2X1 U55 ( .A(\InB<1> ), .B(n99), .Y(n53) );
  AND2X1 U56 ( .A(\InD<9> ), .B(n111), .Y(n54) );
  INVX1 U57 ( .A(n54), .Y(n55) );
  AND2X1 U58 ( .A(\InD<14> ), .B(n111), .Y(n56) );
  INVX1 U59 ( .A(n56), .Y(n57) );
  AND2X1 U60 ( .A(\InB<9> ), .B(n99), .Y(n58) );
  INVX1 U61 ( .A(n58), .Y(n59) );
  AND2X1 U62 ( .A(\InB<14> ), .B(n99), .Y(n60) );
  INVX1 U63 ( .A(n60), .Y(n61) );
  BUFX2 U64 ( .A(n131), .Y(n62) );
  BUFX2 U65 ( .A(n134), .Y(n63) );
  BUFX2 U66 ( .A(n138), .Y(n64) );
  AND2X1 U67 ( .A(\InB<10> ), .B(n99), .Y(n65) );
  INVX1 U68 ( .A(n65), .Y(n66) );
  BUFX2 U69 ( .A(n119), .Y(n67) );
  BUFX2 U70 ( .A(n121), .Y(n68) );
  BUFX2 U71 ( .A(n124), .Y(n69) );
  BUFX2 U72 ( .A(n125), .Y(n70) );
  BUFX2 U73 ( .A(n130), .Y(n71) );
  BUFX2 U74 ( .A(n120), .Y(n72) );
  AND2X1 U75 ( .A(n147), .B(n142), .Y(n73) );
  INVX1 U76 ( .A(n73), .Y(n74) );
  AND2X1 U77 ( .A(\InC<2> ), .B(n113), .Y(n75) );
  INVX1 U78 ( .A(n75), .Y(n76) );
  AND2X1 U79 ( .A(\InB<3> ), .B(n99), .Y(n77) );
  INVX1 U80 ( .A(n77), .Y(n78) );
  AND2X1 U81 ( .A(\InC<4> ), .B(n113), .Y(n79) );
  INVX1 U82 ( .A(n79), .Y(n80) );
  AND2X1 U83 ( .A(\InC<7> ), .B(n113), .Y(n81) );
  INVX1 U84 ( .A(n81), .Y(n82) );
  AND2X1 U85 ( .A(\InC<8> ), .B(n113), .Y(n83) );
  INVX1 U86 ( .A(n83), .Y(n84) );
  OR2X1 U87 ( .A(n133), .B(n136), .Y(n85) );
  INVX1 U88 ( .A(n85), .Y(n86) );
  OR2X1 U89 ( .A(n137), .B(n136), .Y(n87) );
  INVX1 U90 ( .A(n87), .Y(n88) );
  AND2X2 U91 ( .A(n55), .B(n59), .Y(n89) );
  INVX1 U92 ( .A(n89), .Y(n90) );
  AND2X2 U93 ( .A(n57), .B(n61), .Y(n91) );
  INVX1 U94 ( .A(n91), .Y(n92) );
  AND2X2 U95 ( .A(n45), .B(n30), .Y(n93) );
  INVX1 U96 ( .A(n93), .Y(n94) );
  AND2X1 U97 ( .A(\InC<5> ), .B(n113), .Y(n95) );
  INVX1 U98 ( .A(n95), .Y(n96) );
  BUFX2 U99 ( .A(n122), .Y(n97) );
  AND2X1 U100 ( .A(\S<0> ), .B(n116), .Y(n99) );
  INVX1 U101 ( .A(n26), .Y(\Out<12> ) );
  BUFX2 U102 ( .A(n148), .Y(\Out<9> ) );
  OR2X1 U103 ( .A(\S<1> ), .B(\S<0> ), .Y(n147) );
  INVX1 U104 ( .A(n140), .Y(n142) );
  INVX1 U105 ( .A(n103), .Y(\Out<8> ) );
  AND2X2 U106 ( .A(n28), .B(n49), .Y(n103) );
  INVX1 U107 ( .A(n117), .Y(n104) );
  INVX1 U108 ( .A(n118), .Y(n105) );
  INVX1 U109 ( .A(n1), .Y(\Out<6> ) );
  INVX1 U110 ( .A(n5), .Y(\Out<4> ) );
  BUFX2 U111 ( .A(n144), .Y(n108) );
  BUFX2 U112 ( .A(n146), .Y(n109) );
  BUFX2 U113 ( .A(n127), .Y(n110) );
  AND2X1 U114 ( .A(\S<0> ), .B(\S<1> ), .Y(n111) );
  INVX1 U115 ( .A(n111), .Y(n112) );
  AND2X1 U116 ( .A(n115), .B(\S<1> ), .Y(n113) );
  INVX1 U117 ( .A(n113), .Y(n114) );
  INVX1 U118 ( .A(\S<0> ), .Y(n115) );
  INVX1 U119 ( .A(\S<1> ), .Y(n116) );
  INVX1 U120 ( .A(\InA<9> ), .Y(n126) );
  INVX1 U121 ( .A(\InA<13> ), .Y(n141) );
  INVX1 U122 ( .A(\InA<14> ), .Y(n143) );
  INVX1 U123 ( .A(\InA<15> ), .Y(n145) );
  INVX4 U124 ( .A(n147), .Y(n136) );
  AOI22X1 U125 ( .A(\InD<0> ), .B(n111), .C(\InC<0> ), .D(n113), .Y(n117) );
  AOI22X1 U126 ( .A(\InD<1> ), .B(n111), .C(\InC<1> ), .D(n113), .Y(n118) );
  AOI22X1 U127 ( .A(\InD<2> ), .B(n111), .C(\InB<2> ), .D(n99), .Y(n119) );
  AOI22X1 U128 ( .A(\InD<3> ), .B(n111), .C(\InC<3> ), .D(n113), .Y(n120) );
  AOI22X1 U129 ( .A(\InD<4> ), .B(n111), .C(\InB<4> ), .D(n99), .Y(n121) );
  AOI22X1 U130 ( .A(\InB<5> ), .B(n99), .C(\InD<5> ), .D(n111), .Y(n122) );
  NAND3X1 U131 ( .A(n96), .B(n97), .C(n43), .Y(\Out<5> ) );
  AOI22X1 U132 ( .A(\InD<6> ), .B(n111), .C(\InC<6> ), .D(n113), .Y(n123) );
  AOI22X1 U133 ( .A(\InD<7> ), .B(n111), .C(\InB<7> ), .D(n99), .Y(n124) );
  AOI22X1 U134 ( .A(\InD<8> ), .B(n111), .C(\InB<8> ), .D(n99), .Y(n125) );
  AOI21X1 U135 ( .A(\InC<9> ), .B(n113), .C(n90), .Y(n127) );
  AOI22X1 U136 ( .A(n147), .B(n110), .C(n126), .D(n110), .Y(n148) );
  OAI21X1 U137 ( .A(n112), .B(n128), .C(n66), .Y(n129) );
  AOI21X1 U138 ( .A(\InC<10> ), .B(n113), .C(n129), .Y(n130) );
  INVX2 U139 ( .A(\InC<11> ), .Y(n132) );
  AOI22X1 U140 ( .A(\InD<11> ), .B(n111), .C(\InB<11> ), .D(n99), .Y(n131) );
  OAI21X1 U141 ( .A(n114), .B(n132), .C(n62), .Y(n133) );
  INVX2 U142 ( .A(\InC<12> ), .Y(n135) );
  AOI22X1 U143 ( .A(\InD<12> ), .B(n111), .C(\InB<12> ), .D(n99), .Y(n134) );
  OAI21X1 U144 ( .A(n114), .B(n135), .C(n63), .Y(n137) );
  INVX2 U145 ( .A(\InC<13> ), .Y(n139) );
  AOI22X1 U146 ( .A(\InD<13> ), .B(n111), .C(\InB<13> ), .D(n99), .Y(n138) );
  OAI21X1 U147 ( .A(n114), .B(n139), .C(n64), .Y(n140) );
  AOI21X1 U148 ( .A(\InC<14> ), .B(n113), .C(n92), .Y(n144) );
  AOI22X1 U149 ( .A(n147), .B(n108), .C(n108), .D(n143), .Y(\Out<14> ) );
  AOI21X1 U150 ( .A(\InC<15> ), .B(n113), .C(n94), .Y(n146) );
  AOI22X1 U151 ( .A(n147), .B(n109), .C(n109), .D(n145), .Y(\Out<15> ) );
endmodule


module lshifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), Rot_sel, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , Rot_sel;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33,
         n35, n36, n37, n39, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n145, n147, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277;

  AND2X2 U2 ( .A(\Cnt<0> ), .B(\Cnt<1> ), .Y(n7) );
  INVX1 U3 ( .A(\In<4> ), .Y(n248) );
  INVX1 U4 ( .A(\Cnt<2> ), .Y(n209) );
  INVX1 U5 ( .A(\Cnt<3> ), .Y(n203) );
  AND2X1 U6 ( .A(n111), .B(n107), .Y(n27) );
  INVX1 U7 ( .A(\In<0> ), .Y(n212) );
  INVX8 U8 ( .A(n242), .Y(n254) );
  INVX4 U9 ( .A(n7), .Y(n8) );
  INVX1 U10 ( .A(n204), .Y(n1) );
  AND2X2 U11 ( .A(n204), .B(\Cnt<1> ), .Y(n172) );
  OR2X2 U12 ( .A(n78), .B(n3), .Y(\Out<6> ) );
  OR2X2 U13 ( .A(n141), .B(n151), .Y(n3) );
  OR2X2 U14 ( .A(n67), .B(n5), .Y(n4) );
  OR2X2 U15 ( .A(n181), .B(n75), .Y(n5) );
  AND2X2 U16 ( .A(n203), .B(\Cnt<2> ), .Y(n6) );
  AND2X2 U17 ( .A(\Cnt<0> ), .B(n213), .Y(n9) );
  INVX1 U18 ( .A(n9), .Y(n10) );
  AND2X2 U19 ( .A(Rot_sel), .B(n62), .Y(n11) );
  OR2X2 U20 ( .A(n8), .B(n206), .Y(n12) );
  INVX1 U21 ( .A(n12), .Y(n13) );
  AND2X2 U22 ( .A(Rot_sel), .B(n165), .Y(n14) );
  AND2X2 U23 ( .A(n213), .B(n239), .Y(n15) );
  INVX1 U24 ( .A(n15), .Y(n16) );
  AND2X2 U25 ( .A(\In<14> ), .B(n172), .Y(n17) );
  INVX1 U26 ( .A(n17), .Y(n18) );
  AND2X2 U27 ( .A(n109), .B(n104), .Y(n19) );
  INVX1 U28 ( .A(n19), .Y(\Out<0> ) );
  AND2X2 U29 ( .A(\In<0> ), .B(n164), .Y(n21) );
  INVX1 U30 ( .A(n21), .Y(n22) );
  AND2X2 U31 ( .A(\In<15> ), .B(n172), .Y(n23) );
  INVX1 U32 ( .A(n23), .Y(n24) );
  AND2X2 U33 ( .A(n110), .B(n105), .Y(n25) );
  INVX1 U34 ( .A(n25), .Y(\Out<1> ) );
  INVX1 U35 ( .A(n27), .Y(\Out<2> ) );
  OR2X2 U36 ( .A(n8), .B(n245), .Y(n29) );
  INVX1 U37 ( .A(n29), .Y(n30) );
  OR2X2 U38 ( .A(n8), .B(n248), .Y(n31) );
  INVX1 U39 ( .A(n31), .Y(n32) );
  AND2X2 U40 ( .A(n112), .B(n108), .Y(n33) );
  INVX1 U41 ( .A(n33), .Y(\Out<3> ) );
  AND2X2 U42 ( .A(n6), .B(n187), .Y(n35) );
  INVX1 U43 ( .A(n35), .Y(n36) );
  AND2X2 U44 ( .A(n114), .B(n56), .Y(n37) );
  INVX1 U45 ( .A(n37), .Y(\Out<12> ) );
  AND2X2 U46 ( .A(n58), .B(n57), .Y(n39) );
  INVX1 U47 ( .A(n39), .Y(\Out<15> ) );
  BUFX2 U48 ( .A(n264), .Y(n41) );
  BUFX2 U49 ( .A(n261), .Y(n42) );
  BUFX2 U50 ( .A(n263), .Y(n43) );
  BUFX2 U51 ( .A(n219), .Y(n44) );
  BUFX2 U52 ( .A(n224), .Y(n45) );
  BUFX2 U53 ( .A(n231), .Y(n46) );
  BUFX2 U54 ( .A(n234), .Y(n47) );
  BUFX2 U55 ( .A(n237), .Y(n48) );
  BUFX2 U56 ( .A(n246), .Y(n49) );
  BUFX2 U57 ( .A(n252), .Y(n50) );
  BUFX2 U58 ( .A(n255), .Y(n51) );
  AND2X2 U59 ( .A(Rot_sel), .B(n215), .Y(n52) );
  INVX1 U60 ( .A(n52), .Y(n53) );
  AND2X2 U61 ( .A(Rot_sel), .B(n227), .Y(n54) );
  INVX1 U62 ( .A(n54), .Y(n55) );
  BUFX2 U63 ( .A(n270), .Y(n56) );
  BUFX2 U64 ( .A(n276), .Y(n57) );
  BUFX2 U65 ( .A(n277), .Y(n58) );
  BUFX2 U66 ( .A(n259), .Y(n59) );
  OR2X2 U67 ( .A(n200), .B(n201), .Y(n60) );
  INVX1 U68 ( .A(n60), .Y(n61) );
  AND2X2 U69 ( .A(\Cnt<3> ), .B(\Cnt<2> ), .Y(n62) );
  INVX1 U70 ( .A(n247), .Y(n63) );
  INVX1 U71 ( .A(n63), .Y(n64) );
  INVX1 U72 ( .A(n250), .Y(n65) );
  INVX1 U73 ( .A(n65), .Y(n66) );
  AND2X2 U74 ( .A(\In<6> ), .B(n172), .Y(n67) );
  OR2X1 U75 ( .A(n8), .B(n218), .Y(n68) );
  INVX1 U76 ( .A(n68), .Y(n69) );
  OR2X1 U77 ( .A(n8), .B(n241), .Y(n70) );
  INVX1 U78 ( .A(n70), .Y(n71) );
  AND2X2 U79 ( .A(n165), .B(n273), .Y(n72) );
  INVX1 U80 ( .A(n72), .Y(n73) );
  AND2X2 U81 ( .A(n116), .B(n22), .Y(n74) );
  AND2X2 U82 ( .A(\In<5> ), .B(n7), .Y(n75) );
  AND2X2 U83 ( .A(n6), .B(n174), .Y(n76) );
  INVX1 U84 ( .A(n76), .Y(n77) );
  AND2X1 U85 ( .A(n11), .B(n185), .Y(n78) );
  BUFX2 U86 ( .A(n208), .Y(n79) );
  INVX1 U87 ( .A(n220), .Y(n80) );
  INVX1 U88 ( .A(n80), .Y(n81) );
  BUFX2 U89 ( .A(n222), .Y(n82) );
  INVX1 U90 ( .A(n225), .Y(n83) );
  INVX1 U91 ( .A(n83), .Y(n84) );
  BUFX2 U92 ( .A(n232), .Y(n85) );
  BUFX2 U93 ( .A(n235), .Y(n86) );
  BUFX2 U94 ( .A(n238), .Y(n87) );
  INVX1 U95 ( .A(n253), .Y(n88) );
  INVX1 U96 ( .A(n88), .Y(n89) );
  INVX1 U97 ( .A(n256), .Y(n90) );
  INVX1 U98 ( .A(n90), .Y(n91) );
  INVX1 U99 ( .A(n262), .Y(n92) );
  INVX1 U100 ( .A(n92), .Y(n93) );
  BUFX2 U101 ( .A(n268), .Y(n94) );
  BUFX2 U102 ( .A(n267), .Y(n95) );
  INVX1 U103 ( .A(n207), .Y(n96) );
  INVX1 U104 ( .A(n96), .Y(n97) );
  INVX1 U105 ( .A(n221), .Y(n98) );
  INVX1 U106 ( .A(n98), .Y(n99) );
  INVX1 U107 ( .A(n249), .Y(n100) );
  INVX1 U108 ( .A(n100), .Y(n101) );
  INVX1 U109 ( .A(n240), .Y(n102) );
  INVX1 U110 ( .A(n102), .Y(n103) );
  BUFX2 U111 ( .A(n216), .Y(n104) );
  BUFX2 U112 ( .A(n228), .Y(n105) );
  INVX1 U113 ( .A(n243), .Y(n106) );
  INVX1 U114 ( .A(n106), .Y(n107) );
  BUFX2 U115 ( .A(n257), .Y(n108) );
  BUFX2 U116 ( .A(n217), .Y(n109) );
  BUFX2 U117 ( .A(n229), .Y(n110) );
  BUFX2 U118 ( .A(n244), .Y(n111) );
  BUFX2 U119 ( .A(n258), .Y(n112) );
  INVX1 U120 ( .A(n271), .Y(n113) );
  INVX1 U121 ( .A(n113), .Y(n114) );
  AND2X2 U122 ( .A(\In<1> ), .B(n254), .Y(n115) );
  INVX1 U123 ( .A(n115), .Y(n116) );
  OR2X1 U124 ( .A(n8), .B(n223), .Y(n117) );
  INVX1 U125 ( .A(n117), .Y(n118) );
  OR2X2 U126 ( .A(n8), .B(n230), .Y(n119) );
  INVX1 U127 ( .A(n119), .Y(n120) );
  OR2X1 U128 ( .A(n8), .B(n233), .Y(n121) );
  INVX1 U129 ( .A(n121), .Y(n122) );
  OR2X1 U130 ( .A(n8), .B(n236), .Y(n123) );
  INVX1 U131 ( .A(n123), .Y(n124) );
  OR2X1 U132 ( .A(n8), .B(n251), .Y(n125) );
  INVX1 U133 ( .A(n125), .Y(n126) );
  OR2X1 U134 ( .A(n8), .B(n212), .Y(n127) );
  INVX1 U135 ( .A(n127), .Y(n128) );
  AND2X2 U136 ( .A(\In<10> ), .B(n172), .Y(n129) );
  INVX1 U137 ( .A(n129), .Y(n130) );
  AND2X2 U138 ( .A(n11), .B(n4), .Y(n131) );
  INVX1 U139 ( .A(n131), .Y(n132) );
  AND2X2 U140 ( .A(n11), .B(n183), .Y(n133) );
  INVX1 U141 ( .A(n133), .Y(n134) );
  AND2X2 U142 ( .A(n165), .B(n174), .Y(n135) );
  INVX1 U143 ( .A(n135), .Y(n136) );
  AND2X2 U144 ( .A(n62), .B(n174), .Y(n137) );
  INVX1 U145 ( .A(n137), .Y(n138) );
  AND2X1 U146 ( .A(n62), .B(n273), .Y(n139) );
  INVX1 U147 ( .A(n139), .Y(n140) );
  INVX1 U148 ( .A(n260), .Y(n141) );
  AND2X1 U149 ( .A(Rot_sel), .B(n6), .Y(n142) );
  AND2X2 U150 ( .A(n93), .B(n42), .Y(n143) );
  INVX1 U151 ( .A(n143), .Y(\Out<7> ) );
  AND2X2 U152 ( .A(n41), .B(n43), .Y(n145) );
  INVX1 U153 ( .A(n145), .Y(\Out<8> ) );
  AND2X2 U154 ( .A(n94), .B(n95), .Y(n147) );
  INVX1 U155 ( .A(n147), .Y(\Out<11> ) );
  AND2X1 U156 ( .A(\In<15> ), .B(Rot_sel), .Y(n149) );
  INVX1 U157 ( .A(n149), .Y(n150) );
  AND2X1 U158 ( .A(n6), .B(n273), .Y(n151) );
  AND2X2 U159 ( .A(n11), .B(n176), .Y(n152) );
  INVX1 U160 ( .A(n152), .Y(n153) );
  AND2X1 U161 ( .A(n11), .B(n178), .Y(n154) );
  INVX1 U162 ( .A(n154), .Y(n155) );
  AND2X2 U163 ( .A(n165), .B(n189), .Y(n156) );
  INVX1 U164 ( .A(n156), .Y(n157) );
  AND2X1 U165 ( .A(n165), .B(n191), .Y(n158) );
  INVX1 U166 ( .A(n158), .Y(n159) );
  BUFX2 U167 ( .A(n265), .Y(n160) );
  BUFX2 U168 ( .A(n266), .Y(n161) );
  BUFX2 U169 ( .A(n272), .Y(n162) );
  BUFX2 U170 ( .A(n274), .Y(n163) );
  INVX4 U171 ( .A(n10), .Y(n164) );
  AND2X1 U172 ( .A(\Cnt<3> ), .B(n209), .Y(n165) );
  INVX1 U173 ( .A(n269), .Y(n166) );
  INVX1 U174 ( .A(n166), .Y(n167) );
  INVX1 U175 ( .A(n166), .Y(n168) );
  AND2X1 U176 ( .A(\In<9> ), .B(n7), .Y(n169) );
  INVX1 U177 ( .A(n169), .Y(n170) );
  BUFX2 U178 ( .A(n205), .Y(n171) );
  AND2X2 U179 ( .A(n74), .B(n55), .Y(n173) );
  INVX1 U180 ( .A(n173), .Y(n174) );
  AND2X2 U181 ( .A(n81), .B(n44), .Y(n175) );
  INVX1 U182 ( .A(n175), .Y(n176) );
  AND2X2 U183 ( .A(n85), .B(n46), .Y(n177) );
  INVX1 U184 ( .A(n177), .Y(n178) );
  AND2X2 U185 ( .A(n79), .B(n97), .Y(n179) );
  INVX1 U186 ( .A(n179), .Y(n180) );
  INVX1 U187 ( .A(n210), .Y(n181) );
  AND2X2 U188 ( .A(n84), .B(n45), .Y(n182) );
  INVX1 U189 ( .A(n182), .Y(n183) );
  AND2X2 U190 ( .A(n87), .B(n48), .Y(n184) );
  INVX1 U191 ( .A(n184), .Y(n185) );
  AND2X2 U192 ( .A(n16), .B(n53), .Y(n186) );
  INVX1 U193 ( .A(n186), .Y(n187) );
  AND2X2 U194 ( .A(n82), .B(n99), .Y(n188) );
  INVX1 U195 ( .A(n188), .Y(n189) );
  AND2X2 U196 ( .A(n86), .B(n47), .Y(n190) );
  INVX1 U197 ( .A(n190), .Y(n191) );
  AND2X2 U198 ( .A(n64), .B(n49), .Y(n192) );
  INVX1 U199 ( .A(n192), .Y(n193) );
  AND2X2 U200 ( .A(n89), .B(n50), .Y(n194) );
  INVX1 U201 ( .A(n194), .Y(n195) );
  AND2X2 U202 ( .A(n66), .B(n101), .Y(n196) );
  INVX1 U203 ( .A(n196), .Y(n197) );
  AND2X2 U204 ( .A(n91), .B(n51), .Y(n198) );
  INVX1 U205 ( .A(n198), .Y(n199) );
  AND2X2 U206 ( .A(n167), .B(n14), .Y(n200) );
  AND2X2 U207 ( .A(n180), .B(n275), .Y(n201) );
  INVX2 U208 ( .A(n211), .Y(n275) );
  INVX1 U209 ( .A(n213), .Y(n202) );
  INVX1 U210 ( .A(\Cnt<0> ), .Y(n204) );
  INVX1 U211 ( .A(\Cnt<1> ), .Y(n213) );
  OR2X2 U212 ( .A(n202), .B(n1), .Y(n242) );
  AOI22X1 U213 ( .A(\In<11> ), .B(n164), .C(\In<12> ), .D(n254), .Y(n205) );
  NAND3X1 U214 ( .A(n130), .B(n170), .C(n171), .Y(n269) );
  AOI22X1 U215 ( .A(\In<4> ), .B(n254), .C(\In<3> ), .D(n164), .Y(n208) );
  INVX2 U216 ( .A(\In<1> ), .Y(n206) );
  AOI21X1 U217 ( .A(\In<2> ), .B(n172), .C(n13), .Y(n207) );
  AOI22X1 U218 ( .A(n142), .B(n167), .C(n11), .D(n180), .Y(n217) );
  AOI22X1 U219 ( .A(\In<7> ), .B(n164), .C(\In<8> ), .D(n254), .Y(n210) );
  OR2X2 U220 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n211) );
  MUX2X1 U221 ( .B(n212), .A(n150), .S(n1), .Y(n239) );
  INVX2 U222 ( .A(\In<13> ), .Y(n214) );
  OAI21X1 U223 ( .A(n8), .B(n214), .C(n18), .Y(n215) );
  AOI22X1 U224 ( .A(n14), .B(n4), .C(n275), .D(n187), .Y(n216) );
  AOI22X1 U225 ( .A(\In<13> ), .B(n254), .C(\In<12> ), .D(n164), .Y(n220) );
  INVX2 U226 ( .A(\In<10> ), .Y(n218) );
  AOI21X1 U227 ( .A(\In<11> ), .B(n172), .C(n69), .Y(n219) );
  AOI22X1 U228 ( .A(\In<5> ), .B(n254), .C(\In<4> ), .D(n164), .Y(n222) );
  INVX2 U229 ( .A(\In<2> ), .Y(n241) );
  AOI21X1 U230 ( .A(\In<3> ), .B(n172), .C(n71), .Y(n221) );
  AOI22X1 U231 ( .A(n142), .B(n176), .C(n11), .D(n189), .Y(n229) );
  AOI22X1 U232 ( .A(\In<9> ), .B(n254), .C(\In<8> ), .D(n164), .Y(n225) );
  INVX2 U233 ( .A(\In<6> ), .Y(n223) );
  AOI21X1 U234 ( .A(\In<7> ), .B(n172), .C(n118), .Y(n224) );
  INVX2 U235 ( .A(\In<14> ), .Y(n226) );
  OAI21X1 U236 ( .A(n8), .B(n226), .C(n24), .Y(n227) );
  AOI22X1 U237 ( .A(n14), .B(n183), .C(n275), .D(n174), .Y(n228) );
  AOI22X1 U238 ( .A(\In<14> ), .B(n254), .C(\In<13> ), .D(n164), .Y(n232) );
  INVX2 U239 ( .A(\In<11> ), .Y(n230) );
  AOI21X1 U240 ( .A(\In<12> ), .B(n172), .C(n120), .Y(n231) );
  AOI22X1 U241 ( .A(\In<6> ), .B(n254), .C(\In<5> ), .D(n164), .Y(n235) );
  INVX2 U242 ( .A(\In<3> ), .Y(n233) );
  AOI21X1 U243 ( .A(\In<4> ), .B(n172), .C(n122), .Y(n234) );
  AOI22X1 U244 ( .A(n142), .B(n178), .C(n11), .D(n191), .Y(n244) );
  AOI22X1 U245 ( .A(\In<10> ), .B(n254), .C(\In<9> ), .D(n164), .Y(n238) );
  INVX2 U246 ( .A(\In<7> ), .Y(n236) );
  AOI21X1 U247 ( .A(\In<8> ), .B(n172), .C(n124), .Y(n237) );
  AOI22X1 U248 ( .A(\In<1> ), .B(n164), .C(n202), .D(n239), .Y(n240) );
  OAI21X1 U249 ( .A(n242), .B(n241), .C(n103), .Y(n273) );
  AOI22X1 U250 ( .A(n14), .B(n185), .C(n275), .D(n273), .Y(n243) );
  AOI22X1 U251 ( .A(\In<15> ), .B(n254), .C(\In<14> ), .D(n164), .Y(n247) );
  INVX2 U252 ( .A(\In<12> ), .Y(n245) );
  AOI21X1 U253 ( .A(\In<13> ), .B(n172), .C(n30), .Y(n246) );
  AOI22X1 U254 ( .A(\In<7> ), .B(n254), .C(\In<6> ), .D(n164), .Y(n250) );
  AOI21X1 U255 ( .A(\In<5> ), .B(n172), .C(n32), .Y(n249) );
  AOI22X1 U256 ( .A(n142), .B(n193), .C(n11), .D(n197), .Y(n258) );
  AOI22X1 U257 ( .A(\In<11> ), .B(n254), .C(\In<10> ), .D(n164), .Y(n253) );
  INVX2 U258 ( .A(\In<8> ), .Y(n251) );
  AOI21X1 U259 ( .A(\In<9> ), .B(n172), .C(n126), .Y(n252) );
  AOI22X1 U260 ( .A(\In<3> ), .B(n254), .C(\In<2> ), .D(n164), .Y(n256) );
  AOI21X1 U261 ( .A(\In<1> ), .B(n172), .C(n128), .Y(n255) );
  AOI22X1 U262 ( .A(n14), .B(n195), .C(n275), .D(n199), .Y(n257) );
  NAND3X1 U263 ( .A(n61), .B(n36), .C(n132), .Y(\Out<4> ) );
  AOI22X1 U264 ( .A(n14), .B(n176), .C(n275), .D(n189), .Y(n259) );
  NAND3X1 U265 ( .A(n59), .B(n77), .C(n134), .Y(\Out<5> ) );
  AOI22X1 U266 ( .A(n14), .B(n178), .C(n275), .D(n191), .Y(n260) );
  AOI22X1 U267 ( .A(n6), .B(n199), .C(n11), .D(n195), .Y(n262) );
  AOI22X1 U268 ( .A(n14), .B(n193), .C(n275), .D(n197), .Y(n261) );
  AOI22X1 U269 ( .A(n11), .B(n168), .C(n187), .D(n165), .Y(n264) );
  AOI22X1 U270 ( .A(n275), .B(n4), .C(n180), .D(n6), .Y(n263) );
  AOI22X1 U271 ( .A(n275), .B(n183), .C(n6), .D(n189), .Y(n265) );
  NAND3X1 U272 ( .A(n136), .B(n153), .C(n160), .Y(\Out<9> ) );
  AOI22X1 U273 ( .A(n275), .B(n185), .C(n6), .D(n191), .Y(n266) );
  NAND3X1 U274 ( .A(n73), .B(n155), .C(n161), .Y(\Out<10> ) );
  AOI22X1 U275 ( .A(n11), .B(n193), .C(n165), .D(n199), .Y(n268) );
  AOI22X1 U276 ( .A(n275), .B(n195), .C(n6), .D(n197), .Y(n267) );
  AOI22X1 U277 ( .A(n180), .B(n165), .C(n62), .D(n187), .Y(n271) );
  AOI22X1 U278 ( .A(n168), .B(n275), .C(n6), .D(n4), .Y(n270) );
  AOI22X1 U279 ( .A(n275), .B(n176), .C(n6), .D(n183), .Y(n272) );
  NAND3X1 U280 ( .A(n138), .B(n157), .C(n162), .Y(\Out<13> ) );
  AOI22X1 U281 ( .A(n275), .B(n178), .C(n6), .D(n185), .Y(n274) );
  NAND3X1 U282 ( .A(n140), .B(n159), .C(n163), .Y(\Out<14> ) );
  AOI22X1 U283 ( .A(n165), .B(n197), .C(n62), .D(n199), .Y(n277) );
  AOI22X1 U284 ( .A(n275), .B(n193), .C(n6), .D(n195), .Y(n276) );
endmodule


module rshifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), Rot_sel, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , Rot_sel;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n147, n149, n151, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291;

  INVX4 U2 ( .A(n33), .Y(n34) );
  INVX1 U3 ( .A(\In<4> ), .Y(n239) );
  INVX1 U4 ( .A(\In<3> ), .Y(n226) );
  INVX1 U5 ( .A(\Cnt<3> ), .Y(n221) );
  INVX1 U6 ( .A(\In<6> ), .Y(n268) );
  INVX1 U7 ( .A(\In<10> ), .Y(n263) );
  INVX1 U8 ( .A(\In<14> ), .Y(n260) );
  INVX1 U9 ( .A(\In<8> ), .Y(n236) );
  INVX1 U10 ( .A(\In<12> ), .Y(n233) );
  INVX1 U11 ( .A(\In<15> ), .Y(n218) );
  INVX1 U12 ( .A(\In<7> ), .Y(n222) );
  INVX1 U13 ( .A(n257), .Y(n232) );
  INVX1 U14 ( .A(\Cnt<2> ), .Y(n214) );
  AND2X1 U15 ( .A(n75), .B(n81), .Y(n149) );
  AND2X1 U16 ( .A(n77), .B(n83), .Y(n151) );
  INVX8 U17 ( .A(n245), .Y(n267) );
  AND2X2 U18 ( .A(\Cnt<0> ), .B(\Cnt<1> ), .Y(n33) );
  AND2X2 U19 ( .A(\In<13> ), .B(n267), .Y(n50) );
  AND2X2 U20 ( .A(n215), .B(\Cnt<1> ), .Y(n184) );
  AND2X2 U21 ( .A(n3), .B(n29), .Y(n1) );
  INVX1 U22 ( .A(n1), .Y(\Out<15> ) );
  AND2X2 U23 ( .A(n41), .B(n24), .Y(n3) );
  OR2X2 U24 ( .A(n49), .B(n5), .Y(n4) );
  OR2X2 U25 ( .A(n50), .B(n13), .Y(n5) );
  OR2X2 U26 ( .A(n47), .B(n7), .Y(n6) );
  OR2X2 U27 ( .A(n194), .B(n48), .Y(n7) );
  AND2X2 U28 ( .A(n116), .B(n110), .Y(n8) );
  AND2X2 U29 ( .A(\Cnt<0> ), .B(n216), .Y(n9) );
  INVX1 U30 ( .A(n9), .Y(n10) );
  AND2X2 U31 ( .A(n111), .B(n105), .Y(n11) );
  INVX1 U32 ( .A(n11), .Y(\Out<0> ) );
  AND2X2 U33 ( .A(\Cnt<1> ), .B(n232), .Y(n13) );
  AND2X2 U34 ( .A(n113), .B(n108), .Y(n14) );
  INVX1 U35 ( .A(n14), .Y(n15) );
  OR2X2 U36 ( .A(n34), .B(n268), .Y(n16) );
  INVX1 U37 ( .A(n16), .Y(n17) );
  AND2X2 U38 ( .A(n196), .B(n39), .Y(n18) );
  INVX1 U39 ( .A(n18), .Y(n19) );
  AND2X2 U40 ( .A(n114), .B(n106), .Y(n20) );
  INVX1 U41 ( .A(n20), .Y(\Out<5> ) );
  AND2X1 U42 ( .A(n212), .B(n182), .Y(n22) );
  AND2X2 U43 ( .A(n290), .B(n211), .Y(n23) );
  INVX1 U44 ( .A(n23), .Y(n24) );
  BUFX2 U45 ( .A(n278), .Y(n25) );
  BUFX2 U46 ( .A(n223), .Y(n26) );
  AND2X2 U47 ( .A(n212), .B(n244), .Y(n27) );
  INVX1 U48 ( .A(n27), .Y(n28) );
  BUFX2 U49 ( .A(n291), .Y(n29) );
  BUFX2 U50 ( .A(n287), .Y(n30) );
  AND2X2 U51 ( .A(n36), .B(n4), .Y(n31) );
  INVX1 U52 ( .A(n31), .Y(n32) );
  AND2X2 U53 ( .A(\Cnt<3> ), .B(n214), .Y(n35) );
  AND2X1 U54 ( .A(\Cnt<3> ), .B(\Cnt<2> ), .Y(n36) );
  OR2X2 U55 ( .A(n34), .B(n260), .Y(n37) );
  INVX1 U56 ( .A(n37), .Y(n38) );
  AND2X2 U57 ( .A(n212), .B(n36), .Y(n39) );
  AND2X1 U58 ( .A(n191), .B(n39), .Y(n40) );
  INVX1 U59 ( .A(n40), .Y(n41) );
  OR2X1 U60 ( .A(n34), .B(n263), .Y(n42) );
  INVX1 U61 ( .A(n42), .Y(n43) );
  AND2X1 U62 ( .A(n187), .B(n39), .Y(n44) );
  INVX1 U63 ( .A(n44), .Y(n45) );
  BUFX2 U64 ( .A(n255), .Y(n46) );
  AND2X2 U65 ( .A(\In<10> ), .B(n269), .Y(n47) );
  AND2X1 U66 ( .A(\In<11> ), .B(n33), .Y(n48) );
  AND2X1 U67 ( .A(\In<14> ), .B(n266), .Y(n49) );
  AND2X2 U68 ( .A(n36), .B(n193), .Y(n51) );
  INVX1 U69 ( .A(n51), .Y(n52) );
  AND2X2 U70 ( .A(n36), .B(n289), .Y(n53) );
  INVX1 U71 ( .A(n53), .Y(n54) );
  AND2X1 U72 ( .A(n212), .B(n35), .Y(n55) );
  BUFX2 U73 ( .A(n220), .Y(n56) );
  INVX1 U74 ( .A(n224), .Y(n57) );
  INVX1 U75 ( .A(n57), .Y(n58) );
  BUFX2 U76 ( .A(n228), .Y(n59) );
  BUFX2 U77 ( .A(n235), .Y(n60) );
  BUFX2 U78 ( .A(n238), .Y(n61) );
  BUFX2 U79 ( .A(n241), .Y(n62) );
  BUFX2 U80 ( .A(n248), .Y(n63) );
  BUFX2 U81 ( .A(n251), .Y(n64) );
  BUFX2 U82 ( .A(n254), .Y(n65) );
  INVX1 U83 ( .A(n262), .Y(n66) );
  INVX1 U84 ( .A(n66), .Y(n67) );
  INVX1 U85 ( .A(n271), .Y(n68) );
  INVX1 U86 ( .A(n68), .Y(n69) );
  INVX1 U87 ( .A(n277), .Y(n70) );
  INVX1 U88 ( .A(n70), .Y(n71) );
  INVX1 U89 ( .A(n279), .Y(n72) );
  INVX1 U90 ( .A(n72), .Y(n73) );
  INVX1 U91 ( .A(n281), .Y(n74) );
  INVX1 U92 ( .A(n74), .Y(n75) );
  INVX1 U93 ( .A(n286), .Y(n76) );
  INVX1 U94 ( .A(n76), .Y(n77) );
  INVX1 U95 ( .A(n276), .Y(n78) );
  INVX1 U96 ( .A(n78), .Y(n79) );
  INVX1 U97 ( .A(n280), .Y(n80) );
  INVX1 U98 ( .A(n80), .Y(n81) );
  INVX1 U99 ( .A(n285), .Y(n82) );
  INVX1 U100 ( .A(n82), .Y(n83) );
  INVX1 U101 ( .A(n219), .Y(n84) );
  INVX1 U102 ( .A(n84), .Y(n85) );
  BUFX2 U103 ( .A(n227), .Y(n86) );
  INVX1 U104 ( .A(n234), .Y(n87) );
  INVX1 U105 ( .A(n87), .Y(n88) );
  INVX1 U106 ( .A(n237), .Y(n89) );
  INVX1 U107 ( .A(n89), .Y(n90) );
  INVX1 U108 ( .A(n240), .Y(n91) );
  INVX1 U109 ( .A(n91), .Y(n92) );
  INVX1 U110 ( .A(n247), .Y(n93) );
  INVX1 U111 ( .A(n93), .Y(n94) );
  INVX1 U112 ( .A(n250), .Y(n95) );
  INVX1 U113 ( .A(n95), .Y(n96) );
  INVX1 U114 ( .A(n253), .Y(n97) );
  INVX1 U115 ( .A(n97), .Y(n98) );
  INVX1 U116 ( .A(n261), .Y(n99) );
  INVX1 U117 ( .A(n99), .Y(n100) );
  INVX1 U118 ( .A(n270), .Y(n101) );
  INVX1 U119 ( .A(n101), .Y(n102) );
  AND2X2 U120 ( .A(\In<0> ), .B(n184), .Y(n103) );
  INVX1 U121 ( .A(n103), .Y(n104) );
  BUFX2 U122 ( .A(n229), .Y(n105) );
  BUFX2 U123 ( .A(n274), .Y(n106) );
  INVX1 U124 ( .A(n264), .Y(n107) );
  INVX1 U125 ( .A(n107), .Y(n108) );
  AND2X2 U126 ( .A(\In<15> ), .B(n266), .Y(n109) );
  INVX1 U127 ( .A(n109), .Y(n110) );
  BUFX2 U128 ( .A(n230), .Y(n111) );
  INVX1 U129 ( .A(n265), .Y(n112) );
  INVX1 U130 ( .A(n112), .Y(n113) );
  BUFX2 U131 ( .A(n275), .Y(n114) );
  AND2X2 U132 ( .A(\In<14> ), .B(n267), .Y(n115) );
  INVX1 U133 ( .A(n115), .Y(n116) );
  OR2X1 U134 ( .A(n34), .B(n218), .Y(n117) );
  INVX1 U135 ( .A(n117), .Y(n118) );
  OR2X1 U136 ( .A(n34), .B(n222), .Y(n119) );
  INVX1 U137 ( .A(n119), .Y(n120) );
  OR2X1 U138 ( .A(n34), .B(n226), .Y(n121) );
  INVX1 U139 ( .A(n121), .Y(n122) );
  OR2X2 U140 ( .A(n34), .B(n233), .Y(n123) );
  INVX1 U141 ( .A(n123), .Y(n124) );
  OR2X1 U142 ( .A(n34), .B(n236), .Y(n125) );
  INVX1 U143 ( .A(n125), .Y(n126) );
  OR2X1 U144 ( .A(n34), .B(n239), .Y(n127) );
  INVX1 U145 ( .A(n127), .Y(n128) );
  OR2X2 U146 ( .A(n34), .B(n246), .Y(n129) );
  INVX1 U147 ( .A(n129), .Y(n130) );
  OR2X1 U148 ( .A(n34), .B(n249), .Y(n131) );
  INVX1 U149 ( .A(n131), .Y(n132) );
  OR2X1 U150 ( .A(n34), .B(n252), .Y(n133) );
  INVX1 U151 ( .A(n133), .Y(n134) );
  OR2X2 U152 ( .A(n34), .B(n256), .Y(n135) );
  INVX1 U153 ( .A(n135), .Y(n136) );
  AND2X1 U154 ( .A(n290), .B(n187), .Y(n137) );
  INVX1 U155 ( .A(n137), .Y(n138) );
  AND2X1 U156 ( .A(n290), .B(n189), .Y(n139) );
  INVX1 U157 ( .A(n139), .Y(n140) );
  AND2X1 U158 ( .A(n290), .B(n191), .Y(n141) );
  INVX1 U159 ( .A(n141), .Y(n142) );
  AND2X1 U160 ( .A(n189), .B(n39), .Y(n143) );
  INVX1 U161 ( .A(n143), .Y(n144) );
  AND2X2 U162 ( .A(n71), .B(n79), .Y(n145) );
  INVX1 U163 ( .A(n145), .Y(\Out<6> ) );
  AND2X2 U164 ( .A(n73), .B(n25), .Y(n147) );
  INVX1 U165 ( .A(n147), .Y(\Out<7> ) );
  INVX1 U166 ( .A(n149), .Y(\Out<8> ) );
  INVX1 U167 ( .A(n151), .Y(\Out<12> ) );
  AND2X1 U168 ( .A(n35), .B(n187), .Y(n153) );
  INVX1 U169 ( .A(n153), .Y(n154) );
  AND2X2 U170 ( .A(n35), .B(n189), .Y(n155) );
  INVX1 U171 ( .A(n155), .Y(n156) );
  AND2X2 U172 ( .A(n35), .B(n191), .Y(n157) );
  INVX1 U173 ( .A(n157), .Y(n158) );
  AND2X2 U174 ( .A(n6), .B(n182), .Y(n159) );
  INVX1 U175 ( .A(n159), .Y(n160) );
  AND2X1 U176 ( .A(n182), .B(n4), .Y(n161) );
  INVX1 U177 ( .A(n161), .Y(n162) );
  AND2X1 U178 ( .A(n182), .B(n193), .Y(n163) );
  INVX1 U179 ( .A(n163), .Y(n164) );
  AND2X2 U180 ( .A(n182), .B(n211), .Y(n165) );
  INVX1 U181 ( .A(n165), .Y(n166) );
  AND2X1 U182 ( .A(n290), .B(n4), .Y(n167) );
  INVX1 U183 ( .A(n167), .Y(n168) );
  AND2X1 U184 ( .A(n290), .B(n193), .Y(n169) );
  INVX1 U185 ( .A(n169), .Y(n170) );
  INVX1 U186 ( .A(n242), .Y(n171) );
  INVX1 U187 ( .A(n171), .Y(n172) );
  INVX1 U188 ( .A(n272), .Y(n173) );
  INVX1 U189 ( .A(n173), .Y(n174) );
  BUFX2 U190 ( .A(n273), .Y(n175) );
  INVX1 U191 ( .A(n282), .Y(n176) );
  INVX1 U192 ( .A(n176), .Y(n177) );
  BUFX2 U193 ( .A(n283), .Y(n178) );
  BUFX2 U194 ( .A(n284), .Y(n179) );
  INVX1 U195 ( .A(n288), .Y(n180) );
  INVX1 U196 ( .A(n180), .Y(n181) );
  AND2X1 U197 ( .A(n221), .B(\Cnt<2> ), .Y(n182) );
  BUFX2 U198 ( .A(n259), .Y(n183) );
  INVX1 U199 ( .A(n184), .Y(n185) );
  AND2X2 U200 ( .A(n60), .B(n88), .Y(n186) );
  INVX1 U201 ( .A(n186), .Y(n187) );
  AND2X2 U202 ( .A(n63), .B(n94), .Y(n188) );
  INVX1 U203 ( .A(n188), .Y(n189) );
  AND2X2 U204 ( .A(n67), .B(n100), .Y(n190) );
  INVX1 U205 ( .A(n190), .Y(n191) );
  AND2X2 U206 ( .A(n8), .B(n28), .Y(n192) );
  INVX1 U207 ( .A(n192), .Y(n193) );
  INVX1 U208 ( .A(n217), .Y(n194) );
  AND2X2 U209 ( .A(n59), .B(n86), .Y(n195) );
  INVX1 U210 ( .A(n195), .Y(n196) );
  AND2X2 U211 ( .A(n58), .B(n26), .Y(n197) );
  INVX1 U212 ( .A(n197), .Y(n198) );
  AND2X2 U213 ( .A(n61), .B(n90), .Y(n199) );
  INVX1 U214 ( .A(n199), .Y(n200) );
  AND2X2 U215 ( .A(n64), .B(n96), .Y(n201) );
  INVX1 U216 ( .A(n201), .Y(n202) );
  AND2X2 U217 ( .A(n56), .B(n85), .Y(n203) );
  INVX1 U218 ( .A(n203), .Y(n204) );
  AND2X2 U219 ( .A(n62), .B(n92), .Y(n205) );
  INVX1 U220 ( .A(n205), .Y(n206) );
  AND2X2 U221 ( .A(n65), .B(n98), .Y(n207) );
  INVX1 U222 ( .A(n207), .Y(n208) );
  AND2X2 U223 ( .A(n69), .B(n102), .Y(n209) );
  INVX1 U224 ( .A(n209), .Y(n210) );
  OAI21X1 U225 ( .A(n183), .B(n213), .C(n258), .Y(n211) );
  INVX1 U226 ( .A(\Cnt<1> ), .Y(n216) );
  INVX1 U227 ( .A(\Cnt<0> ), .Y(n215) );
  INVX4 U228 ( .A(n185), .Y(n269) );
  INVX4 U229 ( .A(n10), .Y(n266) );
  INVX8 U230 ( .A(n225), .Y(n290) );
  INVX8 U231 ( .A(n213), .Y(n212) );
  INVX8 U232 ( .A(Rot_sel), .Y(n213) );
  OR2X2 U233 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n245) );
  AOI22X1 U234 ( .A(\In<9> ), .B(n266), .C(\In<8> ), .D(n267), .Y(n217) );
  AOI22X1 U235 ( .A(\In<12> ), .B(n267), .C(\In<13> ), .D(n266), .Y(n220) );
  AOI21X1 U236 ( .A(\In<14> ), .B(n269), .C(n118), .Y(n219) );
  AOI22X1 U237 ( .A(n35), .B(n6), .C(n36), .D(n204), .Y(n230) );
  AOI22X1 U238 ( .A(\In<4> ), .B(n267), .C(\In<5> ), .D(n266), .Y(n224) );
  AOI21X1 U239 ( .A(\In<6> ), .B(n269), .C(n120), .Y(n223) );
  OR2X2 U240 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n225) );
  AOI22X1 U241 ( .A(\In<0> ), .B(n267), .C(\In<1> ), .D(n266), .Y(n228) );
  AOI21X1 U242 ( .A(\In<2> ), .B(n269), .C(n122), .Y(n227) );
  AOI22X1 U243 ( .A(n182), .B(n198), .C(n290), .D(n196), .Y(n229) );
  AND2X2 U244 ( .A(n212), .B(\In<0> ), .Y(n231) );
  MUX2X1 U245 ( .B(\In<15> ), .A(n231), .S(\Cnt<0> ), .Y(n257) );
  AOI22X1 U246 ( .A(\In<9> ), .B(n267), .C(\In<10> ), .D(n266), .Y(n235) );
  AOI21X1 U247 ( .A(\In<11> ), .B(n269), .C(n124), .Y(n234) );
  AOI22X1 U248 ( .A(\In<5> ), .B(n267), .C(\In<6> ), .D(n266), .Y(n238) );
  AOI21X1 U249 ( .A(\In<7> ), .B(n269), .C(n126), .Y(n237) );
  AOI22X1 U250 ( .A(\In<1> ), .B(n267), .C(\In<2> ), .D(n266), .Y(n241) );
  AOI21X1 U251 ( .A(\In<3> ), .B(n269), .C(n128), .Y(n240) );
  AOI22X1 U252 ( .A(n182), .B(n200), .C(n290), .D(n206), .Y(n242) );
  NAND3X1 U253 ( .A(n32), .B(n154), .C(n172), .Y(\Out<1> ) );
  INVX2 U254 ( .A(\In<1> ), .Y(n243) );
  OAI21X1 U255 ( .A(n34), .B(n243), .C(n104), .Y(n244) );
  AOI22X1 U256 ( .A(\In<10> ), .B(n267), .C(\In<11> ), .D(n266), .Y(n248) );
  INVX2 U257 ( .A(\In<13> ), .Y(n246) );
  AOI21X1 U258 ( .A(\In<12> ), .B(n269), .C(n130), .Y(n247) );
  AOI22X1 U259 ( .A(\In<6> ), .B(n267), .C(\In<7> ), .D(n266), .Y(n251) );
  INVX2 U260 ( .A(\In<9> ), .Y(n249) );
  AOI21X1 U261 ( .A(\In<8> ), .B(n269), .C(n132), .Y(n250) );
  AOI22X1 U262 ( .A(\In<2> ), .B(n267), .C(\In<3> ), .D(n266), .Y(n254) );
  INVX2 U263 ( .A(\In<5> ), .Y(n252) );
  AOI21X1 U264 ( .A(\In<4> ), .B(n269), .C(n134), .Y(n253) );
  AOI22X1 U265 ( .A(n182), .B(n202), .C(n290), .D(n208), .Y(n255) );
  NAND3X1 U266 ( .A(n52), .B(n156), .C(n46), .Y(\Out<2> ) );
  INVX2 U267 ( .A(\In<2> ), .Y(n256) );
  AOI21X1 U268 ( .A(\In<1> ), .B(n269), .C(n136), .Y(n259) );
  OR2X2 U269 ( .A(n257), .B(\Cnt<1> ), .Y(n258) );
  OAI21X1 U270 ( .A(n183), .B(n213), .C(n258), .Y(n289) );
  AOI22X1 U271 ( .A(\In<11> ), .B(n267), .C(\In<12> ), .D(n266), .Y(n262) );
  AOI21X1 U272 ( .A(\In<13> ), .B(n269), .C(n38), .Y(n261) );
  AOI22X1 U273 ( .A(\In<7> ), .B(n267), .C(\In<8> ), .D(n266), .Y(n265) );
  AOI21X1 U274 ( .A(\In<9> ), .B(n269), .C(n43), .Y(n264) );
  AOI22X1 U275 ( .A(\In<3> ), .B(n267), .C(\In<4> ), .D(n266), .Y(n271) );
  AOI21X1 U276 ( .A(\In<5> ), .B(n269), .C(n17), .Y(n270) );
  AOI22X1 U277 ( .A(n182), .B(n15), .C(n290), .D(n210), .Y(n272) );
  NAND3X1 U278 ( .A(n54), .B(n158), .C(n174), .Y(\Out<3> ) );
  AOI22X1 U279 ( .A(n290), .B(n198), .C(n204), .D(n35), .Y(n273) );
  NAND3X1 U280 ( .A(n19), .B(n160), .C(n175), .Y(\Out<4> ) );
  AOI22X1 U281 ( .A(n182), .B(n187), .C(n206), .D(n39), .Y(n275) );
  AOI22X1 U282 ( .A(n290), .B(n200), .C(n35), .D(n4), .Y(n274) );
  AOI22X1 U283 ( .A(n182), .B(n189), .C(n208), .D(n39), .Y(n277) );
  AOI22X1 U284 ( .A(n290), .B(n202), .C(n35), .D(n193), .Y(n276) );
  AOI22X1 U285 ( .A(n182), .B(n191), .C(n210), .D(n39), .Y(n279) );
  AOI22X1 U286 ( .A(n290), .B(n15), .C(n35), .D(n211), .Y(n278) );
  AOI22X1 U287 ( .A(n198), .B(n39), .C(n196), .D(n55), .Y(n281) );
  AOI22X1 U288 ( .A(n204), .B(n182), .C(n6), .D(n290), .Y(n280) );
  AOI22X1 U289 ( .A(n200), .B(n39), .C(n206), .D(n55), .Y(n282) );
  NAND3X1 U290 ( .A(n138), .B(n162), .C(n177), .Y(\Out<9> ) );
  AOI22X1 U291 ( .A(n202), .B(n39), .C(n208), .D(n55), .Y(n283) );
  NAND3X1 U292 ( .A(n140), .B(n164), .C(n178), .Y(\Out<10> ) );
  AOI22X1 U293 ( .A(n15), .B(n39), .C(n210), .D(n55), .Y(n284) );
  NAND3X1 U294 ( .A(n142), .B(n166), .C(n179), .Y(\Out<11> ) );
  AOI22X1 U295 ( .A(n198), .B(n55), .C(n196), .D(n22), .Y(n286) );
  AOI22X1 U296 ( .A(n204), .B(n290), .C(n6), .D(n39), .Y(n285) );
  AOI22X1 U297 ( .A(n200), .B(n55), .C(n206), .D(n22), .Y(n287) );
  NAND3X1 U298 ( .A(n30), .B(n45), .C(n168), .Y(\Out<13> ) );
  AOI22X1 U299 ( .A(n202), .B(n55), .C(n208), .D(n22), .Y(n288) );
  NAND3X1 U300 ( .A(n144), .B(n170), .C(n181), .Y(\Out<14> ) );
  AOI22X1 U301 ( .A(n15), .B(n55), .C(n210), .D(n22), .Y(n291) );
endmodule


module fulladder1_31 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_30 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_29 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_28 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_27 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_26 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_25 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_24 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_23 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_22 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_21 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_20 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_19 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_18 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_17 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_16 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module cla4_11 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n11,
         n13, n14, n15, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37;

  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n18), .C(n20), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n20), .C(n19), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n16), .C(\G<2> ), .Y(n11) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n13) );
  OAI21X1 U13 ( .A(n9), .B(n20), .C(n19), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n14) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n15) );
  fulladder1_44 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_45 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_46 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n35), .G(n27) );
  fulladder1_47 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  AND2X1 U1 ( .A(n21), .B(n2), .Y(n10) );
  INVX1 U2 ( .A(\G<0> ), .Y(n21) );
  AND2X1 U3 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  INVX1 U4 ( .A(\P<2> ), .Y(n18) );
  AND2X1 U5 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X1 U6 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  INVX1 U7 ( .A(\G<3> ), .Y(n19) );
  AND2X1 U9 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  INVX1 U16 ( .A(\P<3> ), .Y(n20) );
  AND2X1 U17 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U18 ( .A(n1), .Y(n2) );
  BUFX2 U19 ( .A(n15), .Y(n3) );
  INVX1 U20 ( .A(n3), .Y(n17) );
  INVX1 U21 ( .A(n13), .Y(n16) );
  INVX1 U22 ( .A(n11), .Y(n4) );
  INVX1 U23 ( .A(n4), .Y(n5) );
  AND2X1 U24 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U25 ( .A(n6), .Y(n7) );
  INVX1 U26 ( .A(n9), .Y(n8) );
  BUFX2 U27 ( .A(n14), .Y(n9) );
  INVX1 U28 ( .A(n10), .Y(n12) );
  AND2X1 U29 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U30 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U31 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U32 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U33 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U34 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U35 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U36 ( .A(n22), .B(n23), .Y(\G<0> ) );
endmodule


module cla4_10 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n8), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n6), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n10), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_43 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_42 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_41 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_40 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n9), .S(\S<3> ), .P(n38), .G(n30) );
  AND2X1 U1 ( .A(n18), .B(n2), .Y(n12) );
  INVX1 U2 ( .A(\G<0> ), .Y(n18) );
  AND2X1 U3 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  INVX1 U4 ( .A(\P<2> ), .Y(n20) );
  AND2X1 U5 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  INVX1 U6 ( .A(\G<3> ), .Y(n21) );
  AND2X1 U7 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  INVX1 U9 ( .A(\P<3> ), .Y(n22) );
  AND2X2 U16 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U17 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U18 ( .A(n1), .Y(n2) );
  BUFX2 U19 ( .A(n39), .Y(n3) );
  INVX1 U20 ( .A(n3), .Y(n17) );
  BUFX2 U21 ( .A(n41), .Y(n4) );
  INVX1 U22 ( .A(n4), .Y(n19) );
  INVX1 U23 ( .A(n42), .Y(n5) );
  INVX1 U24 ( .A(n5), .Y(n6) );
  AND2X1 U25 ( .A(\P<1> ), .B(\P<0> ), .Y(n7) );
  INVX1 U26 ( .A(n7), .Y(n8) );
  INVX1 U27 ( .A(n10), .Y(n9) );
  BUFX2 U28 ( .A(n40), .Y(n10) );
  INVX1 U29 ( .A(n12), .Y(n16) );
  AND2X1 U30 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U31 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U32 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U33 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U34 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U35 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U36 ( .A(n23), .B(n24), .Y(\G<0> ) );
endmodule


module cla4_9 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n7), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n9), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_39 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_38 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_37 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_36 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n38), .G(n30) );
  AND2X1 U1 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  AND2X1 U2 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  AND2X1 U3 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  INVX1 U4 ( .A(\P<2> ), .Y(n20) );
  INVX1 U5 ( .A(\G<3> ), .Y(n21) );
  AND2X1 U6 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  INVX1 U7 ( .A(\P<3> ), .Y(n22) );
  AND2X2 U9 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U16 ( .A(n1), .Y(n2) );
  BUFX2 U17 ( .A(n39), .Y(n3) );
  INVX1 U18 ( .A(n3), .Y(n17) );
  BUFX2 U19 ( .A(n41), .Y(n4) );
  INVX1 U20 ( .A(n4), .Y(n19) );
  BUFX2 U21 ( .A(n42), .Y(n5) );
  AND2X1 U22 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U23 ( .A(n6), .Y(n7) );
  INVX1 U24 ( .A(n10), .Y(n8) );
  INVX1 U25 ( .A(n8), .Y(n9) );
  BUFX2 U26 ( .A(n40), .Y(n10) );
  AND2X2 U27 ( .A(n2), .B(n18), .Y(n12) );
  INVX1 U28 ( .A(n12), .Y(n16) );
  AND2X1 U29 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U30 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U31 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U32 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U33 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U34 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U35 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U36 ( .A(n23), .B(n24), .Y(\G<0> ) );
  INVX2 U37 ( .A(\G<0> ), .Y(n18) );
endmodule


module cla4_8 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n19), .C(n21), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n21), .C(n20), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n18), .C(\G<2> ), .Y(n41) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n40) );
  OAI21X1 U13 ( .A(n9), .B(n21), .C(n20), .Y(Cout) );
  AOI21X1 U14 ( .A(n16), .B(\P<2> ), .C(\G<2> ), .Y(n39) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n38) );
  fulladder1_35 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_34 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_33 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n1), .S(\S<2> ), .P(n35), .G(n27) );
  fulladder1_32 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  AND2X1 U1 ( .A(Cin), .B(\P<0> ), .Y(n2) );
  AND2X1 U2 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  AND2X1 U3 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X1 U4 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  INVX1 U5 ( .A(\P<2> ), .Y(n19) );
  INVX1 U6 ( .A(\G<3> ), .Y(n20) );
  AND2X1 U7 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  INVX1 U9 ( .A(\P<3> ), .Y(n21) );
  BUFX2 U16 ( .A(n16), .Y(n1) );
  INVX1 U17 ( .A(n38), .Y(n16) );
  INVX1 U18 ( .A(n2), .Y(n3) );
  BUFX2 U19 ( .A(n40), .Y(n4) );
  INVX1 U20 ( .A(n4), .Y(n18) );
  BUFX2 U21 ( .A(n41), .Y(n5) );
  AND2X1 U22 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U23 ( .A(n6), .Y(n7) );
  INVX1 U24 ( .A(n39), .Y(n8) );
  INVX1 U25 ( .A(n8), .Y(n9) );
  AND2X2 U26 ( .A(n3), .B(n17), .Y(n10) );
  INVX1 U27 ( .A(n10), .Y(n12) );
  AND2X1 U28 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U29 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U30 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U31 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U32 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U33 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U34 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U35 ( .A(n22), .B(n23), .Y(\G<0> ) );
  INVX2 U36 ( .A(\G<0> ), .Y(n17) );
endmodule


module rf ( .read1data({\read1data<15> , \read1data<14> , \read1data<13> , 
        \read1data<12> , \read1data<11> , \read1data<10> , \read1data<9> , 
        \read1data<8> , \read1data<7> , \read1data<6> , \read1data<5> , 
        \read1data<4> , \read1data<3> , \read1data<2> , \read1data<1> , 
        \read1data<0> }), .read2data({\read2data<15> , \read2data<14> , 
        \read2data<13> , \read2data<12> , \read2data<11> , \read2data<10> , 
        \read2data<9> , \read2data<8> , \read2data<7> , \read2data<6> , 
        \read2data<5> , \read2data<4> , \read2data<3> , \read2data<2> , 
        \read2data<1> , \read2data<0> }), err, clk, rst, .read1regsel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .read2regsel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .writeregsel({
        \writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   \rf_wr_en<7> , \rf_wr_en<6> , \rf_wr_en<5> , \rf_wr_en<4> ,
         \rf_wr_en<3> , \rf_wr_en<2> , \rf_wr_en<1> , \rf_wr_en<0> ,
         \write_en<7> , \write_en<6> , \write_en<5> , \write_en<4> ,
         \write_en<3> , \write_en<2> , \write_en<1> , \write_en<0> ,
         \reg_in<127> , \reg_in<126> , \reg_in<125> , \reg_in<124> ,
         \reg_in<123> , \reg_in<122> , \reg_in<121> , \reg_in<120> ,
         \reg_in<119> , \reg_in<118> , \reg_in<117> , \reg_in<116> ,
         \reg_in<115> , \reg_in<114> , \reg_in<113> , \reg_in<112> ,
         \reg_in<111> , \reg_in<110> , \reg_in<109> , \reg_in<108> ,
         \reg_in<107> , \reg_in<106> , \reg_in<105> , \reg_in<104> ,
         \reg_in<103> , \reg_in<102> , \reg_in<101> , \reg_in<100> ,
         \reg_in<99> , \reg_in<98> , \reg_in<97> , \reg_in<96> , \reg_in<95> ,
         \reg_in<94> , \reg_in<93> , \reg_in<92> , \reg_in<91> , \reg_in<90> ,
         \reg_in<89> , \reg_in<88> , \reg_in<87> , \reg_in<86> , \reg_in<85> ,
         \reg_in<84> , \reg_in<83> , \reg_in<82> , \reg_in<81> , \reg_in<80> ,
         \reg_in<79> , \reg_in<78> , \reg_in<77> , \reg_in<76> , \reg_in<75> ,
         \reg_in<74> , \reg_in<73> , \reg_in<72> , \reg_in<71> , \reg_in<70> ,
         \reg_in<69> , \reg_in<68> , \reg_in<67> , \reg_in<66> , \reg_in<65> ,
         \reg_in<64> , \reg_in<63> , \reg_in<62> , \reg_in<61> , \reg_in<60> ,
         \reg_in<59> , \reg_in<58> , \reg_in<57> , \reg_in<56> , \reg_in<55> ,
         \reg_in<54> , \reg_in<53> , \reg_in<52> , \reg_in<51> , \reg_in<50> ,
         \reg_in<49> , \reg_in<48> , \reg_in<47> , \reg_in<46> , \reg_in<45> ,
         \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> ,
         \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> ,
         \reg_in<34> , \reg_in<33> , \reg_in<32> , \reg_in<31> , \reg_in<30> ,
         \reg_in<29> , \reg_in<28> , \reg_in<27> , \reg_in<26> , \reg_in<25> ,
         \reg_in<24> , \reg_in<23> , \reg_in<22> , \reg_in<21> , \reg_in<20> ,
         \reg_in<19> , \reg_in<18> , \reg_in<17> , \reg_in<16> , \reg_in<15> ,
         \reg_in<14> , \reg_in<13> , \reg_in<12> , \reg_in<11> , \reg_in<10> ,
         \reg_in<9> , \reg_in<8> , \reg_in<7> , \reg_in<6> , \reg_in<5> ,
         \reg_in<4> , \reg_in<3> , \reg_in<2> , \reg_in<1> , \reg_in<0> ,
         \reg_out<127> , \reg_out<126> , \reg_out<125> , \reg_out<124> ,
         \reg_out<123> , \reg_out<122> , \reg_out<121> , \reg_out<120> ,
         \reg_out<119> , \reg_out<118> , \reg_out<117> , \reg_out<116> ,
         \reg_out<115> , \reg_out<114> , \reg_out<113> , \reg_out<112> ,
         \reg_out<111> , \reg_out<110> , \reg_out<109> , \reg_out<108> ,
         \reg_out<107> , \reg_out<106> , \reg_out<105> , \reg_out<104> ,
         \reg_out<103> , \reg_out<102> , \reg_out<101> , \reg_out<100> ,
         \reg_out<99> , \reg_out<98> , \reg_out<97> , \reg_out<96> ,
         \reg_out<95> , \reg_out<94> , \reg_out<93> , \reg_out<92> ,
         \reg_out<91> , \reg_out<90> , \reg_out<89> , \reg_out<88> ,
         \reg_out<87> , \reg_out<86> , \reg_out<85> , \reg_out<84> ,
         \reg_out<83> , \reg_out<82> , \reg_out<81> , \reg_out<80> ,
         \reg_out<79> , \reg_out<78> , \reg_out<77> , \reg_out<76> ,
         \reg_out<75> , \reg_out<74> , \reg_out<73> , \reg_out<72> ,
         \reg_out<71> , \reg_out<70> , \reg_out<69> , \reg_out<68> ,
         \reg_out<67> , \reg_out<66> , \reg_out<65> , \reg_out<64> ,
         \reg_out<63> , \reg_out<62> , \reg_out<61> , \reg_out<60> ,
         \reg_out<59> , \reg_out<58> , \reg_out<57> , \reg_out<56> ,
         \reg_out<55> , \reg_out<54> , \reg_out<53> , \reg_out<52> ,
         \reg_out<51> , \reg_out<50> , \reg_out<49> , \reg_out<48> ,
         \reg_out<47> , \reg_out<46> , \reg_out<45> , \reg_out<44> ,
         \reg_out<43> , \reg_out<42> , \reg_out<41> , \reg_out<40> ,
         \reg_out<39> , \reg_out<38> , \reg_out<37> , \reg_out<36> ,
         \reg_out<35> , \reg_out<34> , \reg_out<33> , \reg_out<32> ,
         \reg_out<31> , \reg_out<30> , \reg_out<29> , \reg_out<28> ,
         \reg_out<27> , \reg_out<26> , \reg_out<25> , \reg_out<24> ,
         \reg_out<23> , \reg_out<22> , \reg_out<21> , \reg_out<20> ,
         \reg_out<19> , \reg_out<18> , \reg_out<17> , \reg_out<16> ,
         \reg_out<15> , \reg_out<14> , \reg_out<13> , \reg_out<12> ,
         \reg_out<11> , \reg_out<10> , \reg_out<9> , \reg_out<8> ,
         \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , \reg_out<3> ,
         \reg_out<2> , \reg_out<1> , \reg_out<0> , n1, n2, n3, n4;
  assign err = 1'b0;

  register16_0 \registers[0]  ( .d({\reg_in<15> , \reg_in<14> , \reg_in<13> , 
        \reg_in<12> , \reg_in<11> , \reg_in<10> , \reg_in<9> , \reg_in<8> , 
        \reg_in<7> , \reg_in<6> , \reg_in<5> , \reg_in<4> , \reg_in<3> , 
        \reg_in<2> , \reg_in<1> , \reg_in<0> }), .clk(clk), .wr_en(
        \rf_wr_en<0> ), .rst(n3), .q({\reg_out<15> , \reg_out<14> , 
        \reg_out<13> , \reg_out<12> , \reg_out<11> , \reg_out<10> , 
        \reg_out<9> , \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , 
        \reg_out<4> , \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> })
         );
  register16_1 \registers[1]  ( .d({\reg_in<31> , \reg_in<30> , \reg_in<29> , 
        \reg_in<28> , \reg_in<27> , \reg_in<26> , \reg_in<25> , \reg_in<24> , 
        \reg_in<23> , \reg_in<22> , \reg_in<21> , \reg_in<20> , \reg_in<19> , 
        \reg_in<18> , \reg_in<17> , \reg_in<16> }), .clk(clk), .wr_en(
        \rf_wr_en<1> ), .rst(n3), .q({\reg_out<31> , \reg_out<30> , 
        \reg_out<29> , \reg_out<28> , \reg_out<27> , \reg_out<26> , 
        \reg_out<25> , \reg_out<24> , \reg_out<23> , \reg_out<22> , 
        \reg_out<21> , \reg_out<20> , \reg_out<19> , \reg_out<18> , 
        \reg_out<17> , \reg_out<16> }) );
  register16_2 \registers[2]  ( .d({\reg_in<47> , \reg_in<46> , \reg_in<45> , 
        \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> , 
        \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> , 
        \reg_in<34> , \reg_in<33> , \reg_in<32> }), .clk(clk), .wr_en(
        \rf_wr_en<2> ), .rst(n3), .q({\reg_out<47> , \reg_out<46> , 
        \reg_out<45> , \reg_out<44> , \reg_out<43> , \reg_out<42> , 
        \reg_out<41> , \reg_out<40> , \reg_out<39> , \reg_out<38> , 
        \reg_out<37> , \reg_out<36> , \reg_out<35> , \reg_out<34> , 
        \reg_out<33> , \reg_out<32> }) );
  register16_3 \registers[3]  ( .d({\reg_in<63> , \reg_in<62> , \reg_in<61> , 
        \reg_in<60> , \reg_in<59> , \reg_in<58> , \reg_in<57> , \reg_in<56> , 
        \reg_in<55> , \reg_in<54> , \reg_in<53> , \reg_in<52> , \reg_in<51> , 
        \reg_in<50> , \reg_in<49> , \reg_in<48> }), .clk(clk), .wr_en(
        \rf_wr_en<3> ), .rst(n3), .q({\reg_out<63> , \reg_out<62> , 
        \reg_out<61> , \reg_out<60> , \reg_out<59> , \reg_out<58> , 
        \reg_out<57> , \reg_out<56> , \reg_out<55> , \reg_out<54> , 
        \reg_out<53> , \reg_out<52> , \reg_out<51> , \reg_out<50> , 
        \reg_out<49> , \reg_out<48> }) );
  register16_4 \registers[4]  ( .d({\reg_in<79> , \reg_in<78> , \reg_in<77> , 
        \reg_in<76> , \reg_in<75> , \reg_in<74> , \reg_in<73> , \reg_in<72> , 
        \reg_in<71> , \reg_in<70> , \reg_in<69> , \reg_in<68> , \reg_in<67> , 
        \reg_in<66> , \reg_in<65> , \reg_in<64> }), .clk(clk), .wr_en(
        \rf_wr_en<4> ), .rst(n3), .q({\reg_out<79> , \reg_out<78> , 
        \reg_out<77> , \reg_out<76> , \reg_out<75> , \reg_out<74> , 
        \reg_out<73> , \reg_out<72> , \reg_out<71> , \reg_out<70> , 
        \reg_out<69> , \reg_out<68> , \reg_out<67> , \reg_out<66> , 
        \reg_out<65> , \reg_out<64> }) );
  register16_5 \registers[5]  ( .d({\reg_in<95> , \reg_in<94> , \reg_in<93> , 
        \reg_in<92> , \reg_in<91> , \reg_in<90> , \reg_in<89> , \reg_in<88> , 
        \reg_in<87> , \reg_in<86> , \reg_in<85> , \reg_in<84> , \reg_in<83> , 
        \reg_in<82> , \reg_in<81> , \reg_in<80> }), .clk(clk), .wr_en(
        \rf_wr_en<5> ), .rst(n3), .q({\reg_out<95> , \reg_out<94> , 
        \reg_out<93> , \reg_out<92> , \reg_out<91> , \reg_out<90> , 
        \reg_out<89> , \reg_out<88> , \reg_out<87> , \reg_out<86> , 
        \reg_out<85> , \reg_out<84> , \reg_out<83> , \reg_out<82> , 
        \reg_out<81> , \reg_out<80> }) );
  register16_6 \registers[6]  ( .d({\reg_in<111> , \reg_in<110> , 
        \reg_in<109> , \reg_in<108> , \reg_in<107> , \reg_in<106> , 
        \reg_in<105> , \reg_in<104> , \reg_in<103> , \reg_in<102> , 
        \reg_in<101> , \reg_in<100> , \reg_in<99> , \reg_in<98> , \reg_in<97> , 
        \reg_in<96> }), .clk(clk), .wr_en(\rf_wr_en<6> ), .rst(n3), .q({
        \reg_out<111> , \reg_out<110> , \reg_out<109> , \reg_out<108> , 
        \reg_out<107> , \reg_out<106> , \reg_out<105> , \reg_out<104> , 
        \reg_out<103> , \reg_out<102> , \reg_out<101> , \reg_out<100> , 
        \reg_out<99> , \reg_out<98> , \reg_out<97> , \reg_out<96> }) );
  register16_7 \registers[7]  ( .d({\reg_in<127> , \reg_in<126> , 
        \reg_in<125> , \reg_in<124> , \reg_in<123> , \reg_in<122> , 
        \reg_in<121> , \reg_in<120> , \reg_in<119> , \reg_in<118> , 
        \reg_in<117> , \reg_in<116> , \reg_in<115> , \reg_in<114> , 
        \reg_in<113> , \reg_in<112> }), .clk(clk), .wr_en(\rf_wr_en<7> ), 
        .rst(n3), .q({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> }) );
  decoder3to8 wr_dec ( .In({\writeregsel<2> , \writeregsel<1> , n1}), .Out({
        \write_en<7> , \write_en<6> , \write_en<5> , \write_en<4> , 
        \write_en<3> , \write_en<2> , \write_en<1> , \write_en<0> }) );
  mux8to1_16_1 read1_mux ( .In({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> , \reg_out<111> , \reg_out<110> , \reg_out<109> , 
        \reg_out<108> , \reg_out<107> , \reg_out<106> , \reg_out<105> , 
        \reg_out<104> , \reg_out<103> , \reg_out<102> , \reg_out<101> , 
        \reg_out<100> , \reg_out<99> , \reg_out<98> , \reg_out<97> , 
        \reg_out<96> , \reg_out<95> , \reg_out<94> , \reg_out<93> , 
        \reg_out<92> , \reg_out<91> , \reg_out<90> , \reg_out<89> , 
        \reg_out<88> , \reg_out<87> , \reg_out<86> , \reg_out<85> , 
        \reg_out<84> , \reg_out<83> , \reg_out<82> , \reg_out<81> , 
        \reg_out<80> , \reg_out<79> , \reg_out<78> , \reg_out<77> , 
        \reg_out<76> , \reg_out<75> , \reg_out<74> , \reg_out<73> , 
        \reg_out<72> , \reg_out<71> , \reg_out<70> , \reg_out<69> , 
        \reg_out<68> , \reg_out<67> , \reg_out<66> , \reg_out<65> , 
        \reg_out<64> , \reg_out<63> , \reg_out<62> , \reg_out<61> , 
        \reg_out<60> , \reg_out<59> , \reg_out<58> , \reg_out<57> , 
        \reg_out<56> , \reg_out<55> , \reg_out<54> , \reg_out<53> , 
        \reg_out<52> , \reg_out<51> , \reg_out<50> , \reg_out<49> , 
        \reg_out<48> , \reg_out<47> , \reg_out<46> , \reg_out<45> , 
        \reg_out<44> , \reg_out<43> , \reg_out<42> , \reg_out<41> , 
        \reg_out<40> , \reg_out<39> , \reg_out<38> , \reg_out<37> , 
        \reg_out<36> , \reg_out<35> , \reg_out<34> , \reg_out<33> , 
        \reg_out<32> , \reg_out<31> , \reg_out<30> , \reg_out<29> , 
        \reg_out<28> , \reg_out<27> , \reg_out<26> , \reg_out<25> , 
        \reg_out<24> , \reg_out<23> , \reg_out<22> , \reg_out<21> , 
        \reg_out<20> , \reg_out<19> , \reg_out<18> , \reg_out<17> , 
        \reg_out<16> , \reg_out<15> , \reg_out<14> , \reg_out<13> , 
        \reg_out<12> , \reg_out<11> , \reg_out<10> , \reg_out<9> , 
        \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , 
        \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> }), .Sel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .Out({
        \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> , 
        \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> , 
        \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> , 
        \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> }) );
  mux8to1_16_0 read2_mux ( .In({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> , \reg_out<111> , \reg_out<110> , \reg_out<109> , 
        \reg_out<108> , \reg_out<107> , \reg_out<106> , \reg_out<105> , 
        \reg_out<104> , \reg_out<103> , \reg_out<102> , \reg_out<101> , 
        \reg_out<100> , \reg_out<99> , \reg_out<98> , \reg_out<97> , 
        \reg_out<96> , \reg_out<95> , \reg_out<94> , \reg_out<93> , 
        \reg_out<92> , \reg_out<91> , \reg_out<90> , \reg_out<89> , 
        \reg_out<88> , \reg_out<87> , \reg_out<86> , \reg_out<85> , 
        \reg_out<84> , \reg_out<83> , \reg_out<82> , \reg_out<81> , 
        \reg_out<80> , \reg_out<79> , \reg_out<78> , \reg_out<77> , 
        \reg_out<76> , \reg_out<75> , \reg_out<74> , \reg_out<73> , 
        \reg_out<72> , \reg_out<71> , \reg_out<70> , \reg_out<69> , 
        \reg_out<68> , \reg_out<67> , \reg_out<66> , \reg_out<65> , 
        \reg_out<64> , \reg_out<63> , \reg_out<62> , \reg_out<61> , 
        \reg_out<60> , \reg_out<59> , \reg_out<58> , \reg_out<57> , 
        \reg_out<56> , \reg_out<55> , \reg_out<54> , \reg_out<53> , 
        \reg_out<52> , \reg_out<51> , \reg_out<50> , \reg_out<49> , 
        \reg_out<48> , \reg_out<47> , \reg_out<46> , \reg_out<45> , 
        \reg_out<44> , \reg_out<43> , \reg_out<42> , \reg_out<41> , 
        \reg_out<40> , \reg_out<39> , \reg_out<38> , \reg_out<37> , 
        \reg_out<36> , \reg_out<35> , \reg_out<34> , \reg_out<33> , 
        \reg_out<32> , \reg_out<31> , \reg_out<30> , \reg_out<29> , 
        \reg_out<28> , \reg_out<27> , \reg_out<26> , \reg_out<25> , 
        \reg_out<24> , \reg_out<23> , \reg_out<22> , \reg_out<21> , 
        \reg_out<20> , \reg_out<19> , \reg_out<18> , \reg_out<17> , 
        \reg_out<16> , \reg_out<15> , \reg_out<14> , \reg_out<13> , 
        \reg_out<12> , \reg_out<11> , \reg_out<10> , \reg_out<9> , 
        \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , 
        \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> }), .Sel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .Out({
        \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> , 
        \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> , 
        \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> , 
        \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> }) );
  demux1to8_16 wr_demux ( .In({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .S({\writeregsel<2> , 
        \writeregsel<1> , n1}), .Out0({\reg_in<15> , \reg_in<14> , 
        \reg_in<13> , \reg_in<12> , \reg_in<11> , \reg_in<10> , \reg_in<9> , 
        \reg_in<8> , \reg_in<7> , \reg_in<6> , \reg_in<5> , \reg_in<4> , 
        \reg_in<3> , \reg_in<2> , \reg_in<1> , \reg_in<0> }), .Out1({
        \reg_in<31> , \reg_in<30> , \reg_in<29> , \reg_in<28> , \reg_in<27> , 
        \reg_in<26> , \reg_in<25> , \reg_in<24> , \reg_in<23> , \reg_in<22> , 
        \reg_in<21> , \reg_in<20> , \reg_in<19> , \reg_in<18> , \reg_in<17> , 
        \reg_in<16> }), .Out2({\reg_in<47> , \reg_in<46> , \reg_in<45> , 
        \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> , 
        \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> , 
        \reg_in<34> , \reg_in<33> , \reg_in<32> }), .Out3({\reg_in<63> , 
        \reg_in<62> , \reg_in<61> , \reg_in<60> , \reg_in<59> , \reg_in<58> , 
        \reg_in<57> , \reg_in<56> , \reg_in<55> , \reg_in<54> , \reg_in<53> , 
        \reg_in<52> , \reg_in<51> , \reg_in<50> , \reg_in<49> , \reg_in<48> }), 
        .Out4({\reg_in<79> , \reg_in<78> , \reg_in<77> , \reg_in<76> , 
        \reg_in<75> , \reg_in<74> , \reg_in<73> , \reg_in<72> , \reg_in<71> , 
        \reg_in<70> , \reg_in<69> , \reg_in<68> , \reg_in<67> , \reg_in<66> , 
        \reg_in<65> , \reg_in<64> }), .Out5({\reg_in<95> , \reg_in<94> , 
        \reg_in<93> , \reg_in<92> , \reg_in<91> , \reg_in<90> , \reg_in<89> , 
        \reg_in<88> , \reg_in<87> , \reg_in<86> , \reg_in<85> , \reg_in<84> , 
        \reg_in<83> , \reg_in<82> , \reg_in<81> , \reg_in<80> }), .Out6({
        \reg_in<111> , \reg_in<110> , \reg_in<109> , \reg_in<108> , 
        \reg_in<107> , \reg_in<106> , \reg_in<105> , \reg_in<104> , 
        \reg_in<103> , \reg_in<102> , \reg_in<101> , \reg_in<100> , 
        \reg_in<99> , \reg_in<98> , \reg_in<97> , \reg_in<96> }), .Out7({
        \reg_in<127> , \reg_in<126> , \reg_in<125> , \reg_in<124> , 
        \reg_in<123> , \reg_in<122> , \reg_in<121> , \reg_in<120> , 
        \reg_in<119> , \reg_in<118> , \reg_in<117> , \reg_in<116> , 
        \reg_in<115> , \reg_in<114> , \reg_in<113> , \reg_in<112> }) );
  AND2X1 U2 ( .A(\write_en<0> ), .B(write), .Y(\rf_wr_en<0> ) );
  AND2X1 U3 ( .A(\write_en<1> ), .B(write), .Y(\rf_wr_en<1> ) );
  AND2X1 U4 ( .A(\write_en<2> ), .B(write), .Y(\rf_wr_en<2> ) );
  AND2X1 U5 ( .A(\write_en<3> ), .B(write), .Y(\rf_wr_en<3> ) );
  AND2X1 U6 ( .A(\write_en<4> ), .B(write), .Y(\rf_wr_en<4> ) );
  AND2X1 U7 ( .A(\write_en<5> ), .B(write), .Y(\rf_wr_en<5> ) );
  AND2X1 U8 ( .A(\write_en<6> ), .B(write), .Y(\rf_wr_en<6> ) );
  AND2X1 U9 ( .A(\write_en<7> ), .B(write), .Y(\rf_wr_en<7> ) );
  INVX2 U10 ( .A(n2), .Y(n1) );
  INVX1 U11 ( .A(\writeregsel<0> ), .Y(n2) );
  INVX2 U12 ( .A(n4), .Y(n3) );
  INVX1 U13 ( .A(rst), .Y(n4) );
endmodule


module demux1to2_16_1 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), S, .Out0({\Out0<15> , \Out0<14> , 
        \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , \Out0<9> , \Out0<8> , 
        \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , \Out0<3> , \Out0<2> , 
        \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , \Out1<14> , \Out1<13> , 
        \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , \Out1<8> , \Out1<7> , 
        \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , \Out1<2> , \Out1<1> , 
        \Out1<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , S;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> ;
  wire   n1, n2, n3;

  demux1to2_17 \d[0]  ( .In(\In<0> ), .S(n1), .Out0(\Out0<0> ), .Out1(
        \Out1<0> ) );
  demux1to2_18 \d[1]  ( .In(\In<1> ), .S(n2), .Out0(\Out0<1> ), .Out1(
        \Out1<1> ) );
  demux1to2_19 \d[2]  ( .In(\In<2> ), .S(n2), .Out0(\Out0<2> ), .Out1(
        \Out1<2> ) );
  demux1to2_20 \d[3]  ( .In(\In<3> ), .S(n2), .Out0(\Out0<3> ), .Out1(
        \Out1<3> ) );
  demux1to2_21 \d[4]  ( .In(\In<4> ), .S(n2), .Out0(\Out0<4> ), .Out1(
        \Out1<4> ) );
  demux1to2_22 \d[5]  ( .In(\In<5> ), .S(n1), .Out0(\Out0<5> ), .Out1(
        \Out1<5> ) );
  demux1to2_23 \d[6]  ( .In(\In<6> ), .S(n1), .Out0(\Out0<6> ), .Out1(
        \Out1<6> ) );
  demux1to2_24 \d[7]  ( .In(\In<7> ), .S(n1), .Out0(\Out0<7> ), .Out1(
        \Out1<7> ) );
  demux1to2_25 \d[8]  ( .In(\In<8> ), .S(n1), .Out0(\Out0<8> ), .Out1(
        \Out1<8> ) );
  demux1to2_26 \d[9]  ( .In(\In<9> ), .S(n1), .Out0(\Out0<9> ), .Out1(
        \Out1<9> ) );
  demux1to2_27 \d[10]  ( .In(\In<10> ), .S(n1), .Out0(\Out0<10> ), .Out1(
        \Out1<10> ) );
  demux1to2_28 \d[11]  ( .In(\In<11> ), .S(n1), .Out0(\Out0<11> ), .Out1(
        \Out1<11> ) );
  demux1to2_29 \d[12]  ( .In(\In<12> ), .S(n1), .Out0(\Out0<12> ), .Out1(
        \Out1<12> ) );
  demux1to2_30 \d[13]  ( .In(\In<13> ), .S(n1), .Out0(\Out0<13> ), .Out1(
        \Out1<13> ) );
  demux1to2_31 \d[14]  ( .In(\In<14> ), .S(n1), .Out0(\Out0<14> ), .Out1(
        \Out1<14> ) );
  demux1to2_32 \d[15]  ( .In(\In<15> ), .S(n1), .Out0(\Out0<15> ), .Out1(
        \Out1<15> ) );
  INVX8 U1 ( .A(n3), .Y(n1) );
  INVX8 U2 ( .A(n3), .Y(n2) );
  INVX8 U3 ( .A(S), .Y(n3) );
endmodule


module demux1to2_16_0 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), S, .Out0({\Out0<15> , \Out0<14> , 
        \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , \Out0<9> , \Out0<8> , 
        \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , \Out0<3> , \Out0<2> , 
        \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , \Out1<14> , \Out1<13> , 
        \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , \Out1<8> , \Out1<7> , 
        \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , \Out1<2> , \Out1<1> , 
        \Out1<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , S;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> ;
  wire   n1, n2;

  demux1to2_15 \d[0]  ( .In(\In<0> ), .S(n1), .Out0(\Out0<0> ), .Out1(
        \Out1<0> ) );
  demux1to2_14 \d[1]  ( .In(\In<1> ), .S(n1), .Out0(\Out0<1> ), .Out1(
        \Out1<1> ) );
  demux1to2_13 \d[2]  ( .In(\In<2> ), .S(n1), .Out0(\Out0<2> ), .Out1(
        \Out1<2> ) );
  demux1to2_12 \d[3]  ( .In(\In<3> ), .S(n1), .Out0(\Out0<3> ), .Out1(
        \Out1<3> ) );
  demux1to2_11 \d[4]  ( .In(\In<4> ), .S(n1), .Out0(\Out0<4> ), .Out1(
        \Out1<4> ) );
  demux1to2_10 \d[5]  ( .In(\In<5> ), .S(n1), .Out0(\Out0<5> ), .Out1(
        \Out1<5> ) );
  demux1to2_9 \d[6]  ( .In(\In<6> ), .S(n1), .Out0(\Out0<6> ), .Out1(\Out1<6> ) );
  demux1to2_8 \d[7]  ( .In(\In<7> ), .S(n1), .Out0(\Out0<7> ), .Out1(\Out1<7> ) );
  demux1to2_7 \d[8]  ( .In(\In<8> ), .S(n1), .Out0(\Out0<8> ), .Out1(\Out1<8> ) );
  demux1to2_6 \d[9]  ( .In(\In<9> ), .S(n1), .Out0(\Out0<9> ), .Out1(\Out1<9> ) );
  demux1to2_5 \d[10]  ( .In(\In<10> ), .S(n1), .Out0(\Out0<10> ), .Out1(
        \Out1<10> ) );
  demux1to2_4 \d[11]  ( .In(\In<11> ), .S(n1), .Out0(\Out0<11> ), .Out1(
        \Out1<11> ) );
  demux1to2_3 \d[12]  ( .In(\In<12> ), .S(n1), .Out0(\Out0<12> ), .Out1(
        \Out1<12> ) );
  demux1to2_2 \d[13]  ( .In(\In<13> ), .S(n1), .Out0(\Out0<13> ), .Out1(
        \Out1<13> ) );
  demux1to2_1 \d[14]  ( .In(\In<14> ), .S(n1), .Out0(\Out0<14> ), .Out1(
        \Out1<14> ) );
  demux1to2_0 \d[15]  ( .In(\In<15> ), .S(n1), .Out0(\Out0<15> ), .Out1(
        \Out1<15> ) );
  INVX4 U1 ( .A(S), .Y(n2) );
  INVX8 U2 ( .A(n2), .Y(n1) );
endmodule


module cla_or_xor_and ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , 
        \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , 
        \B<3> , \B<2> , \B<1> , \B<0> }), Cin, .Op({\Op<1> , \Op<0> }), .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<1> , \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Cout;
  wire   cla_cout, \op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> ,
         \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> ,
         \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> ,
         \op0_A<1> , \op0_A<0> , \op1_A<15> , \op1_A<14> , \op1_A<13> ,
         \op1_A<12> , \op1_A<11> , \op1_A<10> , \op1_A<9> , \op1_A<8> ,
         \op1_A<7> , \op1_A<6> , \op1_A<5> , \op1_A<4> , \op1_A<3> ,
         \op1_A<2> , \op1_A<1> , \op1_A<0> , \op2_A<15> , \op2_A<14> ,
         \op2_A<13> , \op2_A<12> , \op2_A<11> , \op2_A<10> , \op2_A<9> ,
         \op2_A<8> , \op2_A<7> , \op2_A<6> , \op2_A<5> , \op2_A<4> ,
         \op2_A<3> , \op2_A<2> , \op2_A<1> , \op2_A<0> , \op3_A<15> ,
         \op3_A<14> , \op3_A<13> , \op3_A<12> , \op3_A<11> , \op3_A<10> ,
         \op3_A<9> , \op3_A<8> , \op3_A<7> , \op3_A<6> , \op3_A<5> ,
         \op3_A<4> , \op3_A<3> , \op3_A<2> , \op3_A<1> , \op3_A<0> ,
         \op0_B<15> , \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> ,
         \op0_B<10> , \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> ,
         \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , \op0_B<1> ,
         \op0_B<0> , \op1_B<15> , \op1_B<14> , \op1_B<13> , \op1_B<12> ,
         \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , \op1_B<7> ,
         \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> ,
         \op1_B<1> , \op1_B<0> , \op2_B<15> , \op2_B<14> , \op2_B<13> ,
         \op2_B<12> , \op2_B<11> , \op2_B<10> , \op2_B<9> , \op2_B<8> ,
         \op2_B<7> , \op2_B<6> , \op2_B<5> , \op2_B<4> , \op2_B<3> ,
         \op2_B<2> , \op2_B<1> , \op2_B<0> , \op3_B<15> , \op3_B<14> ,
         \op3_B<13> , \op3_B<12> , \op3_B<11> , \op3_B<10> , \op3_B<9> ,
         \op3_B<8> , \op3_B<7> , \op3_B<6> , \op3_B<5> , \op3_B<4> ,
         \op3_B<3> , \op3_B<2> , \op3_B<1> , \op3_B<0> , \op0_out<15> ,
         \op0_out<14> , \op0_out<13> , \op0_out<12> , \op0_out<11> ,
         \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , \op0_out<6> ,
         \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , \op0_out<1> ,
         \op0_out<0> , \op1_out<13> , \op1_out<12> , \op1_out<11> ,
         \op1_out<10> , \op1_out<6> , \op1_out<5> , \op2_out<15> ,
         \op2_out<14> , \op2_out<13> , \op2_out<12> , \op2_out<11> ,
         \op2_out<10> , \op2_out<9> , \op2_out<8> , \op2_out<7> , \op2_out<6> ,
         \op2_out<5> , \op2_out<4> , \op2_out<3> , \op2_out<2> , \op2_out<1> ,
         \op2_out<0> , \op3_out<15> , \op3_out<14> , \op3_out<13> ,
         \op3_out<12> , \op3_out<11> , \op3_out<10> , \op3_out<9> ,
         \op3_out<8> , \op3_out<7> , \op3_out<6> , \op3_out<5> , \op3_out<4> ,
         \op3_out<3> , \op3_out<2> , \op3_out<1> , \op3_out<0> , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50;

  AND2X2 U15 ( .A(\op3_B<11> ), .B(\op3_A<11> ), .Y(\op3_out<11> ) );
  OR2X2 U29 ( .A(\op1_A<13> ), .B(\op1_B<13> ), .Y(\op1_out<13> ) );
  OR2X2 U30 ( .A(\op1_A<12> ), .B(\op1_B<12> ), .Y(\op1_out<12> ) );
  OR2X2 U31 ( .A(\op1_A<11> ), .B(\op1_B<11> ), .Y(\op1_out<11> ) );
  OR2X2 U32 ( .A(\op1_A<10> ), .B(\op1_B<10> ), .Y(\op1_out<10> ) );
  XOR2X1 U46 ( .A(\op2_B<13> ), .B(\op2_A<13> ), .Y(\op2_out<13> ) );
  XOR2X1 U47 ( .A(\op2_B<12> ), .B(\op2_A<12> ), .Y(\op2_out<12> ) );
  XOR2X1 U48 ( .A(\op2_B<11> ), .B(\op2_A<11> ), .Y(\op2_out<11> ) );
  XOR2X1 U49 ( .A(\op2_B<10> ), .B(\op2_A<10> ), .Y(\op2_out<10> ) );
  demux1to4_16_1 demux0 ( .In({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .S({\Op<1> , \Op<0> }), .Out0({\op0_A<15> , 
        \op0_A<14> , \op0_A<13> , \op0_A<12> , \op0_A<11> , \op0_A<10> , 
        \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , \op0_A<5> , \op0_A<4> , 
        \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .Out1({\op1_A<15> , 
        \op1_A<14> , \op1_A<13> , \op1_A<12> , \op1_A<11> , \op1_A<10> , 
        \op1_A<9> , \op1_A<8> , \op1_A<7> , \op1_A<6> , \op1_A<5> , \op1_A<4> , 
        \op1_A<3> , \op1_A<2> , \op1_A<1> , \op1_A<0> }), .Out2({\op2_A<15> , 
        \op2_A<14> , \op2_A<13> , \op2_A<12> , \op2_A<11> , \op2_A<10> , 
        \op2_A<9> , \op2_A<8> , \op2_A<7> , \op2_A<6> , \op2_A<5> , \op2_A<4> , 
        \op2_A<3> , \op2_A<2> , \op2_A<1> , \op2_A<0> }), .Out3({\op3_A<15> , 
        \op3_A<14> , \op3_A<13> , \op3_A<12> , \op3_A<11> , \op3_A<10> , 
        \op3_A<9> , \op3_A<8> , \op3_A<7> , \op3_A<6> , \op3_A<5> , \op3_A<4> , 
        \op3_A<3> , \op3_A<2> , \op3_A<1> , \op3_A<0> }) );
  demux1to4_16_0 demux1 ( .In({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , 
        \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , 
        \B<2> , \B<1> , \B<0> }), .S({\Op<1> , \Op<0> }), .Out0({\op0_B<15> , 
        \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , \op0_B<10> , 
        \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , 
        \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }), .Out1({\op1_B<15> , 
        \op1_B<14> , \op1_B<13> , \op1_B<12> , \op1_B<11> , \op1_B<10> , 
        \op1_B<9> , \op1_B<8> , \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , 
        \op1_B<3> , \op1_B<2> , \op1_B<1> , \op1_B<0> }), .Out2({\op2_B<15> , 
        \op2_B<14> , \op2_B<13> , \op2_B<12> , \op2_B<11> , \op2_B<10> , 
        \op2_B<9> , \op2_B<8> , \op2_B<7> , \op2_B<6> , \op2_B<5> , \op2_B<4> , 
        \op2_B<3> , \op2_B<2> , \op2_B<1> , \op2_B<0> }), .Out3({\op3_B<15> , 
        \op3_B<14> , \op3_B<13> , \op3_B<12> , \op3_B<11> , \op3_B<10> , 
        \op3_B<9> , \op3_B<8> , \op3_B<7> , \op3_B<6> , \op3_B<5> , \op3_B<4> , 
        \op3_B<3> , \op3_B<2> , \op3_B<1> , \op3_B<0> }) );
  cla16_0 cla0 ( .A({\op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> , 
        \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> , 
        \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> , \op0_A<1> , 
        \op0_A<0> }), .B({\op0_B<15> , \op0_B<14> , \op0_B<13> , \op0_B<12> , 
        \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> , \op0_B<7> , 
        \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , \op0_B<1> , 
        \op0_B<0> }), .Cin(Cin), .S({\op0_out<15> , \op0_out<14> , 
        \op0_out<13> , \op0_out<12> , \op0_out<11> , \op0_out<10> , 
        \op0_out<9> , \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , 
        \op0_out<4> , \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> }), 
        .Cout(cla_cout) );
  mux4to1_16_4 mux0 ( .InA({\op0_out<15> , \op0_out<14> , \op0_out<13> , 
        \op0_out<12> , \op0_out<11> , \op0_out<10> , \op0_out<9> , 
        \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , \op0_out<4> , 
        \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> }), .InB({n2, 
        n12, \op1_out<13> , \op1_out<12> , \op1_out<11> , \op1_out<10> , n10, 
        n20, n18, \op1_out<6> , \op1_out<5> , n16, n8, n14, n6, n4}), .InC({
        \op2_out<15> , \op2_out<14> , \op2_out<13> , \op2_out<12> , 
        \op2_out<11> , \op2_out<10> , \op2_out<9> , \op2_out<8> , \op2_out<7> , 
        \op2_out<6> , \op2_out<5> , \op2_out<4> , \op2_out<3> , \op2_out<2> , 
        \op2_out<1> , \op2_out<0> }), .InD({\op3_out<15> , \op3_out<14> , 
        \op3_out<13> , \op3_out<12> , \op3_out<11> , \op3_out<10> , 
        \op3_out<9> , \op3_out<8> , \op3_out<7> , \op3_out<6> , \op3_out<5> , 
        \op3_out<4> , \op3_out<3> , \op3_out<2> , \op3_out<1> , \op3_out<0> }), 
        .S({n22, n21}), .Out({\Out<15> , \Out<14> , \Out<13> , \Out<12> , 
        \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , 
        \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> }) );
  AND2X1 U2 ( .A(\op3_B<12> ), .B(\op3_A<12> ), .Y(\op3_out<12> ) );
  INVX1 U3 ( .A(\op1_A<7> ), .Y(n40) );
  AND2X1 U4 ( .A(\op3_B<10> ), .B(\op3_A<10> ), .Y(\op3_out<10> ) );
  AND2X1 U5 ( .A(\op3_B<13> ), .B(\op3_A<13> ), .Y(\op3_out<13> ) );
  OR2X1 U6 ( .A(\op1_A<6> ), .B(\op1_B<6> ), .Y(\op1_out<6> ) );
  AND2X2 U7 ( .A(n49), .B(n48), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(n2) );
  OR2X1 U9 ( .A(\op1_A<5> ), .B(\op1_B<5> ), .Y(\op1_out<5> ) );
  AND2X1 U10 ( .A(\op3_B<5> ), .B(\op3_A<5> ), .Y(\op3_out<5> ) );
  AND2X1 U11 ( .A(n31), .B(n30), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(n4) );
  AND2X1 U13 ( .A(n33), .B(n32), .Y(n5) );
  INVX1 U14 ( .A(n5), .Y(n6) );
  AND2X1 U16 ( .A(n37), .B(n36), .Y(n7) );
  INVX1 U17 ( .A(n7), .Y(n8) );
  AND2X1 U18 ( .A(n45), .B(n44), .Y(n9) );
  INVX1 U19 ( .A(n9), .Y(n10) );
  AND2X1 U20 ( .A(n47), .B(n46), .Y(n11) );
  INVX1 U21 ( .A(n11), .Y(n12) );
  INVX1 U22 ( .A(cla_cout), .Y(n50) );
  INVX1 U23 ( .A(\op1_B<15> ), .Y(n49) );
  INVX1 U24 ( .A(\op1_B<14> ), .Y(n47) );
  INVX1 U25 ( .A(\op1_B<9> ), .Y(n45) );
  INVX1 U26 ( .A(\op1_B<8> ), .Y(n43) );
  INVX1 U27 ( .A(\op1_B<7> ), .Y(n41) );
  INVX1 U28 ( .A(\op1_B<4> ), .Y(n39) );
  INVX1 U33 ( .A(\op1_B<3> ), .Y(n37) );
  INVX1 U34 ( .A(\op1_B<2> ), .Y(n35) );
  INVX1 U35 ( .A(\op1_B<1> ), .Y(n33) );
  INVX1 U36 ( .A(\op1_B<0> ), .Y(n31) );
  INVX1 U37 ( .A(\op2_A<15> ), .Y(n29) );
  INVX1 U38 ( .A(\op2_A<14> ), .Y(n28) );
  INVX1 U39 ( .A(\op2_A<8> ), .Y(n27) );
  INVX1 U40 ( .A(\op2_A<4> ), .Y(n26) );
  AND2X1 U41 ( .A(n35), .B(n34), .Y(n13) );
  INVX1 U42 ( .A(n13), .Y(n14) );
  AND2X1 U43 ( .A(n39), .B(n38), .Y(n15) );
  INVX1 U44 ( .A(n15), .Y(n16) );
  AND2X1 U45 ( .A(n41), .B(n40), .Y(n17) );
  INVX1 U50 ( .A(n17), .Y(n18) );
  AND2X1 U51 ( .A(n43), .B(n42), .Y(n19) );
  INVX1 U52 ( .A(n19), .Y(n20) );
  INVX1 U53 ( .A(n23), .Y(n22) );
  BUFX2 U54 ( .A(\Op<0> ), .Y(n21) );
  INVX1 U55 ( .A(\Op<1> ), .Y(n23) );
  AND2X2 U56 ( .A(\op3_A<0> ), .B(\op3_B<0> ), .Y(\op3_out<0> ) );
  AND2X2 U57 ( .A(\op3_A<1> ), .B(\op3_B<1> ), .Y(\op3_out<1> ) );
  AND2X2 U58 ( .A(\op3_A<2> ), .B(\op3_B<2> ), .Y(\op3_out<2> ) );
  AND2X2 U59 ( .A(\op3_A<3> ), .B(\op3_B<3> ), .Y(\op3_out<3> ) );
  AND2X2 U60 ( .A(\op3_A<4> ), .B(\op3_B<4> ), .Y(\op3_out<4> ) );
  AND2X2 U61 ( .A(\op3_A<6> ), .B(\op3_B<6> ), .Y(\op3_out<6> ) );
  AND2X2 U62 ( .A(\op3_A<7> ), .B(\op3_B<7> ), .Y(\op3_out<7> ) );
  AND2X2 U63 ( .A(\op3_A<8> ), .B(\op3_B<8> ), .Y(\op3_out<8> ) );
  AND2X2 U64 ( .A(\op3_A<9> ), .B(\op3_B<9> ), .Y(\op3_out<9> ) );
  AND2X2 U65 ( .A(\op3_A<14> ), .B(\op3_B<14> ), .Y(\op3_out<14> ) );
  AND2X2 U66 ( .A(\op3_A<15> ), .B(\op3_B<15> ), .Y(\op3_out<15> ) );
  XOR2X1 U67 ( .A(\op2_A<0> ), .B(\op2_B<0> ), .Y(\op2_out<0> ) );
  INVX2 U68 ( .A(\op2_A<1> ), .Y(n24) );
  XNOR2X1 U69 ( .A(\op2_B<1> ), .B(n24), .Y(\op2_out<1> ) );
  INVX2 U70 ( .A(\op2_A<2> ), .Y(n25) );
  XNOR2X1 U71 ( .A(\op2_B<2> ), .B(n25), .Y(\op2_out<2> ) );
  XOR2X1 U72 ( .A(\op2_A<3> ), .B(\op2_B<3> ), .Y(\op2_out<3> ) );
  XNOR2X1 U73 ( .A(\op2_B<4> ), .B(n26), .Y(\op2_out<4> ) );
  XOR2X1 U74 ( .A(\op2_A<5> ), .B(\op2_B<5> ), .Y(\op2_out<5> ) );
  XOR2X1 U75 ( .A(\op2_A<6> ), .B(\op2_B<6> ), .Y(\op2_out<6> ) );
  XOR2X1 U76 ( .A(\op2_A<7> ), .B(\op2_B<7> ), .Y(\op2_out<7> ) );
  XNOR2X1 U77 ( .A(\op2_B<8> ), .B(n27), .Y(\op2_out<8> ) );
  XOR2X1 U78 ( .A(\op2_A<9> ), .B(\op2_B<9> ), .Y(\op2_out<9> ) );
  XNOR2X1 U79 ( .A(\op2_B<14> ), .B(n28), .Y(\op2_out<14> ) );
  XNOR2X1 U80 ( .A(\op2_B<15> ), .B(n29), .Y(\op2_out<15> ) );
  INVX2 U81 ( .A(\op1_A<0> ), .Y(n30) );
  INVX2 U82 ( .A(\op1_A<1> ), .Y(n32) );
  INVX2 U83 ( .A(\op1_A<2> ), .Y(n34) );
  INVX2 U84 ( .A(\op1_A<3> ), .Y(n36) );
  INVX2 U85 ( .A(\op1_A<4> ), .Y(n38) );
  INVX2 U86 ( .A(\op1_A<8> ), .Y(n42) );
  INVX2 U87 ( .A(\op1_A<9> ), .Y(n44) );
  INVX2 U88 ( .A(\op1_A<14> ), .Y(n46) );
  INVX2 U89 ( .A(\op1_A<15> ), .Y(n48) );
  NOR3X1 U90 ( .A(n22), .B(n21), .C(n50), .Y(Cout) );
endmodule


module shifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Op({\Op<1> , \Op<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , \Op<1> ,
         \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \ls_out<15> , \ls_out<14> , \ls_out<13> , \ls_out<12> , \ls_out<11> ,
         \ls_out<10> , \ls_out<9> , \ls_out<8> , \ls_out<7> , \ls_out<6> ,
         \ls_out<5> , \ls_out<4> , \ls_out<3> , \ls_out<2> , \ls_out<1> ,
         \ls_out<0> , \rs_out<15> , \rs_out<14> , \rs_out<13> , \rs_out<12> ,
         \rs_out<11> , \rs_out<10> , \rs_out<9> , \rs_out<8> , \rs_out<7> ,
         \rs_out<6> , \rs_out<5> , \rs_out<4> , \rs_out<3> , \rs_out<2> ,
         \rs_out<1> , \rs_out<0> , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38;

  lshifter ls ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Rot_sel(n6), .Out({\ls_out<15> , \ls_out<14> , 
        \ls_out<13> , \ls_out<12> , \ls_out<11> , \ls_out<10> , \ls_out<9> , 
        \ls_out<8> , \ls_out<7> , \ls_out<6> , \ls_out<5> , \ls_out<4> , 
        \ls_out<3> , \ls_out<2> , \ls_out<1> , \ls_out<0> }) );
  rshifter rs ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Rot_sel(n6), .Out({\rs_out<15> , \rs_out<14> , 
        \rs_out<13> , \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> , 
        \rs_out<8> , \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> , 
        \rs_out<3> , \rs_out<2> , \rs_out<1> , \rs_out<0> }) );
  INVX1 U1 ( .A(n9), .Y(n7) );
  INVX1 U2 ( .A(n1), .Y(\Out<0> ) );
  MUX2X1 U3 ( .B(\rs_out<0> ), .A(\ls_out<0> ), .S(n9), .Y(n1) );
  AND2X2 U4 ( .A(n4), .B(n5), .Y(\Out<1> ) );
  BUFX2 U5 ( .A(\rs_out<1> ), .Y(n3) );
  INVX1 U6 ( .A(\rs_out<9> ), .Y(n25) );
  INVX1 U7 ( .A(\rs_out<10> ), .Y(n27) );
  INVX1 U8 ( .A(\rs_out<11> ), .Y(n29) );
  INVX1 U9 ( .A(\rs_out<13> ), .Y(n33) );
  INVX1 U10 ( .A(\rs_out<14> ), .Y(n35) );
  INVX1 U11 ( .A(\rs_out<15> ), .Y(n37) );
  INVX1 U12 ( .A(\ls_out<6> ), .Y(n20) );
  INVX1 U13 ( .A(\ls_out<9> ), .Y(n26) );
  INVX1 U14 ( .A(\ls_out<10> ), .Y(n28) );
  INVX1 U15 ( .A(\ls_out<13> ), .Y(n34) );
  INVX1 U16 ( .A(\ls_out<14> ), .Y(n36) );
  INVX1 U17 ( .A(\rs_out<6> ), .Y(n19) );
  INVX1 U18 ( .A(\rs_out<7> ), .Y(n21) );
  INVX1 U19 ( .A(\rs_out<8> ), .Y(n23) );
  INVX1 U20 ( .A(\rs_out<12> ), .Y(n31) );
  INVX1 U21 ( .A(\ls_out<7> ), .Y(n22) );
  INVX1 U22 ( .A(\ls_out<8> ), .Y(n24) );
  INVX1 U23 ( .A(\ls_out<11> ), .Y(n30) );
  INVX1 U24 ( .A(\ls_out<12> ), .Y(n32) );
  INVX1 U25 ( .A(\ls_out<15> ), .Y(n38) );
  INVX1 U26 ( .A(\ls_out<2> ), .Y(n12) );
  INVX1 U27 ( .A(\rs_out<3> ), .Y(n13) );
  INVX1 U28 ( .A(\ls_out<3> ), .Y(n14) );
  OR2X2 U29 ( .A(n3), .B(n9), .Y(n5) );
  INVX1 U30 ( .A(\rs_out<4> ), .Y(n15) );
  NAND2X1 U31 ( .A(n10), .B(n9), .Y(n4) );
  INVX1 U32 ( .A(n9), .Y(n8) );
  INVX1 U33 ( .A(\ls_out<4> ), .Y(n16) );
  INVX1 U34 ( .A(\ls_out<5> ), .Y(n18) );
  INVX1 U35 ( .A(\rs_out<5> ), .Y(n17) );
  INVX1 U36 ( .A(\ls_out<1> ), .Y(n10) );
  INVX1 U37 ( .A(\rs_out<2> ), .Y(n11) );
  INVX1 U38 ( .A(\Op<1> ), .Y(n9) );
  INVX8 U39 ( .A(\Op<0> ), .Y(n6) );
  MUX2X1 U40 ( .B(n12), .A(n11), .S(n8), .Y(\Out<2> ) );
  MUX2X1 U41 ( .B(n14), .A(n13), .S(n8), .Y(\Out<3> ) );
  MUX2X1 U42 ( .B(n16), .A(n15), .S(n7), .Y(\Out<4> ) );
  MUX2X1 U43 ( .B(n18), .A(n17), .S(n7), .Y(\Out<5> ) );
  MUX2X1 U44 ( .B(n20), .A(n19), .S(n7), .Y(\Out<6> ) );
  MUX2X1 U45 ( .B(n22), .A(n21), .S(n7), .Y(\Out<7> ) );
  MUX2X1 U46 ( .B(n24), .A(n23), .S(n7), .Y(\Out<8> ) );
  MUX2X1 U47 ( .B(n26), .A(n25), .S(n7), .Y(\Out<9> ) );
  MUX2X1 U48 ( .B(n28), .A(n27), .S(n7), .Y(\Out<10> ) );
  MUX2X1 U49 ( .B(n30), .A(n29), .S(n7), .Y(\Out<11> ) );
  MUX2X1 U50 ( .B(n32), .A(n31), .S(n7), .Y(\Out<12> ) );
  MUX2X1 U51 ( .B(n34), .A(n33), .S(n7), .Y(\Out<13> ) );
  MUX2X1 U52 ( .B(n36), .A(n35), .S(n7), .Y(\Out<14> ) );
  MUX2X1 U53 ( .B(n38), .A(n37), .S(n7), .Y(\Out<15> ) );
endmodule


module cla4_7 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n19), .C(n21), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n21), .C(n20), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n18), .C(\G<2> ), .Y(n41) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n40) );
  OAI21X1 U13 ( .A(n9), .B(n21), .C(n20), .Y(Cout) );
  AOI21X1 U14 ( .A(n16), .B(\P<2> ), .C(\G<2> ), .Y(n39) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n38) );
  fulladder1_31 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_30 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_29 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n16), .S(\S<2> ), .P(
        n35), .G(n27) );
  fulladder1_28 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  INVX1 U1 ( .A(\P<2> ), .Y(n19) );
  AND2X1 U2 ( .A(n17), .B(n2), .Y(n10) );
  INVX1 U3 ( .A(\G<0> ), .Y(n17) );
  INVX1 U4 ( .A(\G<3> ), .Y(n20) );
  INVX1 U5 ( .A(\P<3> ), .Y(n21) );
  AND2X1 U6 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  BUFX2 U9 ( .A(n38), .Y(n3) );
  INVX1 U16 ( .A(n3), .Y(n16) );
  INVX1 U17 ( .A(n41), .Y(n4) );
  INVX1 U18 ( .A(n4), .Y(n5) );
  INVX1 U19 ( .A(n40), .Y(n18) );
  AND2X1 U20 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U21 ( .A(n6), .Y(n7) );
  INVX1 U22 ( .A(n9), .Y(n8) );
  BUFX2 U23 ( .A(n39), .Y(n9) );
  INVX1 U24 ( .A(n10), .Y(n12) );
  AND2X1 U25 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U26 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U27 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U28 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U29 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U30 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U31 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U32 ( .A(n22), .B(n23), .Y(\G<0> ) );
endmodule


module cla4_6 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n7), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n9), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_27 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_26 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_25 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_24 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n38), .G(n30) );
  INVX1 U1 ( .A(\P<2> ), .Y(n20) );
  INVX1 U2 ( .A(\G<0> ), .Y(n18) );
  INVX1 U3 ( .A(\G<3> ), .Y(n21) );
  INVX1 U4 ( .A(\P<3> ), .Y(n22) );
  AND2X1 U5 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  BUFX2 U7 ( .A(n39), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(n17) );
  BUFX2 U16 ( .A(n41), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n19) );
  BUFX2 U18 ( .A(n42), .Y(n5) );
  AND2X1 U19 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(n7) );
  INVX1 U21 ( .A(n10), .Y(n8) );
  INVX1 U22 ( .A(n8), .Y(n9) );
  BUFX2 U23 ( .A(n40), .Y(n10) );
  AND2X2 U24 ( .A(n18), .B(n2), .Y(n12) );
  INVX1 U25 ( .A(n12), .Y(n16) );
  AND2X1 U26 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U27 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U28 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U29 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U30 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U31 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U32 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U33 ( .A(n23), .B(n24), .Y(\G<0> ) );
endmodule


module cla4_5 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n7), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n9), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_23 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_22 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_21 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_20 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n38), .G(n30) );
  INVX1 U1 ( .A(\G<0> ), .Y(n18) );
  INVX1 U2 ( .A(\P<2> ), .Y(n20) );
  INVX1 U3 ( .A(\G<3> ), .Y(n21) );
  INVX1 U4 ( .A(\P<3> ), .Y(n22) );
  AND2X1 U5 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  BUFX2 U7 ( .A(n39), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(n17) );
  BUFX2 U16 ( .A(n41), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n19) );
  BUFX2 U18 ( .A(n42), .Y(n5) );
  AND2X1 U19 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(n7) );
  INVX1 U21 ( .A(n10), .Y(n8) );
  INVX1 U22 ( .A(n8), .Y(n9) );
  BUFX2 U23 ( .A(n40), .Y(n10) );
  AND2X2 U24 ( .A(n18), .B(n2), .Y(n12) );
  INVX1 U25 ( .A(n12), .Y(n16) );
  AND2X1 U26 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U27 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U28 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U29 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U30 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U31 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U32 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U33 ( .A(n23), .B(n24), .Y(\G<0> ) );
endmodule


module cla4_4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n19), .C(n21), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n21), .C(n20), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n18), .C(\G<2> ), .Y(n41) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n40) );
  OAI21X1 U13 ( .A(n9), .B(n21), .C(n20), .Y(Cout) );
  AOI21X1 U14 ( .A(n16), .B(\P<2> ), .C(\G<2> ), .Y(n39) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n38) );
  fulladder1_19 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_18 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_17 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n3), .S(\S<2> ), .P(n35), .G(n27) );
  fulladder1_16 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  INVX1 U1 ( .A(\G<0> ), .Y(n17) );
  INVX1 U2 ( .A(\P<2> ), .Y(n19) );
  INVX1 U3 ( .A(\G<3> ), .Y(n20) );
  INVX1 U4 ( .A(\P<3> ), .Y(n21) );
  AND2X1 U5 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  BUFX2 U7 ( .A(n16), .Y(n3) );
  INVX1 U9 ( .A(n38), .Y(n16) );
  BUFX2 U16 ( .A(n40), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n18) );
  BUFX2 U18 ( .A(n41), .Y(n5) );
  AND2X1 U19 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(n7) );
  INVX1 U21 ( .A(n39), .Y(n8) );
  INVX1 U22 ( .A(n8), .Y(n9) );
  AND2X2 U23 ( .A(n17), .B(n2), .Y(n10) );
  INVX1 U24 ( .A(n10), .Y(n12) );
  AND2X1 U25 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U26 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U27 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U28 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U29 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U30 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U31 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U32 ( .A(n22), .B(n23), .Y(\G<0> ) );
endmodule


module dff_388 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_389 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_390 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_391 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_392 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_393 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_394 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_395 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_396 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_397 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_398 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_399 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_400 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_401 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_402 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_403 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_372 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_373 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_374 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_375 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_376 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_377 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_378 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_379 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_380 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_381 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_382 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_383 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_384 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_385 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_386 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_387 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_404 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memory2c ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, \mem<0><7> , \mem<0><6> , \mem<0><5> ,
         \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> ,
         \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> ,
         \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> ,
         \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> ,
         \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> ,
         \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> ,
         \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> ,
         \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> ,
         \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> ,
         \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> ,
         \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> ,
         \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> ,
         \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> ,
         \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> ,
         \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> ,
         \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> ,
         \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> ,
         \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> ,
         \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> ,
         \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> ,
         \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> ,
         \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> ,
         \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> ,
         \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> ,
         \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> ,
         \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> ,
         \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> ,
         \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> ,
         \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> ,
         \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> ,
         \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> ,
         \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> ,
         \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> ,
         \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> ,
         \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> ,
         \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> ,
         \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> ,
         \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> ,
         \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> , \mem<33><4> ,
         \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> , \mem<34><7> ,
         \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> , \mem<34><2> ,
         \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> , \mem<35><5> ,
         \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> , \mem<35><0> ,
         \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> , \mem<36><3> ,
         \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> , \mem<37><6> ,
         \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> , \mem<37><1> ,
         \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> , \mem<38><4> ,
         \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> , \mem<39><7> ,
         \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> , \mem<39><2> ,
         \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> , \mem<40><5> ,
         \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> , \mem<40><0> ,
         \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> , \mem<41><3> ,
         \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> , \mem<42><6> ,
         \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> , \mem<42><1> ,
         \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> , \mem<43><4> ,
         \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> , \mem<44><7> ,
         \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> , \mem<44><2> ,
         \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> , \mem<45><5> ,
         \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> , \mem<45><0> ,
         \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> , \mem<46><3> ,
         \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> , \mem<47><6> ,
         \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> , \mem<47><1> ,
         \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> , \mem<48><4> ,
         \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> , \mem<49><7> ,
         \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> , \mem<49><2> ,
         \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> , \mem<50><5> ,
         \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> , \mem<50><0> ,
         \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> , \mem<51><3> ,
         \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> , \mem<52><6> ,
         \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> , \mem<52><1> ,
         \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> , \mem<53><4> ,
         \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> , \mem<54><7> ,
         \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> , \mem<54><2> ,
         \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> , \mem<55><5> ,
         \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> , \mem<55><0> ,
         \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> , \mem<56><3> ,
         \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> , \mem<57><6> ,
         \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> , \mem<57><1> ,
         \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> , \mem<58><4> ,
         \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> , \mem<59><7> ,
         \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> , \mem<59><2> ,
         \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> , \mem<60><5> ,
         \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> , \mem<60><0> ,
         \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> , \mem<61><3> ,
         \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> , \mem<62><6> ,
         \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> , \mem<62><1> ,
         \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> , \mem<63><4> ,
         \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> , N185, N186,
         N187, N188, N189, N190, N191, N192, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n610, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1367, n1368,
         n1370, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1772, n1774, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1797,
         n1798, n1799, n1800, n1801, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n609, n611, n624, n637, n649, n661, n673, n685, n697,
         n709, n721, n733, n745, n757, n769, n781, n793, n805, n817, n829,
         n841, n853, n865, n877, n889, n901, n913, n925, n937, n949, n961,
         n973, n985, n997, n1009, n1021, n1033, n1045, n1057, n1069, n1081,
         n1093, n1105, n1117, n1129, n1141, n1153, n1165, n1177, n1189, n1201,
         n1213, n1225, n1237, n1249, n1261, n1273, n1285, n1297, n1309, n1321,
         n1333, n1345, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1369, n1371, n1372, n1383, n1384, n1396, n1397, n1409,
         n1410, n1424, n1425, n1436, n1437, n1449, n1450, n1461, n1462, n1476,
         n1477, n1488, n1489, n1501, n1502, n1513, n1514, n1528, n1529, n1540,
         n1541, n1553, n1554, n1565, n1566, n1580, n1581, n1592, n1593, n1605,
         n1606, n1617, n1618, n1632, n1633, n1644, n1645, n1657, n1658, n1669,
         n1670, n1684, n1685, n1696, n1697, n1709, n1710, n1721, n1722, n1736,
         n1737, n1758, n1759, n1771, n1773, n1775, n1776, n1793, n1794, n1795,
         n1796, n1802, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n2327), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2326), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2325), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2324), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2323), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2322), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2321), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2320), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2319), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2318), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2317), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2316), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2315), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2314), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2313), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2312), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2311), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2310), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2309), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2308), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2307), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2306), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2305), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2304), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2303), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2302), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2301), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2300), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2299), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2298), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2297), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2296), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2295), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2294), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2293), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2292), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2291), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2290), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2289), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2288), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2287), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2286), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2285), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2284), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2283), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2282), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2281), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2280), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2279), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2278), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2277), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2276), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2275), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2274), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2273), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2272), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2271), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2270), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2269), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2268), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2267), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2266), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2265), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2264), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2263), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2262), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2261), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2260), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2259), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2258), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2257), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2256), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2255), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2254), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2253), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2252), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2251), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2250), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2249), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2248), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2247), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2246), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2245), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2244), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2243), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2242), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2241), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2240), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2239), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2238), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2237), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2236), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2235), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2234), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2233), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2232), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2231), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2230), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2229), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2228), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2227), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2226), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2225), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2224), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2223), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2222), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2221), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2220), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2219), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2218), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2217), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2216), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2215), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2214), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2213), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2212), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2211), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2210), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2209), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2208), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2207), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2206), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2205), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2204), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2203), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2202), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2201), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2200), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2199), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2198), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2197), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2196), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2195), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2194), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2193), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2192), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2191), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2190), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2189), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2188), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2187), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2186), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2185), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2184), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2183), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2182), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2181), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2180), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2179), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2178), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2177), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2176), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2175), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2174), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2173), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2172), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2171), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2170), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2169), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2168), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2167), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2166), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2165), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2164), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2163), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2162), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2161), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2160), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2159), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2158), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2157), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2156), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2155), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2154), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2153), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2152), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2151), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2150), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2149), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2148), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2147), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2146), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2145), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2144), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2143), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2142), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2141), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2140), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2139), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2138), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2137), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2136), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2135), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2134), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2133), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2132), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2131), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2130), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2129), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2128), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2127), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2126), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2125), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2124), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2123), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2122), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2121), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2120), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2119), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2118), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2117), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2116), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2115), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2114), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2113), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2112), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2111), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2110), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2109), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2108), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2107), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2106), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2105), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2104), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2103), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2102), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2101), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2100), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2099), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2098), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2097), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2096), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2095), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2094), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2093), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2092), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2091), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2090), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2089), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2088), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2087), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2086), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2085), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2084), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2083), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2082), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2081), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2080), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2079), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2078), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2077), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2076), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2075), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2074), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2073), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2072), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n2071), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n2070), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n2069), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n2068), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n2067), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n2066), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n2065), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n2064), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n2063), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n2062), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n2061), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n2060), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n2059), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n2058), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n2057), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n2056), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n2055), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n2054), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n2053), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n2052), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n2051), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n2050), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n2049), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n2048), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n2047), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n2046), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n2045), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n2044), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n2043), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n2042), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n2041), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n2040), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n2039), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n2038), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n2037), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n2036), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n2035), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n2034), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n2033), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n2032), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n2031), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n2030), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n2029), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n2028), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n2027), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n2026), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n2025), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n2024), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n2023), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n2022), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n2021), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n2020), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n2019), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n2018), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n2017), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n2016), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n2015), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n2014), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n2013), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n2012), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n2011), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n2010), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n2009), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n2008), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n2007), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n2006), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n2005), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n2004), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n2003), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n2002), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n2001), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n2000), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n1999), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n1998), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n1997), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n1996), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n1995), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n1994), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n1993), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n1992), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n1991), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n1990), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n1989), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n1988), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n1987), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n1986), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n1985), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n1984), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n1983), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n1982), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n1981), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n1980), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n1979), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n1978), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n1977), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n1976), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n1975), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n1974), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n1973), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n1972), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n1971), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n1970), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n1969), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n1968), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n1967), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n1966), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n1965), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n1964), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n1963), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n1962), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n1961), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n1960), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n1959), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n1958), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n1957), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n1956), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n1955), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n1954), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n1953), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n1952), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n1951), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n1950), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n1949), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n1948), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n1947), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n1946), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n1945), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n1944), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n1943), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n1942), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n1941), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n1940), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n1939), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n1938), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n1937), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n1936), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n1935), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n1934), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n1933), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n1932), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n1931), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n1930), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n1929), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n1928), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n1927), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n1926), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n1925), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n1924), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n1923), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n1922), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n1921), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n1920), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n1919), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n1918), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n1917), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n1916), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n1915), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n1914), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n1913), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n1912), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n1911), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n1910), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n1909), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n1908), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n1907), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n1906), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n1905), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n1904), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n1903), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n1902), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n1901), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n1900), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n1899), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n1898), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n1897), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n1896), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n1895), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n1894), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n1893), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n1892), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n1891), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n1890), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n1889), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n1888), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n1887), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n1886), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n1885), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n1884), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n1883), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n1882), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n1881), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n1880), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n1879), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n1878), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n1877), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n1876), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n1875), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n1874), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n1873), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n1872), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n1871), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n1870), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n1869), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n1868), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n1867), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n1866), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n1865), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n1864), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n1863), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n1862), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n1861), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n1860), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n1859), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n1858), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n1857), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n1856), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n1855), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n1854), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n1853), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n1852), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n1851), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n1850), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n1849), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n1848), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n1847), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n1846), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n1845), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n1844), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n1843), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n1842), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n1841), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n1840), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n1839), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n1838), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n1837), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n1836), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n1835), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n1834), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n1833), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n1832), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n1831), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n1830), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n1829), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n1828), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n1827), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n1826), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n1825), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n1824), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n1823), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n1822), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n1821), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n1820), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n1819), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n1818), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n1817), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n1816), .CLK(clk), .Q(\mem<63><0> ) );
  AND2X2 U132 ( .A(n1376), .B(n1377), .Y(n1375) );
  AND2X2 U133 ( .A(n1381), .B(n1382), .Y(n1380) );
  AND2X2 U135 ( .A(n1388), .B(n1389), .Y(n1387) );
  AND2X2 U136 ( .A(n1393), .B(n1394), .Y(n1392) );
  AND2X2 U137 ( .A(n1401), .B(n1402), .Y(n1400) );
  AND2X2 U138 ( .A(n1407), .B(n1408), .Y(n1406) );
  AND2X2 U140 ( .A(n1414), .B(n1415), .Y(n1413) );
  AND2X2 U141 ( .A(n1419), .B(n1420), .Y(n1418) );
  AND2X2 U142 ( .A(n1429), .B(n1430), .Y(n1428) );
  AND2X2 U143 ( .A(n1434), .B(n1435), .Y(n1433) );
  AND2X2 U145 ( .A(n1441), .B(n1442), .Y(n1440) );
  AND2X2 U146 ( .A(n1446), .B(n1447), .Y(n1445) );
  AND2X2 U147 ( .A(n1454), .B(n1455), .Y(n1453) );
  AND2X2 U148 ( .A(n1459), .B(n1460), .Y(n1458) );
  AND2X2 U150 ( .A(n1466), .B(n1467), .Y(n1465) );
  AND2X2 U151 ( .A(n1471), .B(n1472), .Y(n1470) );
  AND2X2 U152 ( .A(n1481), .B(n1482), .Y(n1480) );
  AND2X2 U153 ( .A(n1486), .B(n1487), .Y(n1485) );
  AND2X2 U155 ( .A(n1493), .B(n1494), .Y(n1492) );
  AND2X2 U156 ( .A(n1498), .B(n1499), .Y(n1497) );
  AND2X2 U157 ( .A(n1506), .B(n1507), .Y(n1505) );
  AND2X2 U158 ( .A(n1511), .B(n1512), .Y(n1510) );
  AND2X2 U160 ( .A(n1518), .B(n1519), .Y(n1517) );
  AND2X2 U161 ( .A(n1523), .B(n1524), .Y(n1522) );
  AND2X2 U162 ( .A(n1533), .B(n1534), .Y(n1532) );
  AND2X2 U163 ( .A(n1538), .B(n1539), .Y(n1537) );
  AND2X2 U165 ( .A(n1545), .B(n1546), .Y(n1544) );
  AND2X2 U166 ( .A(n1550), .B(n1551), .Y(n1549) );
  AND2X2 U167 ( .A(n1558), .B(n1559), .Y(n1557) );
  AND2X2 U168 ( .A(n1563), .B(n1564), .Y(n1562) );
  AND2X2 U170 ( .A(n1570), .B(n1571), .Y(n1569) );
  AND2X2 U171 ( .A(n1575), .B(n1576), .Y(n1574) );
  AND2X2 U172 ( .A(n1585), .B(n1586), .Y(n1584) );
  AND2X2 U173 ( .A(n1590), .B(n1591), .Y(n1589) );
  AND2X2 U175 ( .A(n1597), .B(n1598), .Y(n1596) );
  AND2X2 U176 ( .A(n1602), .B(n1603), .Y(n1601) );
  AND2X2 U177 ( .A(n1610), .B(n1611), .Y(n1609) );
  AND2X2 U178 ( .A(n1615), .B(n1616), .Y(n1614) );
  AND2X2 U180 ( .A(n1622), .B(n1623), .Y(n1621) );
  AND2X2 U181 ( .A(n1627), .B(n1628), .Y(n1626) );
  AND2X2 U182 ( .A(n1637), .B(n1638), .Y(n1636) );
  AND2X2 U183 ( .A(n1642), .B(n1643), .Y(n1641) );
  AND2X2 U185 ( .A(n1649), .B(n1650), .Y(n1648) );
  AND2X2 U186 ( .A(n1654), .B(n1655), .Y(n1653) );
  AND2X2 U187 ( .A(n1662), .B(n1663), .Y(n1661) );
  AND2X2 U188 ( .A(n1667), .B(n1668), .Y(n1666) );
  AND2X2 U190 ( .A(n1674), .B(n1675), .Y(n1673) );
  AND2X2 U191 ( .A(n1679), .B(n1680), .Y(n1678) );
  AND2X2 U192 ( .A(n1689), .B(n1690), .Y(n1688) );
  AND2X2 U193 ( .A(n1694), .B(n1695), .Y(n1693) );
  AND2X2 U195 ( .A(n1701), .B(n1702), .Y(n1700) );
  AND2X2 U196 ( .A(n1706), .B(n1707), .Y(n1705) );
  AND2X2 U197 ( .A(n1714), .B(n1715), .Y(n1713) );
  AND2X2 U198 ( .A(n1719), .B(n1720), .Y(n1718) );
  AND2X2 U200 ( .A(n1726), .B(n1727), .Y(n1725) );
  AND2X2 U201 ( .A(n1731), .B(n1732), .Y(n1730) );
  AND2X2 U208 ( .A(n1741), .B(n1742), .Y(n1740) );
  AND2X2 U209 ( .A(n1753), .B(n1754), .Y(n1752) );
  AND2X2 U212 ( .A(n1763), .B(n1764), .Y(n1762) );
  AND2X2 U213 ( .A(n1768), .B(n1769), .Y(n1767) );
  AND2X2 U214 ( .A(n1780), .B(n1781), .Y(n1779) );
  OR2X2 U215 ( .A(n1785), .B(n1786), .Y(n1784) );
  AND2X2 U216 ( .A(n1791), .B(n1792), .Y(n1790) );
  AND2X2 U218 ( .A(n1800), .B(n1801), .Y(n1799) );
  AND2X2 U219 ( .A(n1806), .B(n1807), .Y(n1805) );
  OAI21X1 U817 ( .A(n598), .B(n3710), .C(n1776), .Y(n1816) );
  AOI22X1 U818 ( .A(\data_in<8> ), .B(n600), .C(\data_in<0> ), .D(n601), .Y(
        n599) );
  OAI21X1 U819 ( .A(n598), .B(n3709), .C(n1775), .Y(n1817) );
  AOI22X1 U820 ( .A(\data_in<9> ), .B(n600), .C(\data_in<1> ), .D(n601), .Y(
        n602) );
  OAI21X1 U821 ( .A(n598), .B(n3708), .C(n1773), .Y(n1818) );
  AOI22X1 U822 ( .A(\data_in<10> ), .B(n600), .C(\data_in<2> ), .D(n601), .Y(
        n603) );
  OAI21X1 U823 ( .A(n598), .B(n3707), .C(n1771), .Y(n1819) );
  AOI22X1 U824 ( .A(\data_in<11> ), .B(n600), .C(\data_in<3> ), .D(n601), .Y(
        n604) );
  OAI21X1 U825 ( .A(n598), .B(n3706), .C(n1759), .Y(n1820) );
  AOI22X1 U826 ( .A(\data_in<12> ), .B(n600), .C(\data_in<4> ), .D(n601), .Y(
        n605) );
  OAI21X1 U827 ( .A(n598), .B(n3705), .C(n1758), .Y(n1821) );
  AOI22X1 U828 ( .A(\data_in<13> ), .B(n600), .C(\data_in<5> ), .D(n601), .Y(
        n606) );
  OAI21X1 U829 ( .A(n598), .B(n3704), .C(n1737), .Y(n1822) );
  AOI22X1 U830 ( .A(\data_in<14> ), .B(n600), .C(\data_in<6> ), .D(n601), .Y(
        n607) );
  OAI21X1 U831 ( .A(n598), .B(n3703), .C(n1736), .Y(n1823) );
  AOI22X1 U832 ( .A(\data_in<15> ), .B(n600), .C(\data_in<7> ), .D(n601), .Y(
        n608) );
  OAI21X1 U833 ( .A(n2454), .B(n612), .C(n2460), .Y(n610) );
  OAI21X1 U834 ( .A(n3175), .B(n3702), .C(n1722), .Y(n1824) );
  AOI22X1 U835 ( .A(n615), .B(\data_in<8> ), .C(n616), .D(\data_in<0> ), .Y(
        n614) );
  OAI21X1 U836 ( .A(n3175), .B(n3701), .C(n1721), .Y(n1825) );
  AOI22X1 U837 ( .A(n615), .B(\data_in<9> ), .C(n616), .D(\data_in<1> ), .Y(
        n617) );
  OAI21X1 U838 ( .A(n3175), .B(n3700), .C(n1710), .Y(n1826) );
  AOI22X1 U839 ( .A(n615), .B(\data_in<10> ), .C(n616), .D(\data_in<2> ), .Y(
        n618) );
  OAI21X1 U840 ( .A(n3175), .B(n3699), .C(n1709), .Y(n1827) );
  AOI22X1 U841 ( .A(n615), .B(\data_in<11> ), .C(n616), .D(\data_in<3> ), .Y(
        n619) );
  OAI21X1 U842 ( .A(n3175), .B(n3698), .C(n1697), .Y(n1828) );
  AOI22X1 U843 ( .A(n615), .B(\data_in<12> ), .C(n616), .D(\data_in<4> ), .Y(
        n620) );
  OAI21X1 U844 ( .A(n3175), .B(n3697), .C(n1696), .Y(n1829) );
  AOI22X1 U845 ( .A(n615), .B(\data_in<13> ), .C(n616), .D(\data_in<5> ), .Y(
        n621) );
  OAI21X1 U846 ( .A(n3175), .B(n3696), .C(n1685), .Y(n1830) );
  AOI22X1 U847 ( .A(n615), .B(\data_in<14> ), .C(n616), .D(\data_in<6> ), .Y(
        n622) );
  OAI21X1 U848 ( .A(n3175), .B(n3695), .C(n1684), .Y(n1831) );
  AOI22X1 U849 ( .A(n615), .B(\data_in<15> ), .C(n616), .D(\data_in<7> ), .Y(
        n623) );
  AOI21X1 U850 ( .A(n2460), .B(n2563), .C(n2452), .Y(n613) );
  OAI21X1 U851 ( .A(n3174), .B(n3694), .C(n1670), .Y(n1832) );
  AOI22X1 U852 ( .A(n628), .B(\data_in<8> ), .C(n629), .D(\data_in<0> ), .Y(
        n627) );
  OAI21X1 U853 ( .A(n3174), .B(n3693), .C(n1669), .Y(n1833) );
  AOI22X1 U854 ( .A(n628), .B(\data_in<9> ), .C(n629), .D(\data_in<1> ), .Y(
        n630) );
  OAI21X1 U855 ( .A(n3174), .B(n3692), .C(n1658), .Y(n1834) );
  AOI22X1 U856 ( .A(n628), .B(\data_in<10> ), .C(n629), .D(\data_in<2> ), .Y(
        n631) );
  OAI21X1 U857 ( .A(n3174), .B(n3691), .C(n1657), .Y(n1835) );
  AOI22X1 U858 ( .A(n628), .B(\data_in<11> ), .C(n629), .D(\data_in<3> ), .Y(
        n632) );
  OAI21X1 U859 ( .A(n3174), .B(n3690), .C(n1645), .Y(n1836) );
  AOI22X1 U860 ( .A(n628), .B(\data_in<12> ), .C(n629), .D(\data_in<4> ), .Y(
        n633) );
  OAI21X1 U861 ( .A(n3174), .B(n3689), .C(n1644), .Y(n1837) );
  AOI22X1 U862 ( .A(n628), .B(\data_in<13> ), .C(n629), .D(\data_in<5> ), .Y(
        n634) );
  OAI21X1 U863 ( .A(n3174), .B(n3688), .C(n1633), .Y(n1838) );
  AOI22X1 U864 ( .A(n628), .B(\data_in<14> ), .C(n629), .D(\data_in<6> ), .Y(
        n635) );
  OAI21X1 U865 ( .A(n3174), .B(n3687), .C(n1632), .Y(n1839) );
  AOI22X1 U866 ( .A(n628), .B(\data_in<15> ), .C(n629), .D(\data_in<7> ), .Y(
        n636) );
  AOI21X1 U867 ( .A(n2563), .B(n2560), .C(n2452), .Y(n626) );
  OAI21X1 U868 ( .A(n3173), .B(n3686), .C(n1618), .Y(n1840) );
  AOI22X1 U869 ( .A(n640), .B(\data_in<8> ), .C(n641), .D(\data_in<0> ), .Y(
        n639) );
  OAI21X1 U870 ( .A(n3173), .B(n3685), .C(n1617), .Y(n1841) );
  AOI22X1 U871 ( .A(n640), .B(\data_in<9> ), .C(n641), .D(\data_in<1> ), .Y(
        n642) );
  OAI21X1 U872 ( .A(n3173), .B(n3684), .C(n1606), .Y(n1842) );
  AOI22X1 U873 ( .A(n640), .B(\data_in<10> ), .C(n641), .D(\data_in<2> ), .Y(
        n643) );
  OAI21X1 U874 ( .A(n3173), .B(n3683), .C(n1605), .Y(n1843) );
  AOI22X1 U875 ( .A(n640), .B(\data_in<11> ), .C(n641), .D(\data_in<3> ), .Y(
        n644) );
  OAI21X1 U876 ( .A(n3173), .B(n3682), .C(n1593), .Y(n1844) );
  AOI22X1 U877 ( .A(n640), .B(\data_in<12> ), .C(n641), .D(\data_in<4> ), .Y(
        n645) );
  OAI21X1 U878 ( .A(n3173), .B(n3681), .C(n1592), .Y(n1845) );
  AOI22X1 U879 ( .A(n640), .B(\data_in<13> ), .C(n641), .D(\data_in<5> ), .Y(
        n646) );
  OAI21X1 U880 ( .A(n3173), .B(n3680), .C(n1581), .Y(n1846) );
  AOI22X1 U881 ( .A(n640), .B(\data_in<14> ), .C(n641), .D(\data_in<6> ), .Y(
        n647) );
  OAI21X1 U882 ( .A(n3173), .B(n3679), .C(n1580), .Y(n1847) );
  AOI22X1 U883 ( .A(n640), .B(\data_in<15> ), .C(n641), .D(\data_in<7> ), .Y(
        n648) );
  AOI21X1 U884 ( .A(n2560), .B(n2561), .C(n2452), .Y(n638) );
  OAI21X1 U885 ( .A(n3172), .B(n3678), .C(n1566), .Y(n1848) );
  AOI22X1 U886 ( .A(n652), .B(\data_in<8> ), .C(n653), .D(\data_in<0> ), .Y(
        n651) );
  OAI21X1 U887 ( .A(n3172), .B(n3677), .C(n1565), .Y(n1849) );
  AOI22X1 U888 ( .A(n652), .B(\data_in<9> ), .C(n653), .D(\data_in<1> ), .Y(
        n654) );
  OAI21X1 U889 ( .A(n3172), .B(n3676), .C(n1554), .Y(n1850) );
  AOI22X1 U890 ( .A(n652), .B(\data_in<10> ), .C(n653), .D(\data_in<2> ), .Y(
        n655) );
  OAI21X1 U891 ( .A(n3172), .B(n3675), .C(n1553), .Y(n1851) );
  AOI22X1 U892 ( .A(n652), .B(\data_in<11> ), .C(n653), .D(\data_in<3> ), .Y(
        n656) );
  OAI21X1 U893 ( .A(n3172), .B(n3674), .C(n1541), .Y(n1852) );
  AOI22X1 U894 ( .A(n652), .B(\data_in<12> ), .C(n653), .D(\data_in<4> ), .Y(
        n657) );
  OAI21X1 U895 ( .A(n3172), .B(n3673), .C(n1540), .Y(n1853) );
  AOI22X1 U896 ( .A(n652), .B(\data_in<13> ), .C(n653), .D(\data_in<5> ), .Y(
        n658) );
  OAI21X1 U897 ( .A(n3172), .B(n3672), .C(n1529), .Y(n1854) );
  AOI22X1 U898 ( .A(n652), .B(\data_in<14> ), .C(n653), .D(\data_in<6> ), .Y(
        n659) );
  OAI21X1 U899 ( .A(n3172), .B(n3671), .C(n1528), .Y(n1855) );
  AOI22X1 U900 ( .A(n652), .B(\data_in<15> ), .C(n653), .D(\data_in<7> ), .Y(
        n660) );
  AOI21X1 U901 ( .A(n2561), .B(n2556), .C(n2452), .Y(n650) );
  OAI21X1 U902 ( .A(n3171), .B(n3670), .C(n1514), .Y(n1856) );
  AOI22X1 U903 ( .A(n664), .B(\data_in<8> ), .C(n665), .D(\data_in<0> ), .Y(
        n663) );
  OAI21X1 U904 ( .A(n3171), .B(n3669), .C(n1513), .Y(n1857) );
  AOI22X1 U905 ( .A(n664), .B(\data_in<9> ), .C(n665), .D(\data_in<1> ), .Y(
        n666) );
  OAI21X1 U906 ( .A(n3171), .B(n3668), .C(n1502), .Y(n1858) );
  AOI22X1 U907 ( .A(n664), .B(\data_in<10> ), .C(n665), .D(\data_in<2> ), .Y(
        n667) );
  OAI21X1 U908 ( .A(n3171), .B(n3667), .C(n1501), .Y(n1859) );
  AOI22X1 U909 ( .A(n664), .B(\data_in<11> ), .C(n665), .D(\data_in<3> ), .Y(
        n668) );
  OAI21X1 U910 ( .A(n3171), .B(n3666), .C(n1489), .Y(n1860) );
  AOI22X1 U911 ( .A(n664), .B(\data_in<12> ), .C(n665), .D(\data_in<4> ), .Y(
        n669) );
  OAI21X1 U912 ( .A(n3171), .B(n3665), .C(n1488), .Y(n1861) );
  AOI22X1 U913 ( .A(n664), .B(\data_in<13> ), .C(n665), .D(\data_in<5> ), .Y(
        n670) );
  OAI21X1 U914 ( .A(n3171), .B(n3664), .C(n1477), .Y(n1862) );
  AOI22X1 U915 ( .A(n664), .B(\data_in<14> ), .C(n665), .D(\data_in<6> ), .Y(
        n671) );
  OAI21X1 U916 ( .A(n3171), .B(n3663), .C(n1476), .Y(n1863) );
  AOI22X1 U917 ( .A(n664), .B(\data_in<15> ), .C(n665), .D(\data_in<7> ), .Y(
        n672) );
  AOI21X1 U918 ( .A(n2556), .B(n2557), .C(n2452), .Y(n662) );
  OAI21X1 U919 ( .A(n3170), .B(n3662), .C(n1462), .Y(n1864) );
  AOI22X1 U920 ( .A(n676), .B(\data_in<8> ), .C(n677), .D(\data_in<0> ), .Y(
        n675) );
  OAI21X1 U921 ( .A(n3170), .B(n3661), .C(n1461), .Y(n1865) );
  AOI22X1 U922 ( .A(n676), .B(\data_in<9> ), .C(n677), .D(\data_in<1> ), .Y(
        n678) );
  OAI21X1 U923 ( .A(n3170), .B(n3660), .C(n1450), .Y(n1866) );
  AOI22X1 U924 ( .A(n676), .B(\data_in<10> ), .C(n677), .D(\data_in<2> ), .Y(
        n679) );
  OAI21X1 U925 ( .A(n3170), .B(n3659), .C(n1449), .Y(n1867) );
  AOI22X1 U926 ( .A(n676), .B(\data_in<11> ), .C(n677), .D(\data_in<3> ), .Y(
        n680) );
  OAI21X1 U927 ( .A(n3170), .B(n3658), .C(n1437), .Y(n1868) );
  AOI22X1 U928 ( .A(n676), .B(\data_in<12> ), .C(n677), .D(\data_in<4> ), .Y(
        n681) );
  OAI21X1 U929 ( .A(n3170), .B(n3657), .C(n1436), .Y(n1869) );
  AOI22X1 U930 ( .A(n676), .B(\data_in<13> ), .C(n677), .D(\data_in<5> ), .Y(
        n682) );
  OAI21X1 U931 ( .A(n3170), .B(n3656), .C(n1425), .Y(n1870) );
  AOI22X1 U932 ( .A(n676), .B(\data_in<14> ), .C(n677), .D(\data_in<6> ), .Y(
        n683) );
  OAI21X1 U933 ( .A(n3170), .B(n3655), .C(n1424), .Y(n1871) );
  AOI22X1 U934 ( .A(n676), .B(\data_in<15> ), .C(n677), .D(\data_in<7> ), .Y(
        n684) );
  AOI21X1 U935 ( .A(n2557), .B(n2552), .C(n2452), .Y(n674) );
  OAI21X1 U936 ( .A(n3169), .B(n3654), .C(n1410), .Y(n1872) );
  AOI22X1 U937 ( .A(n688), .B(\data_in<8> ), .C(n689), .D(\data_in<0> ), .Y(
        n687) );
  OAI21X1 U938 ( .A(n3169), .B(n3653), .C(n1409), .Y(n1873) );
  AOI22X1 U939 ( .A(n688), .B(\data_in<9> ), .C(n689), .D(\data_in<1> ), .Y(
        n690) );
  OAI21X1 U940 ( .A(n3169), .B(n3652), .C(n1397), .Y(n1874) );
  AOI22X1 U941 ( .A(n688), .B(\data_in<10> ), .C(n689), .D(\data_in<2> ), .Y(
        n691) );
  OAI21X1 U942 ( .A(n3169), .B(n3651), .C(n1396), .Y(n1875) );
  AOI22X1 U943 ( .A(n688), .B(\data_in<11> ), .C(n689), .D(\data_in<3> ), .Y(
        n692) );
  OAI21X1 U944 ( .A(n3169), .B(n3650), .C(n1384), .Y(n1876) );
  AOI22X1 U945 ( .A(n688), .B(\data_in<12> ), .C(n689), .D(\data_in<4> ), .Y(
        n693) );
  OAI21X1 U946 ( .A(n3169), .B(n3649), .C(n1383), .Y(n1877) );
  AOI22X1 U947 ( .A(n688), .B(\data_in<13> ), .C(n689), .D(\data_in<5> ), .Y(
        n694) );
  OAI21X1 U948 ( .A(n3169), .B(n3648), .C(n1372), .Y(n1878) );
  AOI22X1 U949 ( .A(n688), .B(\data_in<14> ), .C(n689), .D(\data_in<6> ), .Y(
        n695) );
  OAI21X1 U950 ( .A(n3169), .B(n3647), .C(n1371), .Y(n1879) );
  AOI22X1 U951 ( .A(n688), .B(\data_in<15> ), .C(n689), .D(\data_in<7> ), .Y(
        n696) );
  AOI21X1 U952 ( .A(n2552), .B(n2553), .C(n3179), .Y(n686) );
  OAI21X1 U953 ( .A(n3168), .B(n3646), .C(n1369), .Y(n1880) );
  AOI22X1 U954 ( .A(n700), .B(\data_in<8> ), .C(n701), .D(\data_in<0> ), .Y(
        n699) );
  OAI21X1 U955 ( .A(n3168), .B(n3645), .C(n1366), .Y(n1881) );
  AOI22X1 U956 ( .A(n700), .B(\data_in<9> ), .C(n701), .D(\data_in<1> ), .Y(
        n702) );
  OAI21X1 U957 ( .A(n3168), .B(n3644), .C(n1365), .Y(n1882) );
  AOI22X1 U958 ( .A(n700), .B(\data_in<10> ), .C(n701), .D(\data_in<2> ), .Y(
        n703) );
  OAI21X1 U959 ( .A(n3168), .B(n3643), .C(n1364), .Y(n1883) );
  AOI22X1 U960 ( .A(n700), .B(\data_in<11> ), .C(n701), .D(\data_in<3> ), .Y(
        n704) );
  OAI21X1 U961 ( .A(n3168), .B(n3642), .C(n1363), .Y(n1884) );
  AOI22X1 U962 ( .A(n700), .B(\data_in<12> ), .C(n701), .D(\data_in<4> ), .Y(
        n705) );
  OAI21X1 U963 ( .A(n3168), .B(n3641), .C(n1362), .Y(n1885) );
  AOI22X1 U964 ( .A(n700), .B(\data_in<13> ), .C(n701), .D(\data_in<5> ), .Y(
        n706) );
  OAI21X1 U965 ( .A(n3168), .B(n3640), .C(n1361), .Y(n1886) );
  AOI22X1 U966 ( .A(n700), .B(\data_in<14> ), .C(n701), .D(\data_in<6> ), .Y(
        n707) );
  OAI21X1 U967 ( .A(n3168), .B(n3639), .C(n1360), .Y(n1887) );
  AOI22X1 U968 ( .A(n700), .B(\data_in<15> ), .C(n701), .D(\data_in<7> ), .Y(
        n708) );
  AOI21X1 U969 ( .A(n2553), .B(n2578), .C(n3179), .Y(n698) );
  OAI21X1 U970 ( .A(n3167), .B(n3638), .C(n1359), .Y(n1888) );
  AOI22X1 U971 ( .A(n712), .B(\data_in<8> ), .C(n713), .D(\data_in<0> ), .Y(
        n711) );
  OAI21X1 U972 ( .A(n3167), .B(n3637), .C(n1358), .Y(n1889) );
  AOI22X1 U973 ( .A(n712), .B(\data_in<9> ), .C(n713), .D(\data_in<1> ), .Y(
        n714) );
  OAI21X1 U974 ( .A(n3167), .B(n3636), .C(n1357), .Y(n1890) );
  AOI22X1 U975 ( .A(n712), .B(\data_in<10> ), .C(n713), .D(\data_in<2> ), .Y(
        n715) );
  OAI21X1 U976 ( .A(n3167), .B(n3635), .C(n1345), .Y(n1891) );
  AOI22X1 U977 ( .A(n712), .B(\data_in<11> ), .C(n713), .D(\data_in<3> ), .Y(
        n716) );
  OAI21X1 U978 ( .A(n3167), .B(n3634), .C(n1333), .Y(n1892) );
  AOI22X1 U979 ( .A(n712), .B(\data_in<12> ), .C(n713), .D(\data_in<4> ), .Y(
        n717) );
  OAI21X1 U980 ( .A(n3167), .B(n3633), .C(n1321), .Y(n1893) );
  AOI22X1 U981 ( .A(n712), .B(\data_in<13> ), .C(n713), .D(\data_in<5> ), .Y(
        n718) );
  OAI21X1 U982 ( .A(n3167), .B(n3632), .C(n1309), .Y(n1894) );
  AOI22X1 U983 ( .A(n712), .B(\data_in<14> ), .C(n713), .D(\data_in<6> ), .Y(
        n719) );
  OAI21X1 U984 ( .A(n3167), .B(n3631), .C(n1297), .Y(n1895) );
  AOI22X1 U985 ( .A(n712), .B(\data_in<15> ), .C(n713), .D(\data_in<7> ), .Y(
        n720) );
  AOI21X1 U986 ( .A(n2578), .B(n2579), .C(n3179), .Y(n710) );
  OAI21X1 U987 ( .A(n3166), .B(n3630), .C(n1285), .Y(n1896) );
  AOI22X1 U988 ( .A(n724), .B(\data_in<8> ), .C(n725), .D(\data_in<0> ), .Y(
        n723) );
  OAI21X1 U989 ( .A(n3166), .B(n3629), .C(n1273), .Y(n1897) );
  AOI22X1 U990 ( .A(n724), .B(\data_in<9> ), .C(n725), .D(\data_in<1> ), .Y(
        n726) );
  OAI21X1 U991 ( .A(n3166), .B(n3628), .C(n1261), .Y(n1898) );
  AOI22X1 U992 ( .A(n724), .B(\data_in<10> ), .C(n725), .D(\data_in<2> ), .Y(
        n727) );
  OAI21X1 U993 ( .A(n3166), .B(n3627), .C(n1249), .Y(n1899) );
  AOI22X1 U994 ( .A(n724), .B(\data_in<11> ), .C(n725), .D(\data_in<3> ), .Y(
        n728) );
  OAI21X1 U995 ( .A(n3166), .B(n3626), .C(n1237), .Y(n1900) );
  AOI22X1 U996 ( .A(n724), .B(\data_in<12> ), .C(n725), .D(\data_in<4> ), .Y(
        n729) );
  OAI21X1 U997 ( .A(n3166), .B(n3625), .C(n1225), .Y(n1901) );
  AOI22X1 U998 ( .A(n724), .B(\data_in<13> ), .C(n725), .D(\data_in<5> ), .Y(
        n730) );
  OAI21X1 U999 ( .A(n3166), .B(n3624), .C(n1213), .Y(n1902) );
  AOI22X1 U1000 ( .A(n724), .B(\data_in<14> ), .C(n725), .D(\data_in<6> ), .Y(
        n731) );
  OAI21X1 U1001 ( .A(n3166), .B(n3623), .C(n1201), .Y(n1903) );
  AOI22X1 U1002 ( .A(n724), .B(\data_in<15> ), .C(n725), .D(\data_in<7> ), .Y(
        n732) );
  AOI21X1 U1003 ( .A(n2579), .B(n2574), .C(n3179), .Y(n722) );
  OAI21X1 U1004 ( .A(n3165), .B(n3622), .C(n1189), .Y(n1904) );
  AOI22X1 U1005 ( .A(n736), .B(\data_in<8> ), .C(n737), .D(\data_in<0> ), .Y(
        n735) );
  OAI21X1 U1006 ( .A(n3165), .B(n3621), .C(n1177), .Y(n1905) );
  AOI22X1 U1007 ( .A(n736), .B(\data_in<9> ), .C(n737), .D(\data_in<1> ), .Y(
        n738) );
  OAI21X1 U1008 ( .A(n3165), .B(n3620), .C(n1165), .Y(n1906) );
  AOI22X1 U1009 ( .A(n736), .B(\data_in<10> ), .C(n737), .D(\data_in<2> ), .Y(
        n739) );
  OAI21X1 U1010 ( .A(n3165), .B(n3619), .C(n1153), .Y(n1907) );
  AOI22X1 U1011 ( .A(n736), .B(\data_in<11> ), .C(n737), .D(\data_in<3> ), .Y(
        n740) );
  OAI21X1 U1012 ( .A(n3165), .B(n3618), .C(n1141), .Y(n1908) );
  AOI22X1 U1013 ( .A(n736), .B(\data_in<12> ), .C(n737), .D(\data_in<4> ), .Y(
        n741) );
  OAI21X1 U1014 ( .A(n3165), .B(n3617), .C(n1129), .Y(n1909) );
  AOI22X1 U1015 ( .A(n736), .B(\data_in<13> ), .C(n737), .D(\data_in<5> ), .Y(
        n742) );
  OAI21X1 U1016 ( .A(n3165), .B(n3616), .C(n1117), .Y(n1910) );
  AOI22X1 U1017 ( .A(n736), .B(\data_in<14> ), .C(n737), .D(\data_in<6> ), .Y(
        n743) );
  OAI21X1 U1018 ( .A(n3165), .B(n3615), .C(n1105), .Y(n1911) );
  AOI22X1 U1019 ( .A(n736), .B(\data_in<15> ), .C(n737), .D(\data_in<7> ), .Y(
        n744) );
  AOI21X1 U1020 ( .A(n2574), .B(n2575), .C(n3179), .Y(n734) );
  OAI21X1 U1021 ( .A(n3164), .B(n3614), .C(n1093), .Y(n1912) );
  AOI22X1 U1022 ( .A(n748), .B(\data_in<8> ), .C(n749), .D(\data_in<0> ), .Y(
        n747) );
  OAI21X1 U1023 ( .A(n3164), .B(n3613), .C(n1081), .Y(n1913) );
  AOI22X1 U1024 ( .A(n748), .B(\data_in<9> ), .C(n749), .D(\data_in<1> ), .Y(
        n750) );
  OAI21X1 U1025 ( .A(n3164), .B(n3612), .C(n1069), .Y(n1914) );
  AOI22X1 U1026 ( .A(n748), .B(\data_in<10> ), .C(n749), .D(\data_in<2> ), .Y(
        n751) );
  OAI21X1 U1027 ( .A(n3164), .B(n3611), .C(n1057), .Y(n1915) );
  AOI22X1 U1028 ( .A(n748), .B(\data_in<11> ), .C(n749), .D(\data_in<3> ), .Y(
        n752) );
  OAI21X1 U1029 ( .A(n3164), .B(n3610), .C(n1045), .Y(n1916) );
  AOI22X1 U1030 ( .A(n748), .B(\data_in<12> ), .C(n749), .D(\data_in<4> ), .Y(
        n753) );
  OAI21X1 U1031 ( .A(n3164), .B(n3609), .C(n1033), .Y(n1917) );
  AOI22X1 U1032 ( .A(n748), .B(\data_in<13> ), .C(n749), .D(\data_in<5> ), .Y(
        n754) );
  OAI21X1 U1033 ( .A(n3164), .B(n3608), .C(n1021), .Y(n1918) );
  AOI22X1 U1034 ( .A(n748), .B(\data_in<14> ), .C(n749), .D(\data_in<6> ), .Y(
        n755) );
  OAI21X1 U1035 ( .A(n3164), .B(n3607), .C(n1009), .Y(n1919) );
  AOI22X1 U1036 ( .A(n748), .B(\data_in<15> ), .C(n749), .D(\data_in<7> ), .Y(
        n756) );
  AOI21X1 U1037 ( .A(n2575), .B(n2570), .C(n3179), .Y(n746) );
  OAI21X1 U1038 ( .A(n3163), .B(n3606), .C(n997), .Y(n1920) );
  AOI22X1 U1039 ( .A(n760), .B(\data_in<8> ), .C(n761), .D(\data_in<0> ), .Y(
        n759) );
  OAI21X1 U1040 ( .A(n3163), .B(n3605), .C(n985), .Y(n1921) );
  AOI22X1 U1041 ( .A(n760), .B(\data_in<9> ), .C(n761), .D(\data_in<1> ), .Y(
        n762) );
  OAI21X1 U1042 ( .A(n3163), .B(n3604), .C(n973), .Y(n1922) );
  AOI22X1 U1043 ( .A(n760), .B(\data_in<10> ), .C(n761), .D(\data_in<2> ), .Y(
        n763) );
  OAI21X1 U1044 ( .A(n3163), .B(n3603), .C(n961), .Y(n1923) );
  AOI22X1 U1045 ( .A(n760), .B(\data_in<11> ), .C(n761), .D(\data_in<3> ), .Y(
        n764) );
  OAI21X1 U1046 ( .A(n3163), .B(n3602), .C(n949), .Y(n1924) );
  AOI22X1 U1047 ( .A(n760), .B(\data_in<12> ), .C(n761), .D(\data_in<4> ), .Y(
        n765) );
  OAI21X1 U1048 ( .A(n3163), .B(n3601), .C(n937), .Y(n1925) );
  AOI22X1 U1049 ( .A(n760), .B(\data_in<13> ), .C(n761), .D(\data_in<5> ), .Y(
        n766) );
  OAI21X1 U1050 ( .A(n3163), .B(n3600), .C(n925), .Y(n1926) );
  AOI22X1 U1051 ( .A(n760), .B(\data_in<14> ), .C(n761), .D(\data_in<6> ), .Y(
        n767) );
  OAI21X1 U1052 ( .A(n3163), .B(n3599), .C(n913), .Y(n1927) );
  AOI22X1 U1053 ( .A(n760), .B(\data_in<15> ), .C(n761), .D(\data_in<7> ), .Y(
        n768) );
  AOI21X1 U1054 ( .A(n2570), .B(n2571), .C(n3179), .Y(n758) );
  OAI21X1 U1055 ( .A(n3162), .B(n3598), .C(n901), .Y(n1928) );
  AOI22X1 U1056 ( .A(n772), .B(\data_in<8> ), .C(n773), .D(\data_in<0> ), .Y(
        n771) );
  OAI21X1 U1057 ( .A(n3162), .B(n3597), .C(n889), .Y(n1929) );
  AOI22X1 U1058 ( .A(n772), .B(\data_in<9> ), .C(n773), .D(\data_in<1> ), .Y(
        n774) );
  OAI21X1 U1059 ( .A(n3162), .B(n3596), .C(n877), .Y(n1930) );
  AOI22X1 U1060 ( .A(n772), .B(\data_in<10> ), .C(n773), .D(\data_in<2> ), .Y(
        n775) );
  OAI21X1 U1061 ( .A(n3162), .B(n3595), .C(n865), .Y(n1931) );
  AOI22X1 U1062 ( .A(n772), .B(\data_in<11> ), .C(n773), .D(\data_in<3> ), .Y(
        n776) );
  OAI21X1 U1063 ( .A(n3162), .B(n3594), .C(n853), .Y(n1932) );
  AOI22X1 U1064 ( .A(n772), .B(\data_in<12> ), .C(n773), .D(\data_in<4> ), .Y(
        n777) );
  OAI21X1 U1065 ( .A(n3162), .B(n3593), .C(n841), .Y(n1933) );
  AOI22X1 U1066 ( .A(n772), .B(\data_in<13> ), .C(n773), .D(\data_in<5> ), .Y(
        n778) );
  OAI21X1 U1067 ( .A(n3162), .B(n3592), .C(n829), .Y(n1934) );
  AOI22X1 U1068 ( .A(n772), .B(\data_in<14> ), .C(n773), .D(\data_in<6> ), .Y(
        n779) );
  OAI21X1 U1069 ( .A(n3162), .B(n3591), .C(n817), .Y(n1935) );
  AOI22X1 U1070 ( .A(n772), .B(\data_in<15> ), .C(n773), .D(\data_in<7> ), .Y(
        n780) );
  AOI21X1 U1071 ( .A(n2571), .B(n2566), .C(n3179), .Y(n770) );
  OAI21X1 U1072 ( .A(n3161), .B(n3590), .C(n805), .Y(n1936) );
  AOI22X1 U1073 ( .A(n784), .B(\data_in<8> ), .C(n785), .D(\data_in<0> ), .Y(
        n783) );
  OAI21X1 U1074 ( .A(n3161), .B(n3589), .C(n793), .Y(n1937) );
  AOI22X1 U1075 ( .A(n784), .B(\data_in<9> ), .C(n785), .D(\data_in<1> ), .Y(
        n786) );
  OAI21X1 U1076 ( .A(n3161), .B(n3588), .C(n781), .Y(n1938) );
  AOI22X1 U1077 ( .A(n784), .B(\data_in<10> ), .C(n785), .D(\data_in<2> ), .Y(
        n787) );
  OAI21X1 U1078 ( .A(n3161), .B(n3587), .C(n769), .Y(n1939) );
  AOI22X1 U1079 ( .A(n784), .B(\data_in<11> ), .C(n785), .D(\data_in<3> ), .Y(
        n788) );
  OAI21X1 U1080 ( .A(n3161), .B(n3586), .C(n757), .Y(n1940) );
  AOI22X1 U1081 ( .A(n784), .B(\data_in<12> ), .C(n785), .D(\data_in<4> ), .Y(
        n789) );
  OAI21X1 U1082 ( .A(n3161), .B(n3585), .C(n745), .Y(n1941) );
  AOI22X1 U1083 ( .A(n784), .B(\data_in<13> ), .C(n785), .D(\data_in<5> ), .Y(
        n790) );
  OAI21X1 U1084 ( .A(n3161), .B(n3584), .C(n733), .Y(n1942) );
  AOI22X1 U1085 ( .A(n784), .B(\data_in<14> ), .C(n785), .D(\data_in<6> ), .Y(
        n791) );
  OAI21X1 U1086 ( .A(n3161), .B(n3583), .C(n721), .Y(n1943) );
  AOI22X1 U1087 ( .A(n784), .B(\data_in<15> ), .C(n785), .D(\data_in<7> ), .Y(
        n792) );
  AOI21X1 U1088 ( .A(n2566), .B(n2567), .C(n3179), .Y(n782) );
  OAI21X1 U1089 ( .A(n3160), .B(n3582), .C(n709), .Y(n1944) );
  AOI22X1 U1090 ( .A(n796), .B(\data_in<8> ), .C(n797), .D(\data_in<0> ), .Y(
        n795) );
  OAI21X1 U1091 ( .A(n3160), .B(n3581), .C(n697), .Y(n1945) );
  AOI22X1 U1092 ( .A(n796), .B(\data_in<9> ), .C(n797), .D(\data_in<1> ), .Y(
        n798) );
  OAI21X1 U1093 ( .A(n3160), .B(n3580), .C(n685), .Y(n1946) );
  AOI22X1 U1094 ( .A(n796), .B(\data_in<10> ), .C(n797), .D(\data_in<2> ), .Y(
        n799) );
  OAI21X1 U1095 ( .A(n3160), .B(n3579), .C(n673), .Y(n1947) );
  AOI22X1 U1096 ( .A(n796), .B(\data_in<11> ), .C(n797), .D(\data_in<3> ), .Y(
        n800) );
  OAI21X1 U1097 ( .A(n3160), .B(n3578), .C(n661), .Y(n1948) );
  AOI22X1 U1098 ( .A(n796), .B(\data_in<12> ), .C(n797), .D(\data_in<4> ), .Y(
        n801) );
  OAI21X1 U1099 ( .A(n3160), .B(n3577), .C(n649), .Y(n1949) );
  AOI22X1 U1100 ( .A(n796), .B(\data_in<13> ), .C(n797), .D(\data_in<5> ), .Y(
        n802) );
  OAI21X1 U1101 ( .A(n3160), .B(n3576), .C(n637), .Y(n1950) );
  AOI22X1 U1102 ( .A(n796), .B(\data_in<14> ), .C(n797), .D(\data_in<6> ), .Y(
        n803) );
  OAI21X1 U1103 ( .A(n3160), .B(n3575), .C(n624), .Y(n1951) );
  AOI22X1 U1104 ( .A(n796), .B(\data_in<15> ), .C(n797), .D(\data_in<7> ), .Y(
        n804) );
  AOI21X1 U1105 ( .A(n2567), .B(n2532), .C(n3179), .Y(n794) );
  OAI21X1 U1106 ( .A(n3159), .B(n3574), .C(n611), .Y(n1952) );
  AOI22X1 U1107 ( .A(n808), .B(\data_in<8> ), .C(n809), .D(\data_in<0> ), .Y(
        n807) );
  OAI21X1 U1108 ( .A(n3159), .B(n3573), .C(n609), .Y(n1953) );
  AOI22X1 U1109 ( .A(n808), .B(\data_in<9> ), .C(n809), .D(\data_in<1> ), .Y(
        n810) );
  OAI21X1 U1110 ( .A(n3159), .B(n3572), .C(n597), .Y(n1954) );
  AOI22X1 U1111 ( .A(n808), .B(\data_in<10> ), .C(n809), .D(\data_in<2> ), .Y(
        n811) );
  OAI21X1 U1112 ( .A(n3159), .B(n3571), .C(n596), .Y(n1955) );
  AOI22X1 U1113 ( .A(n808), .B(\data_in<11> ), .C(n809), .D(\data_in<3> ), .Y(
        n812) );
  OAI21X1 U1114 ( .A(n3159), .B(n3570), .C(n595), .Y(n1956) );
  AOI22X1 U1115 ( .A(n808), .B(\data_in<12> ), .C(n809), .D(\data_in<4> ), .Y(
        n813) );
  OAI21X1 U1116 ( .A(n3159), .B(n3569), .C(n594), .Y(n1957) );
  AOI22X1 U1117 ( .A(n808), .B(\data_in<13> ), .C(n809), .D(\data_in<5> ), .Y(
        n814) );
  OAI21X1 U1118 ( .A(n3159), .B(n3568), .C(n593), .Y(n1958) );
  AOI22X1 U1119 ( .A(n808), .B(\data_in<14> ), .C(n809), .D(\data_in<6> ), .Y(
        n815) );
  OAI21X1 U1120 ( .A(n3159), .B(n3567), .C(n592), .Y(n1959) );
  AOI22X1 U1121 ( .A(n808), .B(\data_in<15> ), .C(n809), .D(\data_in<7> ), .Y(
        n816) );
  AOI21X1 U1122 ( .A(n2532), .B(n2533), .C(n3179), .Y(n806) );
  OAI21X1 U1123 ( .A(n3158), .B(n3566), .C(n591), .Y(n1960) );
  AOI22X1 U1124 ( .A(n820), .B(\data_in<8> ), .C(n821), .D(\data_in<0> ), .Y(
        n819) );
  OAI21X1 U1125 ( .A(n3158), .B(n3565), .C(n590), .Y(n1961) );
  AOI22X1 U1126 ( .A(n820), .B(\data_in<9> ), .C(n821), .D(\data_in<1> ), .Y(
        n822) );
  OAI21X1 U1127 ( .A(n3158), .B(n3564), .C(n589), .Y(n1962) );
  AOI22X1 U1128 ( .A(n820), .B(\data_in<10> ), .C(n821), .D(\data_in<2> ), .Y(
        n823) );
  OAI21X1 U1129 ( .A(n3158), .B(n3563), .C(n588), .Y(n1963) );
  AOI22X1 U1130 ( .A(n820), .B(\data_in<11> ), .C(n821), .D(\data_in<3> ), .Y(
        n824) );
  OAI21X1 U1131 ( .A(n3158), .B(n3562), .C(n587), .Y(n1964) );
  AOI22X1 U1132 ( .A(n820), .B(\data_in<12> ), .C(n821), .D(\data_in<4> ), .Y(
        n825) );
  OAI21X1 U1133 ( .A(n3158), .B(n3561), .C(n586), .Y(n1965) );
  AOI22X1 U1134 ( .A(n820), .B(\data_in<13> ), .C(n821), .D(\data_in<5> ), .Y(
        n826) );
  OAI21X1 U1135 ( .A(n3158), .B(n3560), .C(n585), .Y(n1966) );
  AOI22X1 U1136 ( .A(n820), .B(\data_in<14> ), .C(n821), .D(\data_in<6> ), .Y(
        n827) );
  OAI21X1 U1137 ( .A(n3158), .B(n3559), .C(n584), .Y(n1967) );
  AOI22X1 U1138 ( .A(n820), .B(\data_in<15> ), .C(n821), .D(\data_in<7> ), .Y(
        n828) );
  AOI21X1 U1139 ( .A(n2533), .B(n2528), .C(n3179), .Y(n818) );
  OAI21X1 U1140 ( .A(n3157), .B(n3558), .C(n583), .Y(n1968) );
  AOI22X1 U1141 ( .A(n832), .B(\data_in<8> ), .C(n833), .D(\data_in<0> ), .Y(
        n831) );
  OAI21X1 U1142 ( .A(n3157), .B(n3557), .C(n582), .Y(n1969) );
  AOI22X1 U1143 ( .A(n832), .B(\data_in<9> ), .C(n833), .D(\data_in<1> ), .Y(
        n834) );
  OAI21X1 U1144 ( .A(n3157), .B(n3556), .C(n581), .Y(n1970) );
  AOI22X1 U1145 ( .A(n832), .B(\data_in<10> ), .C(n833), .D(\data_in<2> ), .Y(
        n835) );
  OAI21X1 U1146 ( .A(n3157), .B(n3555), .C(n580), .Y(n1971) );
  AOI22X1 U1147 ( .A(n832), .B(\data_in<11> ), .C(n833), .D(\data_in<3> ), .Y(
        n836) );
  OAI21X1 U1148 ( .A(n3157), .B(n3554), .C(n579), .Y(n1972) );
  AOI22X1 U1149 ( .A(n832), .B(\data_in<12> ), .C(n833), .D(\data_in<4> ), .Y(
        n837) );
  OAI21X1 U1150 ( .A(n3157), .B(n3553), .C(n578), .Y(n1973) );
  AOI22X1 U1151 ( .A(n832), .B(\data_in<13> ), .C(n833), .D(\data_in<5> ), .Y(
        n838) );
  OAI21X1 U1152 ( .A(n3157), .B(n3552), .C(n577), .Y(n1974) );
  AOI22X1 U1153 ( .A(n832), .B(\data_in<14> ), .C(n833), .D(\data_in<6> ), .Y(
        n839) );
  OAI21X1 U1154 ( .A(n3157), .B(n3551), .C(n576), .Y(n1975) );
  AOI22X1 U1155 ( .A(n832), .B(\data_in<15> ), .C(n833), .D(\data_in<7> ), .Y(
        n840) );
  AOI21X1 U1156 ( .A(n2528), .B(n2529), .C(n3179), .Y(n830) );
  OAI21X1 U1157 ( .A(n3156), .B(n3550), .C(n575), .Y(n1976) );
  AOI22X1 U1158 ( .A(n844), .B(\data_in<8> ), .C(n845), .D(\data_in<0> ), .Y(
        n843) );
  OAI21X1 U1159 ( .A(n3156), .B(n3549), .C(n574), .Y(n1977) );
  AOI22X1 U1160 ( .A(n844), .B(\data_in<9> ), .C(n845), .D(\data_in<1> ), .Y(
        n846) );
  OAI21X1 U1161 ( .A(n3156), .B(n3548), .C(n573), .Y(n1978) );
  AOI22X1 U1162 ( .A(n844), .B(\data_in<10> ), .C(n845), .D(\data_in<2> ), .Y(
        n847) );
  OAI21X1 U1163 ( .A(n3156), .B(n3547), .C(n572), .Y(n1979) );
  AOI22X1 U1164 ( .A(n844), .B(\data_in<11> ), .C(n845), .D(\data_in<3> ), .Y(
        n848) );
  OAI21X1 U1165 ( .A(n3156), .B(n3546), .C(n571), .Y(n1980) );
  AOI22X1 U1166 ( .A(n844), .B(\data_in<12> ), .C(n845), .D(\data_in<4> ), .Y(
        n849) );
  OAI21X1 U1167 ( .A(n3156), .B(n3545), .C(n570), .Y(n1981) );
  AOI22X1 U1168 ( .A(n844), .B(\data_in<13> ), .C(n845), .D(\data_in<5> ), .Y(
        n850) );
  OAI21X1 U1169 ( .A(n3156), .B(n3544), .C(n569), .Y(n1982) );
  AOI22X1 U1170 ( .A(n844), .B(\data_in<14> ), .C(n845), .D(\data_in<6> ), .Y(
        n851) );
  OAI21X1 U1171 ( .A(n3156), .B(n3543), .C(n568), .Y(n1983) );
  AOI22X1 U1172 ( .A(n844), .B(\data_in<15> ), .C(n845), .D(\data_in<7> ), .Y(
        n852) );
  AOI21X1 U1173 ( .A(n2529), .B(n2524), .C(n3179), .Y(n842) );
  OAI21X1 U1174 ( .A(n3155), .B(n3542), .C(n567), .Y(n1984) );
  AOI22X1 U1175 ( .A(n856), .B(\data_in<8> ), .C(n857), .D(\data_in<0> ), .Y(
        n855) );
  OAI21X1 U1176 ( .A(n3155), .B(n3541), .C(n566), .Y(n1985) );
  AOI22X1 U1177 ( .A(n856), .B(\data_in<9> ), .C(n857), .D(\data_in<1> ), .Y(
        n858) );
  OAI21X1 U1178 ( .A(n3155), .B(n3540), .C(n565), .Y(n1986) );
  AOI22X1 U1179 ( .A(n856), .B(\data_in<10> ), .C(n857), .D(\data_in<2> ), .Y(
        n859) );
  OAI21X1 U1180 ( .A(n3155), .B(n3539), .C(n564), .Y(n1987) );
  AOI22X1 U1181 ( .A(n856), .B(\data_in<11> ), .C(n857), .D(\data_in<3> ), .Y(
        n860) );
  OAI21X1 U1182 ( .A(n3155), .B(n3538), .C(n563), .Y(n1988) );
  AOI22X1 U1183 ( .A(n856), .B(\data_in<12> ), .C(n857), .D(\data_in<4> ), .Y(
        n861) );
  OAI21X1 U1184 ( .A(n3155), .B(n3537), .C(n562), .Y(n1989) );
  AOI22X1 U1185 ( .A(n856), .B(\data_in<13> ), .C(n857), .D(\data_in<5> ), .Y(
        n862) );
  OAI21X1 U1186 ( .A(n3155), .B(n3536), .C(n561), .Y(n1990) );
  AOI22X1 U1187 ( .A(n856), .B(\data_in<14> ), .C(n857), .D(\data_in<6> ), .Y(
        n863) );
  OAI21X1 U1188 ( .A(n3155), .B(n3535), .C(n560), .Y(n1991) );
  AOI22X1 U1189 ( .A(n856), .B(\data_in<15> ), .C(n857), .D(\data_in<7> ), .Y(
        n864) );
  AOI21X1 U1190 ( .A(n2524), .B(n2525), .C(n3178), .Y(n854) );
  OAI21X1 U1191 ( .A(n3154), .B(n3534), .C(n559), .Y(n1992) );
  AOI22X1 U1192 ( .A(n868), .B(\data_in<8> ), .C(n869), .D(\data_in<0> ), .Y(
        n867) );
  OAI21X1 U1193 ( .A(n3154), .B(n3533), .C(n558), .Y(n1993) );
  AOI22X1 U1194 ( .A(n868), .B(\data_in<9> ), .C(n869), .D(\data_in<1> ), .Y(
        n870) );
  OAI21X1 U1195 ( .A(n3154), .B(n3532), .C(n557), .Y(n1994) );
  AOI22X1 U1196 ( .A(n868), .B(\data_in<10> ), .C(n869), .D(\data_in<2> ), .Y(
        n871) );
  OAI21X1 U1197 ( .A(n3154), .B(n3531), .C(n556), .Y(n1995) );
  AOI22X1 U1198 ( .A(n868), .B(\data_in<11> ), .C(n869), .D(\data_in<3> ), .Y(
        n872) );
  OAI21X1 U1199 ( .A(n3154), .B(n3530), .C(n555), .Y(n1996) );
  AOI22X1 U1200 ( .A(n868), .B(\data_in<12> ), .C(n869), .D(\data_in<4> ), .Y(
        n873) );
  OAI21X1 U1201 ( .A(n3154), .B(n3529), .C(n554), .Y(n1997) );
  AOI22X1 U1202 ( .A(n868), .B(\data_in<13> ), .C(n869), .D(\data_in<5> ), .Y(
        n874) );
  OAI21X1 U1203 ( .A(n3154), .B(n3528), .C(n553), .Y(n1998) );
  AOI22X1 U1204 ( .A(n868), .B(\data_in<14> ), .C(n869), .D(\data_in<6> ), .Y(
        n875) );
  OAI21X1 U1205 ( .A(n3154), .B(n3527), .C(n552), .Y(n1999) );
  AOI22X1 U1206 ( .A(n868), .B(\data_in<15> ), .C(n869), .D(\data_in<7> ), .Y(
        n876) );
  AOI21X1 U1207 ( .A(n2525), .B(n2520), .C(n3178), .Y(n866) );
  OAI21X1 U1208 ( .A(n3153), .B(n3526), .C(n551), .Y(n2000) );
  AOI22X1 U1209 ( .A(n880), .B(\data_in<8> ), .C(n881), .D(\data_in<0> ), .Y(
        n879) );
  OAI21X1 U1210 ( .A(n3153), .B(n3525), .C(n550), .Y(n2001) );
  AOI22X1 U1211 ( .A(n880), .B(\data_in<9> ), .C(n881), .D(\data_in<1> ), .Y(
        n882) );
  OAI21X1 U1212 ( .A(n3153), .B(n3524), .C(n549), .Y(n2002) );
  AOI22X1 U1213 ( .A(n880), .B(\data_in<10> ), .C(n881), .D(\data_in<2> ), .Y(
        n883) );
  OAI21X1 U1214 ( .A(n3153), .B(n3523), .C(n548), .Y(n2003) );
  AOI22X1 U1215 ( .A(n880), .B(\data_in<11> ), .C(n881), .D(\data_in<3> ), .Y(
        n884) );
  OAI21X1 U1216 ( .A(n3153), .B(n3522), .C(n547), .Y(n2004) );
  AOI22X1 U1217 ( .A(n880), .B(\data_in<12> ), .C(n881), .D(\data_in<4> ), .Y(
        n885) );
  OAI21X1 U1218 ( .A(n3153), .B(n3521), .C(n546), .Y(n2005) );
  AOI22X1 U1219 ( .A(n880), .B(\data_in<13> ), .C(n881), .D(\data_in<5> ), .Y(
        n886) );
  OAI21X1 U1220 ( .A(n3153), .B(n3520), .C(n545), .Y(n2006) );
  AOI22X1 U1221 ( .A(n880), .B(\data_in<14> ), .C(n881), .D(\data_in<6> ), .Y(
        n887) );
  OAI21X1 U1222 ( .A(n3153), .B(n3519), .C(n544), .Y(n2007) );
  AOI22X1 U1223 ( .A(n880), .B(\data_in<15> ), .C(n881), .D(\data_in<7> ), .Y(
        n888) );
  AOI21X1 U1224 ( .A(n2520), .B(n2521), .C(n3178), .Y(n878) );
  OAI21X1 U1225 ( .A(n3152), .B(n3518), .C(n543), .Y(n2008) );
  AOI22X1 U1226 ( .A(n892), .B(\data_in<8> ), .C(n893), .D(\data_in<0> ), .Y(
        n891) );
  OAI21X1 U1227 ( .A(n3152), .B(n3517), .C(n542), .Y(n2009) );
  AOI22X1 U1228 ( .A(n892), .B(\data_in<9> ), .C(n893), .D(\data_in<1> ), .Y(
        n894) );
  OAI21X1 U1229 ( .A(n3152), .B(n3516), .C(n541), .Y(n2010) );
  AOI22X1 U1230 ( .A(n892), .B(\data_in<10> ), .C(n893), .D(\data_in<2> ), .Y(
        n895) );
  OAI21X1 U1231 ( .A(n3152), .B(n3515), .C(n540), .Y(n2011) );
  AOI22X1 U1232 ( .A(n892), .B(\data_in<11> ), .C(n893), .D(\data_in<3> ), .Y(
        n896) );
  OAI21X1 U1233 ( .A(n3152), .B(n3514), .C(n539), .Y(n2012) );
  AOI22X1 U1234 ( .A(n892), .B(\data_in<12> ), .C(n893), .D(\data_in<4> ), .Y(
        n897) );
  OAI21X1 U1235 ( .A(n3152), .B(n3513), .C(n538), .Y(n2013) );
  AOI22X1 U1236 ( .A(n892), .B(\data_in<13> ), .C(n893), .D(\data_in<5> ), .Y(
        n898) );
  OAI21X1 U1237 ( .A(n3152), .B(n3512), .C(n537), .Y(n2014) );
  AOI22X1 U1238 ( .A(n892), .B(\data_in<14> ), .C(n893), .D(\data_in<6> ), .Y(
        n899) );
  OAI21X1 U1239 ( .A(n3152), .B(n3511), .C(n536), .Y(n2015) );
  AOI22X1 U1240 ( .A(n892), .B(\data_in<15> ), .C(n893), .D(\data_in<7> ), .Y(
        n900) );
  AOI21X1 U1241 ( .A(n2521), .B(n2548), .C(n3178), .Y(n890) );
  OAI21X1 U1242 ( .A(n3151), .B(n3510), .C(n535), .Y(n2016) );
  AOI22X1 U1243 ( .A(n904), .B(\data_in<8> ), .C(n905), .D(\data_in<0> ), .Y(
        n903) );
  OAI21X1 U1244 ( .A(n3151), .B(n3509), .C(n534), .Y(n2017) );
  AOI22X1 U1245 ( .A(n904), .B(\data_in<9> ), .C(n905), .D(\data_in<1> ), .Y(
        n906) );
  OAI21X1 U1246 ( .A(n3151), .B(n3508), .C(n533), .Y(n2018) );
  AOI22X1 U1247 ( .A(n904), .B(\data_in<10> ), .C(n905), .D(\data_in<2> ), .Y(
        n907) );
  OAI21X1 U1248 ( .A(n3151), .B(n3507), .C(n532), .Y(n2019) );
  AOI22X1 U1249 ( .A(n904), .B(\data_in<11> ), .C(n905), .D(\data_in<3> ), .Y(
        n908) );
  OAI21X1 U1250 ( .A(n3151), .B(n3506), .C(n531), .Y(n2020) );
  AOI22X1 U1251 ( .A(n904), .B(\data_in<12> ), .C(n905), .D(\data_in<4> ), .Y(
        n909) );
  OAI21X1 U1252 ( .A(n3151), .B(n3505), .C(n530), .Y(n2021) );
  AOI22X1 U1253 ( .A(n904), .B(\data_in<13> ), .C(n905), .D(\data_in<5> ), .Y(
        n910) );
  OAI21X1 U1254 ( .A(n3151), .B(n3504), .C(n529), .Y(n2022) );
  AOI22X1 U1255 ( .A(n904), .B(\data_in<14> ), .C(n905), .D(\data_in<6> ), .Y(
        n911) );
  OAI21X1 U1256 ( .A(n3151), .B(n3503), .C(n528), .Y(n2023) );
  AOI22X1 U1257 ( .A(n904), .B(\data_in<15> ), .C(n905), .D(\data_in<7> ), .Y(
        n912) );
  AOI21X1 U1258 ( .A(n2548), .B(n2549), .C(n3178), .Y(n902) );
  OAI21X1 U1259 ( .A(n3150), .B(n3502), .C(n527), .Y(n2024) );
  AOI22X1 U1260 ( .A(n916), .B(\data_in<8> ), .C(n917), .D(\data_in<0> ), .Y(
        n915) );
  OAI21X1 U1261 ( .A(n3150), .B(n3501), .C(n526), .Y(n2025) );
  AOI22X1 U1262 ( .A(n916), .B(\data_in<9> ), .C(n917), .D(\data_in<1> ), .Y(
        n918) );
  OAI21X1 U1263 ( .A(n3150), .B(n3500), .C(n525), .Y(n2026) );
  AOI22X1 U1264 ( .A(n916), .B(\data_in<10> ), .C(n917), .D(\data_in<2> ), .Y(
        n919) );
  OAI21X1 U1265 ( .A(n3150), .B(n3499), .C(n524), .Y(n2027) );
  AOI22X1 U1266 ( .A(n916), .B(\data_in<11> ), .C(n917), .D(\data_in<3> ), .Y(
        n920) );
  OAI21X1 U1267 ( .A(n3150), .B(n3498), .C(n523), .Y(n2028) );
  AOI22X1 U1268 ( .A(n916), .B(\data_in<12> ), .C(n917), .D(\data_in<4> ), .Y(
        n921) );
  OAI21X1 U1269 ( .A(n3150), .B(n3497), .C(n522), .Y(n2029) );
  AOI22X1 U1270 ( .A(n916), .B(\data_in<13> ), .C(n917), .D(\data_in<5> ), .Y(
        n922) );
  OAI21X1 U1271 ( .A(n3150), .B(n3496), .C(n521), .Y(n2030) );
  AOI22X1 U1272 ( .A(n916), .B(\data_in<14> ), .C(n917), .D(\data_in<6> ), .Y(
        n923) );
  OAI21X1 U1273 ( .A(n3150), .B(n3495), .C(n520), .Y(n2031) );
  AOI22X1 U1274 ( .A(n916), .B(\data_in<15> ), .C(n917), .D(\data_in<7> ), .Y(
        n924) );
  AOI21X1 U1275 ( .A(n2549), .B(n2544), .C(n3178), .Y(n914) );
  OAI21X1 U1276 ( .A(n3149), .B(n3494), .C(n519), .Y(n2032) );
  AOI22X1 U1277 ( .A(n928), .B(\data_in<8> ), .C(n929), .D(\data_in<0> ), .Y(
        n927) );
  OAI21X1 U1278 ( .A(n3149), .B(n3493), .C(n518), .Y(n2033) );
  AOI22X1 U1279 ( .A(n928), .B(\data_in<9> ), .C(n929), .D(\data_in<1> ), .Y(
        n930) );
  OAI21X1 U1280 ( .A(n3149), .B(n3492), .C(n517), .Y(n2034) );
  AOI22X1 U1281 ( .A(n928), .B(\data_in<10> ), .C(n929), .D(\data_in<2> ), .Y(
        n931) );
  OAI21X1 U1282 ( .A(n3149), .B(n3491), .C(n516), .Y(n2035) );
  AOI22X1 U1283 ( .A(n928), .B(\data_in<11> ), .C(n929), .D(\data_in<3> ), .Y(
        n932) );
  OAI21X1 U1284 ( .A(n3149), .B(n3490), .C(n515), .Y(n2036) );
  AOI22X1 U1285 ( .A(n928), .B(\data_in<12> ), .C(n929), .D(\data_in<4> ), .Y(
        n933) );
  OAI21X1 U1286 ( .A(n3149), .B(n3489), .C(n514), .Y(n2037) );
  AOI22X1 U1287 ( .A(n928), .B(\data_in<13> ), .C(n929), .D(\data_in<5> ), .Y(
        n934) );
  OAI21X1 U1288 ( .A(n3149), .B(n3488), .C(n513), .Y(n2038) );
  AOI22X1 U1289 ( .A(n928), .B(\data_in<14> ), .C(n929), .D(\data_in<6> ), .Y(
        n935) );
  OAI21X1 U1290 ( .A(n3149), .B(n3487), .C(n512), .Y(n2039) );
  AOI22X1 U1291 ( .A(n928), .B(\data_in<15> ), .C(n929), .D(\data_in<7> ), .Y(
        n936) );
  AOI21X1 U1292 ( .A(n2544), .B(n2545), .C(n3178), .Y(n926) );
  OAI21X1 U1293 ( .A(n3148), .B(n3486), .C(n511), .Y(n2040) );
  AOI22X1 U1294 ( .A(n940), .B(\data_in<8> ), .C(n941), .D(\data_in<0> ), .Y(
        n939) );
  OAI21X1 U1295 ( .A(n3148), .B(n3485), .C(n510), .Y(n2041) );
  AOI22X1 U1296 ( .A(n940), .B(\data_in<9> ), .C(n941), .D(\data_in<1> ), .Y(
        n942) );
  OAI21X1 U1297 ( .A(n3148), .B(n3484), .C(n509), .Y(n2042) );
  AOI22X1 U1298 ( .A(n940), .B(\data_in<10> ), .C(n941), .D(\data_in<2> ), .Y(
        n943) );
  OAI21X1 U1299 ( .A(n3148), .B(n3483), .C(n508), .Y(n2043) );
  AOI22X1 U1300 ( .A(n940), .B(\data_in<11> ), .C(n941), .D(\data_in<3> ), .Y(
        n944) );
  OAI21X1 U1301 ( .A(n3148), .B(n3482), .C(n507), .Y(n2044) );
  AOI22X1 U1302 ( .A(n940), .B(\data_in<12> ), .C(n941), .D(\data_in<4> ), .Y(
        n945) );
  OAI21X1 U1303 ( .A(n3148), .B(n3481), .C(n506), .Y(n2045) );
  AOI22X1 U1304 ( .A(n940), .B(\data_in<13> ), .C(n941), .D(\data_in<5> ), .Y(
        n946) );
  OAI21X1 U1305 ( .A(n3148), .B(n3480), .C(n505), .Y(n2046) );
  AOI22X1 U1306 ( .A(n940), .B(\data_in<14> ), .C(n941), .D(\data_in<6> ), .Y(
        n947) );
  OAI21X1 U1307 ( .A(n3148), .B(n3479), .C(n504), .Y(n2047) );
  AOI22X1 U1308 ( .A(n940), .B(\data_in<15> ), .C(n941), .D(\data_in<7> ), .Y(
        n948) );
  AOI21X1 U1309 ( .A(n2545), .B(n2540), .C(n3178), .Y(n938) );
  OAI21X1 U1310 ( .A(n3147), .B(n3478), .C(n503), .Y(n2048) );
  AOI22X1 U1311 ( .A(n952), .B(\data_in<8> ), .C(n953), .D(\data_in<0> ), .Y(
        n951) );
  OAI21X1 U1312 ( .A(n3147), .B(n3477), .C(n502), .Y(n2049) );
  AOI22X1 U1313 ( .A(n952), .B(\data_in<9> ), .C(n953), .D(\data_in<1> ), .Y(
        n954) );
  OAI21X1 U1314 ( .A(n3147), .B(n3476), .C(n501), .Y(n2050) );
  AOI22X1 U1315 ( .A(n952), .B(\data_in<10> ), .C(n953), .D(\data_in<2> ), .Y(
        n955) );
  OAI21X1 U1316 ( .A(n3147), .B(n3475), .C(n500), .Y(n2051) );
  AOI22X1 U1317 ( .A(n952), .B(\data_in<11> ), .C(n953), .D(\data_in<3> ), .Y(
        n956) );
  OAI21X1 U1318 ( .A(n3147), .B(n3474), .C(n499), .Y(n2052) );
  AOI22X1 U1319 ( .A(n952), .B(\data_in<12> ), .C(n953), .D(\data_in<4> ), .Y(
        n957) );
  OAI21X1 U1320 ( .A(n3147), .B(n3473), .C(n498), .Y(n2053) );
  AOI22X1 U1321 ( .A(n952), .B(\data_in<13> ), .C(n953), .D(\data_in<5> ), .Y(
        n958) );
  OAI21X1 U1322 ( .A(n3147), .B(n3472), .C(n497), .Y(n2054) );
  AOI22X1 U1323 ( .A(n952), .B(\data_in<14> ), .C(n953), .D(\data_in<6> ), .Y(
        n959) );
  OAI21X1 U1324 ( .A(n3147), .B(n3471), .C(n496), .Y(n2055) );
  AOI22X1 U1325 ( .A(n952), .B(\data_in<15> ), .C(n953), .D(\data_in<7> ), .Y(
        n960) );
  AOI21X1 U1326 ( .A(n2540), .B(n2541), .C(n3178), .Y(n950) );
  OAI21X1 U1327 ( .A(n3146), .B(n3470), .C(n495), .Y(n2056) );
  AOI22X1 U1328 ( .A(n964), .B(\data_in<8> ), .C(n965), .D(\data_in<0> ), .Y(
        n963) );
  OAI21X1 U1329 ( .A(n3146), .B(n3469), .C(n494), .Y(n2057) );
  AOI22X1 U1330 ( .A(n964), .B(\data_in<9> ), .C(n965), .D(\data_in<1> ), .Y(
        n966) );
  OAI21X1 U1331 ( .A(n3146), .B(n3468), .C(n493), .Y(n2058) );
  AOI22X1 U1332 ( .A(n964), .B(\data_in<10> ), .C(n965), .D(\data_in<2> ), .Y(
        n967) );
  OAI21X1 U1333 ( .A(n3146), .B(n3467), .C(n492), .Y(n2059) );
  AOI22X1 U1334 ( .A(n964), .B(\data_in<11> ), .C(n965), .D(\data_in<3> ), .Y(
        n968) );
  OAI21X1 U1335 ( .A(n3146), .B(n3466), .C(n491), .Y(n2060) );
  AOI22X1 U1336 ( .A(n964), .B(\data_in<12> ), .C(n965), .D(\data_in<4> ), .Y(
        n969) );
  OAI21X1 U1337 ( .A(n3146), .B(n3465), .C(n490), .Y(n2061) );
  AOI22X1 U1338 ( .A(n964), .B(\data_in<13> ), .C(n965), .D(\data_in<5> ), .Y(
        n970) );
  OAI21X1 U1339 ( .A(n3146), .B(n3464), .C(n489), .Y(n2062) );
  AOI22X1 U1340 ( .A(n964), .B(\data_in<14> ), .C(n965), .D(\data_in<6> ), .Y(
        n971) );
  OAI21X1 U1341 ( .A(n3146), .B(n3463), .C(n488), .Y(n2063) );
  AOI22X1 U1342 ( .A(n964), .B(\data_in<15> ), .C(n965), .D(\data_in<7> ), .Y(
        n972) );
  AOI21X1 U1343 ( .A(n2541), .B(n2535), .C(n3178), .Y(n962) );
  OAI21X1 U1344 ( .A(n3145), .B(n3462), .C(n487), .Y(n2064) );
  AOI22X1 U1345 ( .A(n976), .B(\data_in<8> ), .C(n977), .D(\data_in<0> ), .Y(
        n975) );
  OAI21X1 U1346 ( .A(n3145), .B(n3461), .C(n486), .Y(n2065) );
  AOI22X1 U1347 ( .A(n976), .B(\data_in<9> ), .C(n977), .D(\data_in<1> ), .Y(
        n978) );
  OAI21X1 U1348 ( .A(n3145), .B(n3460), .C(n485), .Y(n2066) );
  AOI22X1 U1349 ( .A(n976), .B(\data_in<10> ), .C(n977), .D(\data_in<2> ), .Y(
        n979) );
  OAI21X1 U1350 ( .A(n3145), .B(n3459), .C(n484), .Y(n2067) );
  AOI22X1 U1351 ( .A(n976), .B(\data_in<11> ), .C(n977), .D(\data_in<3> ), .Y(
        n980) );
  OAI21X1 U1352 ( .A(n3145), .B(n3458), .C(n483), .Y(n2068) );
  AOI22X1 U1353 ( .A(n976), .B(\data_in<12> ), .C(n977), .D(\data_in<4> ), .Y(
        n981) );
  OAI21X1 U1354 ( .A(n3145), .B(n3457), .C(n482), .Y(n2069) );
  AOI22X1 U1355 ( .A(n976), .B(\data_in<13> ), .C(n977), .D(\data_in<5> ), .Y(
        n982) );
  OAI21X1 U1356 ( .A(n3145), .B(n3456), .C(n481), .Y(n2070) );
  AOI22X1 U1357 ( .A(n976), .B(\data_in<14> ), .C(n977), .D(\data_in<6> ), .Y(
        n983) );
  OAI21X1 U1358 ( .A(n3145), .B(n3455), .C(n480), .Y(n2071) );
  AOI22X1 U1359 ( .A(n976), .B(\data_in<15> ), .C(n977), .D(\data_in<7> ), .Y(
        n984) );
  AOI21X1 U1360 ( .A(n2535), .B(n2538), .C(n3178), .Y(n974) );
  OAI21X1 U1361 ( .A(n3144), .B(n3454), .C(n479), .Y(n2072) );
  AOI22X1 U1362 ( .A(n988), .B(\data_in<8> ), .C(n989), .D(\data_in<0> ), .Y(
        n987) );
  OAI21X1 U1363 ( .A(n3144), .B(n3453), .C(n478), .Y(n2073) );
  AOI22X1 U1364 ( .A(n988), .B(\data_in<9> ), .C(n989), .D(\data_in<1> ), .Y(
        n990) );
  OAI21X1 U1365 ( .A(n3144), .B(n3452), .C(n477), .Y(n2074) );
  AOI22X1 U1366 ( .A(n988), .B(\data_in<10> ), .C(n989), .D(\data_in<2> ), .Y(
        n991) );
  OAI21X1 U1367 ( .A(n3144), .B(n3451), .C(n476), .Y(n2075) );
  AOI22X1 U1368 ( .A(n988), .B(\data_in<11> ), .C(n989), .D(\data_in<3> ), .Y(
        n992) );
  OAI21X1 U1369 ( .A(n3144), .B(n3450), .C(n475), .Y(n2076) );
  AOI22X1 U1370 ( .A(n988), .B(\data_in<12> ), .C(n989), .D(\data_in<4> ), .Y(
        n993) );
  OAI21X1 U1371 ( .A(n3144), .B(n3449), .C(n474), .Y(n2077) );
  AOI22X1 U1372 ( .A(n988), .B(\data_in<13> ), .C(n989), .D(\data_in<5> ), .Y(
        n994) );
  OAI21X1 U1373 ( .A(n3144), .B(n3448), .C(n473), .Y(n2078) );
  AOI22X1 U1374 ( .A(n988), .B(\data_in<14> ), .C(n989), .D(\data_in<6> ), .Y(
        n995) );
  OAI21X1 U1375 ( .A(n3144), .B(n3447), .C(n472), .Y(n2079) );
  AOI22X1 U1376 ( .A(n988), .B(\data_in<15> ), .C(n989), .D(\data_in<7> ), .Y(
        n996) );
  AOI21X1 U1377 ( .A(n2538), .B(n2474), .C(n3178), .Y(n986) );
  OAI21X1 U1378 ( .A(n3143), .B(n3446), .C(n471), .Y(n2080) );
  AOI22X1 U1379 ( .A(n1000), .B(\data_in<8> ), .C(n1001), .D(\data_in<0> ), 
        .Y(n999) );
  OAI21X1 U1380 ( .A(n3143), .B(n3445), .C(n470), .Y(n2081) );
  AOI22X1 U1381 ( .A(n1000), .B(\data_in<9> ), .C(n1001), .D(\data_in<1> ), 
        .Y(n1002) );
  OAI21X1 U1382 ( .A(n3143), .B(n3444), .C(n469), .Y(n2082) );
  AOI22X1 U1383 ( .A(n1000), .B(\data_in<10> ), .C(n1001), .D(\data_in<2> ), 
        .Y(n1003) );
  OAI21X1 U1384 ( .A(n3143), .B(n3443), .C(n468), .Y(n2083) );
  AOI22X1 U1385 ( .A(n1000), .B(\data_in<11> ), .C(n1001), .D(\data_in<3> ), 
        .Y(n1004) );
  OAI21X1 U1386 ( .A(n3143), .B(n3442), .C(n467), .Y(n2084) );
  AOI22X1 U1387 ( .A(n1000), .B(\data_in<12> ), .C(n1001), .D(\data_in<4> ), 
        .Y(n1005) );
  OAI21X1 U1388 ( .A(n3143), .B(n3441), .C(n466), .Y(n2085) );
  AOI22X1 U1389 ( .A(n1000), .B(\data_in<13> ), .C(n1001), .D(\data_in<5> ), 
        .Y(n1006) );
  OAI21X1 U1390 ( .A(n3143), .B(n3440), .C(n465), .Y(n2086) );
  AOI22X1 U1391 ( .A(n1000), .B(\data_in<14> ), .C(n1001), .D(\data_in<6> ), 
        .Y(n1007) );
  OAI21X1 U1392 ( .A(n3143), .B(n3439), .C(n464), .Y(n2087) );
  AOI22X1 U1393 ( .A(n1000), .B(\data_in<15> ), .C(n1001), .D(\data_in<7> ), 
        .Y(n1008) );
  AOI21X1 U1394 ( .A(n2474), .B(n2475), .C(n3178), .Y(n998) );
  OAI21X1 U1395 ( .A(n3142), .B(n3438), .C(n463), .Y(n2088) );
  AOI22X1 U1396 ( .A(n1012), .B(\data_in<8> ), .C(n1013), .D(\data_in<0> ), 
        .Y(n1011) );
  OAI21X1 U1397 ( .A(n3142), .B(n3437), .C(n462), .Y(n2089) );
  AOI22X1 U1398 ( .A(n1012), .B(\data_in<9> ), .C(n1013), .D(\data_in<1> ), 
        .Y(n1014) );
  OAI21X1 U1399 ( .A(n3142), .B(n3436), .C(n461), .Y(n2090) );
  AOI22X1 U1400 ( .A(n1012), .B(\data_in<10> ), .C(n1013), .D(\data_in<2> ), 
        .Y(n1015) );
  OAI21X1 U1401 ( .A(n3142), .B(n3435), .C(n460), .Y(n2091) );
  AOI22X1 U1402 ( .A(n1012), .B(\data_in<11> ), .C(n1013), .D(\data_in<3> ), 
        .Y(n1016) );
  OAI21X1 U1403 ( .A(n3142), .B(n3434), .C(n459), .Y(n2092) );
  AOI22X1 U1404 ( .A(n1012), .B(\data_in<12> ), .C(n1013), .D(\data_in<4> ), 
        .Y(n1017) );
  OAI21X1 U1405 ( .A(n3142), .B(n3433), .C(n458), .Y(n2093) );
  AOI22X1 U1406 ( .A(n1012), .B(\data_in<13> ), .C(n1013), .D(\data_in<5> ), 
        .Y(n1018) );
  OAI21X1 U1407 ( .A(n3142), .B(n3432), .C(n457), .Y(n2094) );
  AOI22X1 U1408 ( .A(n1012), .B(\data_in<14> ), .C(n1013), .D(\data_in<6> ), 
        .Y(n1019) );
  OAI21X1 U1409 ( .A(n3142), .B(n3431), .C(n456), .Y(n2095) );
  AOI22X1 U1410 ( .A(n1012), .B(\data_in<15> ), .C(n1013), .D(\data_in<7> ), 
        .Y(n1020) );
  AOI21X1 U1411 ( .A(n2475), .B(n2470), .C(n3178), .Y(n1010) );
  OAI21X1 U1412 ( .A(n3141), .B(n3430), .C(n455), .Y(n2096) );
  AOI22X1 U1413 ( .A(n1024), .B(\data_in<8> ), .C(n1025), .D(\data_in<0> ), 
        .Y(n1023) );
  OAI21X1 U1414 ( .A(n3141), .B(n3429), .C(n454), .Y(n2097) );
  AOI22X1 U1415 ( .A(n1024), .B(\data_in<9> ), .C(n1025), .D(\data_in<1> ), 
        .Y(n1026) );
  OAI21X1 U1416 ( .A(n3141), .B(n3428), .C(n453), .Y(n2098) );
  AOI22X1 U1417 ( .A(n1024), .B(\data_in<10> ), .C(n1025), .D(\data_in<2> ), 
        .Y(n1027) );
  OAI21X1 U1418 ( .A(n3141), .B(n3427), .C(n452), .Y(n2099) );
  AOI22X1 U1419 ( .A(n1024), .B(\data_in<11> ), .C(n1025), .D(\data_in<3> ), 
        .Y(n1028) );
  OAI21X1 U1420 ( .A(n3141), .B(n3426), .C(n451), .Y(n2100) );
  AOI22X1 U1421 ( .A(n1024), .B(\data_in<12> ), .C(n1025), .D(\data_in<4> ), 
        .Y(n1029) );
  OAI21X1 U1422 ( .A(n3141), .B(n3425), .C(n450), .Y(n2101) );
  AOI22X1 U1423 ( .A(n1024), .B(\data_in<13> ), .C(n1025), .D(\data_in<5> ), 
        .Y(n1030) );
  OAI21X1 U1424 ( .A(n3141), .B(n3424), .C(n449), .Y(n2102) );
  AOI22X1 U1425 ( .A(n1024), .B(\data_in<14> ), .C(n1025), .D(\data_in<6> ), 
        .Y(n1031) );
  OAI21X1 U1426 ( .A(n3141), .B(n3423), .C(n448), .Y(n2103) );
  AOI22X1 U1427 ( .A(n1024), .B(\data_in<15> ), .C(n1025), .D(\data_in<7> ), 
        .Y(n1032) );
  AOI21X1 U1428 ( .A(n2470), .B(n2471), .C(n3177), .Y(n1022) );
  OAI21X1 U1429 ( .A(n3140), .B(n3422), .C(n447), .Y(n2104) );
  AOI22X1 U1430 ( .A(n1036), .B(\data_in<8> ), .C(n1037), .D(\data_in<0> ), 
        .Y(n1035) );
  OAI21X1 U1431 ( .A(n3140), .B(n3421), .C(n446), .Y(n2105) );
  AOI22X1 U1432 ( .A(n1036), .B(\data_in<9> ), .C(n1037), .D(\data_in<1> ), 
        .Y(n1038) );
  OAI21X1 U1433 ( .A(n3140), .B(n3420), .C(n445), .Y(n2106) );
  AOI22X1 U1434 ( .A(n1036), .B(\data_in<10> ), .C(n1037), .D(\data_in<2> ), 
        .Y(n1039) );
  OAI21X1 U1435 ( .A(n3140), .B(n3419), .C(n444), .Y(n2107) );
  AOI22X1 U1436 ( .A(n1036), .B(\data_in<11> ), .C(n1037), .D(\data_in<3> ), 
        .Y(n1040) );
  OAI21X1 U1437 ( .A(n3140), .B(n3418), .C(n443), .Y(n2108) );
  AOI22X1 U1438 ( .A(n1036), .B(\data_in<12> ), .C(n1037), .D(\data_in<4> ), 
        .Y(n1041) );
  OAI21X1 U1439 ( .A(n3140), .B(n3417), .C(n442), .Y(n2109) );
  AOI22X1 U1440 ( .A(n1036), .B(\data_in<13> ), .C(n1037), .D(\data_in<5> ), 
        .Y(n1042) );
  OAI21X1 U1441 ( .A(n3140), .B(n3416), .C(n441), .Y(n2110) );
  AOI22X1 U1442 ( .A(n1036), .B(\data_in<14> ), .C(n1037), .D(\data_in<6> ), 
        .Y(n1043) );
  OAI21X1 U1443 ( .A(n3140), .B(n3415), .C(n440), .Y(n2111) );
  AOI22X1 U1444 ( .A(n1036), .B(\data_in<15> ), .C(n1037), .D(\data_in<7> ), 
        .Y(n1044) );
  AOI21X1 U1445 ( .A(n2471), .B(n2466), .C(n3177), .Y(n1034) );
  OAI21X1 U1446 ( .A(n3139), .B(n3414), .C(n439), .Y(n2112) );
  AOI22X1 U1447 ( .A(n1048), .B(\data_in<8> ), .C(n1049), .D(\data_in<0> ), 
        .Y(n1047) );
  OAI21X1 U1448 ( .A(n3139), .B(n3413), .C(n438), .Y(n2113) );
  AOI22X1 U1449 ( .A(n1048), .B(\data_in<9> ), .C(n1049), .D(\data_in<1> ), 
        .Y(n1050) );
  OAI21X1 U1450 ( .A(n3139), .B(n3412), .C(n437), .Y(n2114) );
  AOI22X1 U1451 ( .A(n1048), .B(\data_in<10> ), .C(n1049), .D(\data_in<2> ), 
        .Y(n1051) );
  OAI21X1 U1452 ( .A(n3139), .B(n3411), .C(n436), .Y(n2115) );
  AOI22X1 U1453 ( .A(n1048), .B(\data_in<11> ), .C(n1049), .D(\data_in<3> ), 
        .Y(n1052) );
  OAI21X1 U1454 ( .A(n3139), .B(n3410), .C(n435), .Y(n2116) );
  AOI22X1 U1455 ( .A(n1048), .B(\data_in<12> ), .C(n1049), .D(\data_in<4> ), 
        .Y(n1053) );
  OAI21X1 U1456 ( .A(n3139), .B(n3409), .C(n434), .Y(n2117) );
  AOI22X1 U1457 ( .A(n1048), .B(\data_in<13> ), .C(n1049), .D(\data_in<5> ), 
        .Y(n1054) );
  OAI21X1 U1458 ( .A(n3139), .B(n3408), .C(n433), .Y(n2118) );
  AOI22X1 U1459 ( .A(n1048), .B(\data_in<14> ), .C(n1049), .D(\data_in<6> ), 
        .Y(n1055) );
  OAI21X1 U1460 ( .A(n3139), .B(n3407), .C(n432), .Y(n2119) );
  AOI22X1 U1461 ( .A(n1048), .B(\data_in<15> ), .C(n1049), .D(\data_in<7> ), 
        .Y(n1056) );
  AOI21X1 U1462 ( .A(n2466), .B(n2467), .C(n3177), .Y(n1046) );
  OAI21X1 U1463 ( .A(n3138), .B(n3406), .C(n431), .Y(n2120) );
  AOI22X1 U1464 ( .A(n1060), .B(\data_in<8> ), .C(n1061), .D(\data_in<0> ), 
        .Y(n1059) );
  OAI21X1 U1465 ( .A(n3138), .B(n3405), .C(n430), .Y(n2121) );
  AOI22X1 U1466 ( .A(n1060), .B(\data_in<9> ), .C(n1061), .D(\data_in<1> ), 
        .Y(n1062) );
  OAI21X1 U1467 ( .A(n3138), .B(n3404), .C(n429), .Y(n2122) );
  AOI22X1 U1468 ( .A(n1060), .B(\data_in<10> ), .C(n1061), .D(\data_in<2> ), 
        .Y(n1063) );
  OAI21X1 U1469 ( .A(n3138), .B(n3403), .C(n428), .Y(n2123) );
  AOI22X1 U1470 ( .A(n1060), .B(\data_in<11> ), .C(n1061), .D(\data_in<3> ), 
        .Y(n1064) );
  OAI21X1 U1471 ( .A(n3138), .B(n3402), .C(n427), .Y(n2124) );
  AOI22X1 U1472 ( .A(n1060), .B(\data_in<12> ), .C(n1061), .D(\data_in<4> ), 
        .Y(n1065) );
  OAI21X1 U1473 ( .A(n3138), .B(n3401), .C(n426), .Y(n2125) );
  AOI22X1 U1474 ( .A(n1060), .B(\data_in<13> ), .C(n1061), .D(\data_in<5> ), 
        .Y(n1066) );
  OAI21X1 U1475 ( .A(n3138), .B(n3400), .C(n425), .Y(n2126) );
  AOI22X1 U1476 ( .A(n1060), .B(\data_in<14> ), .C(n1061), .D(\data_in<6> ), 
        .Y(n1067) );
  OAI21X1 U1477 ( .A(n3138), .B(n3399), .C(n424), .Y(n2127) );
  AOI22X1 U1478 ( .A(n1060), .B(\data_in<15> ), .C(n1061), .D(\data_in<7> ), 
        .Y(n1068) );
  AOI21X1 U1479 ( .A(n2467), .B(n2462), .C(n3177), .Y(n1058) );
  OAI21X1 U1480 ( .A(n3137), .B(n3398), .C(n423), .Y(n2128) );
  AOI22X1 U1481 ( .A(n1072), .B(\data_in<8> ), .C(n1073), .D(\data_in<0> ), 
        .Y(n1071) );
  OAI21X1 U1482 ( .A(n3137), .B(n3397), .C(n422), .Y(n2129) );
  AOI22X1 U1483 ( .A(n1072), .B(\data_in<9> ), .C(n1073), .D(\data_in<1> ), 
        .Y(n1074) );
  OAI21X1 U1484 ( .A(n3137), .B(n3396), .C(n421), .Y(n2130) );
  AOI22X1 U1485 ( .A(n1072), .B(\data_in<10> ), .C(n1073), .D(\data_in<2> ), 
        .Y(n1075) );
  OAI21X1 U1486 ( .A(n3137), .B(n3395), .C(n420), .Y(n2131) );
  AOI22X1 U1487 ( .A(n1072), .B(\data_in<11> ), .C(n1073), .D(\data_in<3> ), 
        .Y(n1076) );
  OAI21X1 U1488 ( .A(n3137), .B(n3394), .C(n419), .Y(n2132) );
  AOI22X1 U1489 ( .A(n1072), .B(\data_in<12> ), .C(n1073), .D(\data_in<4> ), 
        .Y(n1077) );
  OAI21X1 U1490 ( .A(n3137), .B(n3393), .C(n418), .Y(n2133) );
  AOI22X1 U1491 ( .A(n1072), .B(\data_in<13> ), .C(n1073), .D(\data_in<5> ), 
        .Y(n1078) );
  OAI21X1 U1492 ( .A(n3137), .B(n3392), .C(n417), .Y(n2134) );
  AOI22X1 U1493 ( .A(n1072), .B(\data_in<14> ), .C(n1073), .D(\data_in<6> ), 
        .Y(n1079) );
  OAI21X1 U1494 ( .A(n3137), .B(n3391), .C(n416), .Y(n2135) );
  AOI22X1 U1495 ( .A(n1072), .B(\data_in<15> ), .C(n1073), .D(\data_in<7> ), 
        .Y(n1080) );
  AOI21X1 U1496 ( .A(n2462), .B(n2463), .C(n3177), .Y(n1070) );
  OAI21X1 U1497 ( .A(n3136), .B(n3390), .C(n415), .Y(n2136) );
  AOI22X1 U1498 ( .A(n1084), .B(\data_in<8> ), .C(n1085), .D(\data_in<0> ), 
        .Y(n1083) );
  OAI21X1 U1499 ( .A(n3136), .B(n3389), .C(n414), .Y(n2137) );
  AOI22X1 U1500 ( .A(n1084), .B(\data_in<9> ), .C(n1085), .D(\data_in<1> ), 
        .Y(n1086) );
  OAI21X1 U1501 ( .A(n3136), .B(n3388), .C(n413), .Y(n2138) );
  AOI22X1 U1502 ( .A(n1084), .B(\data_in<10> ), .C(n1085), .D(\data_in<2> ), 
        .Y(n1087) );
  OAI21X1 U1503 ( .A(n3136), .B(n3387), .C(n412), .Y(n2139) );
  AOI22X1 U1504 ( .A(n1084), .B(\data_in<11> ), .C(n1085), .D(\data_in<3> ), 
        .Y(n1088) );
  OAI21X1 U1505 ( .A(n3136), .B(n3386), .C(n411), .Y(n2140) );
  AOI22X1 U1506 ( .A(n1084), .B(\data_in<12> ), .C(n1085), .D(\data_in<4> ), 
        .Y(n1089) );
  OAI21X1 U1507 ( .A(n3136), .B(n3385), .C(n410), .Y(n2141) );
  AOI22X1 U1508 ( .A(n1084), .B(\data_in<13> ), .C(n1085), .D(\data_in<5> ), 
        .Y(n1090) );
  OAI21X1 U1509 ( .A(n3136), .B(n3384), .C(n409), .Y(n2142) );
  AOI22X1 U1510 ( .A(n1084), .B(\data_in<14> ), .C(n1085), .D(\data_in<6> ), 
        .Y(n1091) );
  OAI21X1 U1511 ( .A(n3136), .B(n3383), .C(n408), .Y(n2143) );
  AOI22X1 U1512 ( .A(n1084), .B(\data_in<15> ), .C(n1085), .D(\data_in<7> ), 
        .Y(n1092) );
  AOI21X1 U1513 ( .A(n2463), .B(n2490), .C(n3177), .Y(n1082) );
  OAI21X1 U1514 ( .A(n3135), .B(n3382), .C(n407), .Y(n2144) );
  AOI22X1 U1515 ( .A(n1096), .B(\data_in<8> ), .C(n1097), .D(\data_in<0> ), 
        .Y(n1095) );
  OAI21X1 U1516 ( .A(n3135), .B(n3381), .C(n406), .Y(n2145) );
  AOI22X1 U1517 ( .A(n1096), .B(\data_in<9> ), .C(n1097), .D(\data_in<1> ), 
        .Y(n1098) );
  OAI21X1 U1518 ( .A(n3135), .B(n3380), .C(n405), .Y(n2146) );
  AOI22X1 U1519 ( .A(n1096), .B(\data_in<10> ), .C(n1097), .D(\data_in<2> ), 
        .Y(n1099) );
  OAI21X1 U1520 ( .A(n3135), .B(n3379), .C(n404), .Y(n2147) );
  AOI22X1 U1521 ( .A(n1096), .B(\data_in<11> ), .C(n1097), .D(\data_in<3> ), 
        .Y(n1100) );
  OAI21X1 U1522 ( .A(n3135), .B(n3378), .C(n403), .Y(n2148) );
  AOI22X1 U1523 ( .A(n1096), .B(\data_in<12> ), .C(n1097), .D(\data_in<4> ), 
        .Y(n1101) );
  OAI21X1 U1524 ( .A(n3135), .B(n3377), .C(n402), .Y(n2149) );
  AOI22X1 U1525 ( .A(n1096), .B(\data_in<13> ), .C(n1097), .D(\data_in<5> ), 
        .Y(n1102) );
  OAI21X1 U1526 ( .A(n3135), .B(n3376), .C(n401), .Y(n2150) );
  AOI22X1 U1527 ( .A(n1096), .B(\data_in<14> ), .C(n1097), .D(\data_in<6> ), 
        .Y(n1103) );
  OAI21X1 U1528 ( .A(n3135), .B(n3375), .C(n400), .Y(n2151) );
  AOI22X1 U1529 ( .A(n1096), .B(\data_in<15> ), .C(n1097), .D(\data_in<7> ), 
        .Y(n1104) );
  AOI21X1 U1530 ( .A(n2490), .B(n2491), .C(n3177), .Y(n1094) );
  OAI21X1 U1531 ( .A(n3134), .B(n3374), .C(n399), .Y(n2152) );
  AOI22X1 U1532 ( .A(n1108), .B(\data_in<8> ), .C(n1109), .D(\data_in<0> ), 
        .Y(n1107) );
  OAI21X1 U1533 ( .A(n3134), .B(n3373), .C(n398), .Y(n2153) );
  AOI22X1 U1534 ( .A(n1108), .B(\data_in<9> ), .C(n1109), .D(\data_in<1> ), 
        .Y(n1110) );
  OAI21X1 U1535 ( .A(n3134), .B(n3372), .C(n397), .Y(n2154) );
  AOI22X1 U1536 ( .A(n1108), .B(\data_in<10> ), .C(n1109), .D(\data_in<2> ), 
        .Y(n1111) );
  OAI21X1 U1537 ( .A(n3134), .B(n3371), .C(n396), .Y(n2155) );
  AOI22X1 U1538 ( .A(n1108), .B(\data_in<11> ), .C(n1109), .D(\data_in<3> ), 
        .Y(n1112) );
  OAI21X1 U1539 ( .A(n3134), .B(n3370), .C(n395), .Y(n2156) );
  AOI22X1 U1540 ( .A(n1108), .B(\data_in<12> ), .C(n1109), .D(\data_in<4> ), 
        .Y(n1113) );
  OAI21X1 U1541 ( .A(n3134), .B(n3369), .C(n394), .Y(n2157) );
  AOI22X1 U1542 ( .A(n1108), .B(\data_in<13> ), .C(n1109), .D(\data_in<5> ), 
        .Y(n1114) );
  OAI21X1 U1543 ( .A(n3134), .B(n3368), .C(n393), .Y(n2158) );
  AOI22X1 U1544 ( .A(n1108), .B(\data_in<14> ), .C(n1109), .D(\data_in<6> ), 
        .Y(n1115) );
  OAI21X1 U1545 ( .A(n3134), .B(n3367), .C(n392), .Y(n2159) );
  AOI22X1 U1546 ( .A(n1108), .B(\data_in<15> ), .C(n1109), .D(\data_in<7> ), 
        .Y(n1116) );
  AOI21X1 U1547 ( .A(n2491), .B(n2486), .C(n3177), .Y(n1106) );
  OAI21X1 U1548 ( .A(n3133), .B(n3366), .C(n391), .Y(n2160) );
  AOI22X1 U1549 ( .A(n1120), .B(\data_in<8> ), .C(n1121), .D(\data_in<0> ), 
        .Y(n1119) );
  OAI21X1 U1550 ( .A(n3133), .B(n3365), .C(n390), .Y(n2161) );
  AOI22X1 U1551 ( .A(n1120), .B(\data_in<9> ), .C(n1121), .D(\data_in<1> ), 
        .Y(n1122) );
  OAI21X1 U1552 ( .A(n3133), .B(n3364), .C(n389), .Y(n2162) );
  AOI22X1 U1553 ( .A(n1120), .B(\data_in<10> ), .C(n1121), .D(\data_in<2> ), 
        .Y(n1123) );
  OAI21X1 U1554 ( .A(n3133), .B(n3363), .C(n388), .Y(n2163) );
  AOI22X1 U1555 ( .A(n1120), .B(\data_in<11> ), .C(n1121), .D(\data_in<3> ), 
        .Y(n1124) );
  OAI21X1 U1556 ( .A(n3133), .B(n3362), .C(n387), .Y(n2164) );
  AOI22X1 U1557 ( .A(n1120), .B(\data_in<12> ), .C(n1121), .D(\data_in<4> ), 
        .Y(n1125) );
  OAI21X1 U1558 ( .A(n3133), .B(n3361), .C(n386), .Y(n2165) );
  AOI22X1 U1559 ( .A(n1120), .B(\data_in<13> ), .C(n1121), .D(\data_in<5> ), 
        .Y(n1126) );
  OAI21X1 U1560 ( .A(n3133), .B(n3360), .C(n385), .Y(n2166) );
  AOI22X1 U1561 ( .A(n1120), .B(\data_in<14> ), .C(n1121), .D(\data_in<6> ), 
        .Y(n1127) );
  OAI21X1 U1562 ( .A(n3133), .B(n3359), .C(n384), .Y(n2167) );
  AOI22X1 U1563 ( .A(n1120), .B(\data_in<15> ), .C(n1121), .D(\data_in<7> ), 
        .Y(n1128) );
  AOI21X1 U1564 ( .A(n2486), .B(n2487), .C(n3177), .Y(n1118) );
  OAI21X1 U1565 ( .A(n3132), .B(n3358), .C(n383), .Y(n2168) );
  AOI22X1 U1566 ( .A(n1132), .B(\data_in<8> ), .C(n1133), .D(\data_in<0> ), 
        .Y(n1131) );
  OAI21X1 U1567 ( .A(n3132), .B(n3357), .C(n382), .Y(n2169) );
  AOI22X1 U1568 ( .A(n1132), .B(\data_in<9> ), .C(n1133), .D(\data_in<1> ), 
        .Y(n1134) );
  OAI21X1 U1569 ( .A(n3132), .B(n3356), .C(n381), .Y(n2170) );
  AOI22X1 U1570 ( .A(n1132), .B(\data_in<10> ), .C(n1133), .D(\data_in<2> ), 
        .Y(n1135) );
  OAI21X1 U1571 ( .A(n3132), .B(n3355), .C(n380), .Y(n2171) );
  AOI22X1 U1572 ( .A(n1132), .B(\data_in<11> ), .C(n1133), .D(\data_in<3> ), 
        .Y(n1136) );
  OAI21X1 U1573 ( .A(n3132), .B(n3354), .C(n379), .Y(n2172) );
  AOI22X1 U1574 ( .A(n1132), .B(\data_in<12> ), .C(n1133), .D(\data_in<4> ), 
        .Y(n1137) );
  OAI21X1 U1575 ( .A(n3132), .B(n3353), .C(n378), .Y(n2173) );
  AOI22X1 U1576 ( .A(n1132), .B(\data_in<13> ), .C(n1133), .D(\data_in<5> ), 
        .Y(n1138) );
  OAI21X1 U1577 ( .A(n3132), .B(n3352), .C(n377), .Y(n2174) );
  AOI22X1 U1578 ( .A(n1132), .B(\data_in<14> ), .C(n1133), .D(\data_in<6> ), 
        .Y(n1139) );
  OAI21X1 U1579 ( .A(n3132), .B(n3351), .C(n376), .Y(n2175) );
  AOI22X1 U1580 ( .A(n1132), .B(\data_in<15> ), .C(n1133), .D(\data_in<7> ), 
        .Y(n1140) );
  AOI21X1 U1581 ( .A(n2487), .B(n2482), .C(n3177), .Y(n1130) );
  OAI21X1 U1582 ( .A(n3131), .B(n3350), .C(n375), .Y(n2176) );
  AOI22X1 U1583 ( .A(n1144), .B(\data_in<8> ), .C(n1145), .D(\data_in<0> ), 
        .Y(n1143) );
  OAI21X1 U1584 ( .A(n3131), .B(n3349), .C(n374), .Y(n2177) );
  AOI22X1 U1585 ( .A(n1144), .B(\data_in<9> ), .C(n1145), .D(\data_in<1> ), 
        .Y(n1146) );
  OAI21X1 U1586 ( .A(n3131), .B(n3348), .C(n373), .Y(n2178) );
  AOI22X1 U1587 ( .A(n1144), .B(\data_in<10> ), .C(n1145), .D(\data_in<2> ), 
        .Y(n1147) );
  OAI21X1 U1588 ( .A(n3131), .B(n3347), .C(n372), .Y(n2179) );
  AOI22X1 U1589 ( .A(n1144), .B(\data_in<11> ), .C(n1145), .D(\data_in<3> ), 
        .Y(n1148) );
  OAI21X1 U1590 ( .A(n3131), .B(n3346), .C(n371), .Y(n2180) );
  AOI22X1 U1591 ( .A(n1144), .B(\data_in<12> ), .C(n1145), .D(\data_in<4> ), 
        .Y(n1149) );
  OAI21X1 U1592 ( .A(n3131), .B(n3345), .C(n370), .Y(n2181) );
  AOI22X1 U1593 ( .A(n1144), .B(\data_in<13> ), .C(n1145), .D(\data_in<5> ), 
        .Y(n1150) );
  OAI21X1 U1594 ( .A(n3131), .B(n3344), .C(n369), .Y(n2182) );
  AOI22X1 U1595 ( .A(n1144), .B(\data_in<14> ), .C(n1145), .D(\data_in<6> ), 
        .Y(n1151) );
  OAI21X1 U1596 ( .A(n3131), .B(n3343), .C(n368), .Y(n2183) );
  AOI22X1 U1597 ( .A(n1144), .B(\data_in<15> ), .C(n1145), .D(\data_in<7> ), 
        .Y(n1152) );
  AOI21X1 U1598 ( .A(n2482), .B(n2483), .C(n3177), .Y(n1142) );
  OAI21X1 U1599 ( .A(n3130), .B(n3342), .C(n367), .Y(n2184) );
  AOI22X1 U1600 ( .A(n1156), .B(\data_in<8> ), .C(n1157), .D(\data_in<0> ), 
        .Y(n1155) );
  OAI21X1 U1601 ( .A(n3130), .B(n3341), .C(n366), .Y(n2185) );
  AOI22X1 U1602 ( .A(n1156), .B(\data_in<9> ), .C(n1157), .D(\data_in<1> ), 
        .Y(n1158) );
  OAI21X1 U1603 ( .A(n3130), .B(n3340), .C(n365), .Y(n2186) );
  AOI22X1 U1604 ( .A(n1156), .B(\data_in<10> ), .C(n1157), .D(\data_in<2> ), 
        .Y(n1159) );
  OAI21X1 U1605 ( .A(n3130), .B(n3339), .C(n364), .Y(n2187) );
  AOI22X1 U1606 ( .A(n1156), .B(\data_in<11> ), .C(n1157), .D(\data_in<3> ), 
        .Y(n1160) );
  OAI21X1 U1607 ( .A(n3130), .B(n3338), .C(n363), .Y(n2188) );
  AOI22X1 U1608 ( .A(n1156), .B(\data_in<12> ), .C(n1157), .D(\data_in<4> ), 
        .Y(n1161) );
  OAI21X1 U1609 ( .A(n3130), .B(n3337), .C(n362), .Y(n2189) );
  AOI22X1 U1610 ( .A(n1156), .B(\data_in<13> ), .C(n1157), .D(\data_in<5> ), 
        .Y(n1162) );
  OAI21X1 U1611 ( .A(n3130), .B(n3336), .C(n361), .Y(n2190) );
  AOI22X1 U1612 ( .A(n1156), .B(\data_in<14> ), .C(n1157), .D(\data_in<6> ), 
        .Y(n1163) );
  OAI21X1 U1613 ( .A(n3130), .B(n3335), .C(n360), .Y(n2191) );
  AOI22X1 U1614 ( .A(n1156), .B(\data_in<15> ), .C(n1157), .D(\data_in<7> ), 
        .Y(n1164) );
  AOI21X1 U1615 ( .A(n2483), .B(n2478), .C(n3177), .Y(n1154) );
  OAI21X1 U1616 ( .A(n3129), .B(n3334), .C(n359), .Y(n2192) );
  AOI22X1 U1617 ( .A(n1168), .B(\data_in<8> ), .C(n1169), .D(\data_in<0> ), 
        .Y(n1167) );
  OAI21X1 U1618 ( .A(n3129), .B(n3333), .C(n358), .Y(n2193) );
  AOI22X1 U1619 ( .A(n1168), .B(\data_in<9> ), .C(n1169), .D(\data_in<1> ), 
        .Y(n1170) );
  OAI21X1 U1620 ( .A(n3129), .B(n3332), .C(n357), .Y(n2194) );
  AOI22X1 U1621 ( .A(n1168), .B(\data_in<10> ), .C(n1169), .D(\data_in<2> ), 
        .Y(n1171) );
  OAI21X1 U1622 ( .A(n3129), .B(n3331), .C(n356), .Y(n2195) );
  AOI22X1 U1623 ( .A(n1168), .B(\data_in<11> ), .C(n1169), .D(\data_in<3> ), 
        .Y(n1172) );
  OAI21X1 U1624 ( .A(n3129), .B(n3330), .C(n355), .Y(n2196) );
  AOI22X1 U1625 ( .A(n1168), .B(\data_in<12> ), .C(n1169), .D(\data_in<4> ), 
        .Y(n1173) );
  OAI21X1 U1626 ( .A(n3129), .B(n3329), .C(n354), .Y(n2197) );
  AOI22X1 U1627 ( .A(n1168), .B(\data_in<13> ), .C(n1169), .D(\data_in<5> ), 
        .Y(n1174) );
  OAI21X1 U1628 ( .A(n3129), .B(n3328), .C(n353), .Y(n2198) );
  AOI22X1 U1629 ( .A(n1168), .B(\data_in<14> ), .C(n1169), .D(\data_in<6> ), 
        .Y(n1175) );
  OAI21X1 U1630 ( .A(n3129), .B(n3327), .C(n352), .Y(n2199) );
  AOI22X1 U1631 ( .A(n1168), .B(\data_in<15> ), .C(n1169), .D(\data_in<7> ), 
        .Y(n1176) );
  AOI21X1 U1632 ( .A(n2478), .B(n2479), .C(n3177), .Y(n1166) );
  OAI21X1 U1633 ( .A(n3128), .B(n3326), .C(n351), .Y(n2200) );
  AOI22X1 U1634 ( .A(n1180), .B(\data_in<8> ), .C(n1181), .D(\data_in<0> ), 
        .Y(n1179) );
  OAI21X1 U1635 ( .A(n3128), .B(n3325), .C(n350), .Y(n2201) );
  AOI22X1 U1636 ( .A(n1180), .B(\data_in<9> ), .C(n1181), .D(\data_in<1> ), 
        .Y(n1182) );
  OAI21X1 U1637 ( .A(n3128), .B(n3324), .C(n349), .Y(n2202) );
  AOI22X1 U1638 ( .A(n1180), .B(\data_in<10> ), .C(n1181), .D(\data_in<2> ), 
        .Y(n1183) );
  OAI21X1 U1639 ( .A(n3128), .B(n3323), .C(n348), .Y(n2203) );
  AOI22X1 U1640 ( .A(n1180), .B(\data_in<11> ), .C(n1181), .D(\data_in<3> ), 
        .Y(n1184) );
  OAI21X1 U1641 ( .A(n3128), .B(n3322), .C(n347), .Y(n2204) );
  AOI22X1 U1642 ( .A(n1180), .B(\data_in<12> ), .C(n1181), .D(\data_in<4> ), 
        .Y(n1185) );
  OAI21X1 U1643 ( .A(n3128), .B(n3321), .C(n346), .Y(n2205) );
  AOI22X1 U1644 ( .A(n1180), .B(\data_in<13> ), .C(n1181), .D(\data_in<5> ), 
        .Y(n1186) );
  OAI21X1 U1645 ( .A(n3128), .B(n3320), .C(n345), .Y(n2206) );
  AOI22X1 U1646 ( .A(n1180), .B(\data_in<14> ), .C(n1181), .D(\data_in<6> ), 
        .Y(n1187) );
  OAI21X1 U1647 ( .A(n3128), .B(n3319), .C(n344), .Y(n2207) );
  AOI22X1 U1648 ( .A(n1180), .B(\data_in<15> ), .C(n1181), .D(\data_in<7> ), 
        .Y(n1188) );
  AOI21X1 U1649 ( .A(n2479), .B(n2506), .C(n3177), .Y(n1178) );
  OAI21X1 U1650 ( .A(n3127), .B(n3318), .C(n343), .Y(n2208) );
  AOI22X1 U1651 ( .A(n1192), .B(\data_in<8> ), .C(n1193), .D(\data_in<0> ), 
        .Y(n1191) );
  OAI21X1 U1652 ( .A(n3127), .B(n3317), .C(n342), .Y(n2209) );
  AOI22X1 U1653 ( .A(n1192), .B(\data_in<9> ), .C(n1193), .D(\data_in<1> ), 
        .Y(n1194) );
  OAI21X1 U1654 ( .A(n3127), .B(n3316), .C(n341), .Y(n2210) );
  AOI22X1 U1655 ( .A(n1192), .B(\data_in<10> ), .C(n1193), .D(\data_in<2> ), 
        .Y(n1195) );
  OAI21X1 U1656 ( .A(n3127), .B(n3315), .C(n340), .Y(n2211) );
  AOI22X1 U1657 ( .A(n1192), .B(\data_in<11> ), .C(n1193), .D(\data_in<3> ), 
        .Y(n1196) );
  OAI21X1 U1658 ( .A(n3127), .B(n3314), .C(n339), .Y(n2212) );
  AOI22X1 U1659 ( .A(n1192), .B(\data_in<12> ), .C(n1193), .D(\data_in<4> ), 
        .Y(n1197) );
  OAI21X1 U1660 ( .A(n3127), .B(n3313), .C(n338), .Y(n2213) );
  AOI22X1 U1661 ( .A(n1192), .B(\data_in<13> ), .C(n1193), .D(\data_in<5> ), 
        .Y(n1198) );
  OAI21X1 U1662 ( .A(n3127), .B(n3312), .C(n337), .Y(n2214) );
  AOI22X1 U1663 ( .A(n1192), .B(\data_in<14> ), .C(n1193), .D(\data_in<6> ), 
        .Y(n1199) );
  OAI21X1 U1664 ( .A(n3127), .B(n3311), .C(n336), .Y(n2215) );
  AOI22X1 U1665 ( .A(n1192), .B(\data_in<15> ), .C(n1193), .D(\data_in<7> ), 
        .Y(n1200) );
  AOI21X1 U1666 ( .A(n2506), .B(n2508), .C(n3176), .Y(n1190) );
  OAI21X1 U1667 ( .A(n3126), .B(n3310), .C(n335), .Y(n2216) );
  AOI22X1 U1668 ( .A(n1204), .B(\data_in<8> ), .C(n1205), .D(\data_in<0> ), 
        .Y(n1203) );
  OAI21X1 U1669 ( .A(n3126), .B(n3309), .C(n334), .Y(n2217) );
  AOI22X1 U1670 ( .A(n1204), .B(\data_in<9> ), .C(n1205), .D(\data_in<1> ), 
        .Y(n1206) );
  OAI21X1 U1671 ( .A(n3126), .B(n3308), .C(n333), .Y(n2218) );
  AOI22X1 U1672 ( .A(n1204), .B(\data_in<10> ), .C(n1205), .D(\data_in<2> ), 
        .Y(n1207) );
  OAI21X1 U1673 ( .A(n3126), .B(n3307), .C(n332), .Y(n2219) );
  AOI22X1 U1674 ( .A(n1204), .B(\data_in<11> ), .C(n1205), .D(\data_in<3> ), 
        .Y(n1208) );
  OAI21X1 U1675 ( .A(n3126), .B(n3306), .C(n331), .Y(n2220) );
  AOI22X1 U1676 ( .A(n1204), .B(\data_in<12> ), .C(n1205), .D(\data_in<4> ), 
        .Y(n1209) );
  OAI21X1 U1677 ( .A(n3126), .B(n3305), .C(n330), .Y(n2221) );
  AOI22X1 U1678 ( .A(n1204), .B(\data_in<13> ), .C(n1205), .D(\data_in<5> ), 
        .Y(n1210) );
  OAI21X1 U1679 ( .A(n3126), .B(n3304), .C(n329), .Y(n2222) );
  AOI22X1 U1680 ( .A(n1204), .B(\data_in<14> ), .C(n1205), .D(\data_in<6> ), 
        .Y(n1211) );
  OAI21X1 U1681 ( .A(n3126), .B(n3303), .C(n328), .Y(n2223) );
  AOI22X1 U1682 ( .A(n1204), .B(\data_in<15> ), .C(n1205), .D(\data_in<7> ), 
        .Y(n1212) );
  AOI21X1 U1683 ( .A(n2508), .B(n2502), .C(n3176), .Y(n1202) );
  OAI21X1 U1684 ( .A(n3125), .B(n3302), .C(n327), .Y(n2224) );
  AOI22X1 U1685 ( .A(n1216), .B(\data_in<8> ), .C(n1217), .D(\data_in<0> ), 
        .Y(n1215) );
  OAI21X1 U1686 ( .A(n3125), .B(n3301), .C(n326), .Y(n2225) );
  AOI22X1 U1687 ( .A(n1216), .B(\data_in<9> ), .C(n1217), .D(\data_in<1> ), 
        .Y(n1218) );
  OAI21X1 U1688 ( .A(n3125), .B(n3300), .C(n325), .Y(n2226) );
  AOI22X1 U1689 ( .A(n1216), .B(\data_in<10> ), .C(n1217), .D(\data_in<2> ), 
        .Y(n1219) );
  OAI21X1 U1690 ( .A(n3125), .B(n3299), .C(n324), .Y(n2227) );
  AOI22X1 U1691 ( .A(n1216), .B(\data_in<11> ), .C(n1217), .D(\data_in<3> ), 
        .Y(n1220) );
  OAI21X1 U1692 ( .A(n3125), .B(n3298), .C(n323), .Y(n2228) );
  AOI22X1 U1693 ( .A(n1216), .B(\data_in<12> ), .C(n1217), .D(\data_in<4> ), 
        .Y(n1221) );
  OAI21X1 U1694 ( .A(n3125), .B(n3297), .C(n322), .Y(n2229) );
  AOI22X1 U1695 ( .A(n1216), .B(\data_in<13> ), .C(n1217), .D(\data_in<5> ), 
        .Y(n1222) );
  OAI21X1 U1696 ( .A(n3125), .B(n3296), .C(n321), .Y(n2230) );
  AOI22X1 U1697 ( .A(n1216), .B(\data_in<14> ), .C(n1217), .D(\data_in<6> ), 
        .Y(n1223) );
  OAI21X1 U1698 ( .A(n3125), .B(n3295), .C(n320), .Y(n2231) );
  AOI22X1 U1699 ( .A(n1216), .B(\data_in<15> ), .C(n1217), .D(\data_in<7> ), 
        .Y(n1224) );
  AOI21X1 U1700 ( .A(n2502), .B(n2504), .C(n3176), .Y(n1214) );
  OAI21X1 U1701 ( .A(n3124), .B(n3294), .C(n319), .Y(n2232) );
  AOI22X1 U1702 ( .A(n1228), .B(\data_in<8> ), .C(n1229), .D(\data_in<0> ), 
        .Y(n1227) );
  OAI21X1 U1703 ( .A(n3124), .B(n3293), .C(n318), .Y(n2233) );
  AOI22X1 U1704 ( .A(n1228), .B(\data_in<9> ), .C(n1229), .D(\data_in<1> ), 
        .Y(n1230) );
  OAI21X1 U1705 ( .A(n3124), .B(n3292), .C(n317), .Y(n2234) );
  AOI22X1 U1706 ( .A(n1228), .B(\data_in<10> ), .C(n1229), .D(\data_in<2> ), 
        .Y(n1231) );
  OAI21X1 U1707 ( .A(n3124), .B(n3291), .C(n316), .Y(n2235) );
  AOI22X1 U1708 ( .A(n1228), .B(\data_in<11> ), .C(n1229), .D(\data_in<3> ), 
        .Y(n1232) );
  OAI21X1 U1709 ( .A(n3124), .B(n3290), .C(n315), .Y(n2236) );
  AOI22X1 U1710 ( .A(n1228), .B(\data_in<12> ), .C(n1229), .D(\data_in<4> ), 
        .Y(n1233) );
  OAI21X1 U1711 ( .A(n3124), .B(n3289), .C(n314), .Y(n2237) );
  AOI22X1 U1712 ( .A(n1228), .B(\data_in<13> ), .C(n1229), .D(\data_in<5> ), 
        .Y(n1234) );
  OAI21X1 U1713 ( .A(n3124), .B(n3288), .C(n313), .Y(n2238) );
  AOI22X1 U1714 ( .A(n1228), .B(\data_in<14> ), .C(n1229), .D(\data_in<6> ), 
        .Y(n1235) );
  OAI21X1 U1715 ( .A(n3124), .B(n3287), .C(n312), .Y(n2239) );
  AOI22X1 U1716 ( .A(n1228), .B(\data_in<15> ), .C(n1229), .D(\data_in<7> ), 
        .Y(n1236) );
  AOI21X1 U1717 ( .A(n2504), .B(n2498), .C(n3176), .Y(n1226) );
  OAI21X1 U1718 ( .A(n3123), .B(n3286), .C(n311), .Y(n2240) );
  AOI22X1 U1719 ( .A(n1240), .B(\data_in<8> ), .C(n1241), .D(\data_in<0> ), 
        .Y(n1239) );
  OAI21X1 U1720 ( .A(n3123), .B(n3285), .C(n310), .Y(n2241) );
  AOI22X1 U1721 ( .A(n1240), .B(\data_in<9> ), .C(n1241), .D(\data_in<1> ), 
        .Y(n1242) );
  OAI21X1 U1722 ( .A(n3123), .B(n3284), .C(n309), .Y(n2242) );
  AOI22X1 U1723 ( .A(n1240), .B(\data_in<10> ), .C(n1241), .D(\data_in<2> ), 
        .Y(n1243) );
  OAI21X1 U1724 ( .A(n3123), .B(n3283), .C(n308), .Y(n2243) );
  AOI22X1 U1725 ( .A(n1240), .B(\data_in<11> ), .C(n1241), .D(\data_in<3> ), 
        .Y(n1244) );
  OAI21X1 U1726 ( .A(n3123), .B(n3282), .C(n307), .Y(n2244) );
  AOI22X1 U1727 ( .A(n1240), .B(\data_in<12> ), .C(n1241), .D(\data_in<4> ), 
        .Y(n1245) );
  OAI21X1 U1728 ( .A(n3123), .B(n3281), .C(n306), .Y(n2245) );
  AOI22X1 U1729 ( .A(n1240), .B(\data_in<13> ), .C(n1241), .D(\data_in<5> ), 
        .Y(n1246) );
  OAI21X1 U1730 ( .A(n3123), .B(n3280), .C(n305), .Y(n2246) );
  AOI22X1 U1731 ( .A(n1240), .B(\data_in<14> ), .C(n1241), .D(\data_in<6> ), 
        .Y(n1247) );
  OAI21X1 U1732 ( .A(n3123), .B(n3279), .C(n304), .Y(n2247) );
  AOI22X1 U1733 ( .A(n1240), .B(\data_in<15> ), .C(n1241), .D(\data_in<7> ), 
        .Y(n1248) );
  AOI21X1 U1734 ( .A(n2498), .B(n2500), .C(n3176), .Y(n1238) );
  OAI21X1 U1735 ( .A(n3122), .B(n3278), .C(n303), .Y(n2248) );
  AOI22X1 U1736 ( .A(n1252), .B(\data_in<8> ), .C(n1253), .D(\data_in<0> ), 
        .Y(n1251) );
  OAI21X1 U1737 ( .A(n3122), .B(n3277), .C(n302), .Y(n2249) );
  AOI22X1 U1738 ( .A(n1252), .B(\data_in<9> ), .C(n1253), .D(\data_in<1> ), 
        .Y(n1254) );
  OAI21X1 U1739 ( .A(n3122), .B(n3276), .C(n301), .Y(n2250) );
  AOI22X1 U1740 ( .A(n1252), .B(\data_in<10> ), .C(n1253), .D(\data_in<2> ), 
        .Y(n1255) );
  OAI21X1 U1741 ( .A(n3122), .B(n3275), .C(n300), .Y(n2251) );
  AOI22X1 U1742 ( .A(n1252), .B(\data_in<11> ), .C(n1253), .D(\data_in<3> ), 
        .Y(n1256) );
  OAI21X1 U1743 ( .A(n3122), .B(n3274), .C(n299), .Y(n2252) );
  AOI22X1 U1744 ( .A(n1252), .B(\data_in<12> ), .C(n1253), .D(\data_in<4> ), 
        .Y(n1257) );
  OAI21X1 U1745 ( .A(n3122), .B(n3273), .C(n298), .Y(n2253) );
  AOI22X1 U1746 ( .A(n1252), .B(\data_in<13> ), .C(n1253), .D(\data_in<5> ), 
        .Y(n1258) );
  OAI21X1 U1747 ( .A(n3122), .B(n3272), .C(n297), .Y(n2254) );
  AOI22X1 U1748 ( .A(n1252), .B(\data_in<14> ), .C(n1253), .D(\data_in<6> ), 
        .Y(n1259) );
  OAI21X1 U1749 ( .A(n3122), .B(n3271), .C(n296), .Y(n2255) );
  AOI22X1 U1750 ( .A(n1252), .B(\data_in<15> ), .C(n1253), .D(\data_in<7> ), 
        .Y(n1260) );
  AOI21X1 U1751 ( .A(n2500), .B(n2494), .C(n3176), .Y(n1250) );
  OAI21X1 U1752 ( .A(n3121), .B(n3270), .C(n295), .Y(n2256) );
  AOI22X1 U1753 ( .A(n1264), .B(\data_in<8> ), .C(n1265), .D(\data_in<0> ), 
        .Y(n1263) );
  OAI21X1 U1754 ( .A(n3121), .B(n3269), .C(n294), .Y(n2257) );
  AOI22X1 U1755 ( .A(n1264), .B(\data_in<9> ), .C(n1265), .D(\data_in<1> ), 
        .Y(n1266) );
  OAI21X1 U1756 ( .A(n3121), .B(n3268), .C(n293), .Y(n2258) );
  AOI22X1 U1757 ( .A(n1264), .B(\data_in<10> ), .C(n1265), .D(\data_in<2> ), 
        .Y(n1267) );
  OAI21X1 U1758 ( .A(n3121), .B(n3267), .C(n292), .Y(n2259) );
  AOI22X1 U1759 ( .A(n1264), .B(\data_in<11> ), .C(n1265), .D(\data_in<3> ), 
        .Y(n1268) );
  OAI21X1 U1760 ( .A(n3121), .B(n3266), .C(n291), .Y(n2260) );
  AOI22X1 U1761 ( .A(n1264), .B(\data_in<12> ), .C(n1265), .D(\data_in<4> ), 
        .Y(n1269) );
  OAI21X1 U1762 ( .A(n3121), .B(n3265), .C(n290), .Y(n2261) );
  AOI22X1 U1763 ( .A(n1264), .B(\data_in<13> ), .C(n1265), .D(\data_in<5> ), 
        .Y(n1270) );
  OAI21X1 U1764 ( .A(n3121), .B(n3264), .C(n289), .Y(n2262) );
  AOI22X1 U1765 ( .A(n1264), .B(\data_in<14> ), .C(n1265), .D(\data_in<6> ), 
        .Y(n1271) );
  OAI21X1 U1766 ( .A(n3121), .B(n3263), .C(n288), .Y(n2263) );
  AOI22X1 U1767 ( .A(n1264), .B(\data_in<15> ), .C(n1265), .D(\data_in<7> ), 
        .Y(n1272) );
  AOI21X1 U1768 ( .A(n2494), .B(n2496), .C(n3176), .Y(n1262) );
  OAI21X1 U1769 ( .A(n3120), .B(n3262), .C(n287), .Y(n2264) );
  AOI22X1 U1770 ( .A(n1276), .B(\data_in<8> ), .C(n1277), .D(\data_in<0> ), 
        .Y(n1275) );
  OAI21X1 U1771 ( .A(n3120), .B(n3261), .C(n286), .Y(n2265) );
  AOI22X1 U1772 ( .A(n1276), .B(\data_in<9> ), .C(n1277), .D(\data_in<1> ), 
        .Y(n1278) );
  OAI21X1 U1773 ( .A(n3120), .B(n3260), .C(n285), .Y(n2266) );
  AOI22X1 U1774 ( .A(n1276), .B(\data_in<10> ), .C(n1277), .D(\data_in<2> ), 
        .Y(n1279) );
  OAI21X1 U1775 ( .A(n3120), .B(n3259), .C(n284), .Y(n2267) );
  AOI22X1 U1776 ( .A(n1276), .B(\data_in<11> ), .C(n1277), .D(\data_in<3> ), 
        .Y(n1280) );
  OAI21X1 U1777 ( .A(n3120), .B(n3258), .C(n283), .Y(n2268) );
  AOI22X1 U1778 ( .A(n1276), .B(\data_in<12> ), .C(n1277), .D(\data_in<4> ), 
        .Y(n1281) );
  OAI21X1 U1779 ( .A(n3120), .B(n3257), .C(n282), .Y(n2269) );
  AOI22X1 U1780 ( .A(n1276), .B(\data_in<13> ), .C(n1277), .D(\data_in<5> ), 
        .Y(n1282) );
  OAI21X1 U1781 ( .A(n3120), .B(n3256), .C(n281), .Y(n2270) );
  AOI22X1 U1782 ( .A(n1276), .B(\data_in<14> ), .C(n1277), .D(\data_in<6> ), 
        .Y(n1283) );
  OAI21X1 U1783 ( .A(n3120), .B(n3255), .C(n280), .Y(n2271) );
  AOI22X1 U1784 ( .A(n1276), .B(\data_in<15> ), .C(n1277), .D(\data_in<7> ), 
        .Y(n1284) );
  AOI21X1 U1785 ( .A(n2496), .B(n2516), .C(n3176), .Y(n1274) );
  OAI21X1 U1786 ( .A(n3119), .B(n3254), .C(n279), .Y(n2272) );
  AOI22X1 U1787 ( .A(n1288), .B(\data_in<8> ), .C(n1289), .D(\data_in<0> ), 
        .Y(n1287) );
  OAI21X1 U1788 ( .A(n3119), .B(n3253), .C(n278), .Y(n2273) );
  AOI22X1 U1789 ( .A(n1288), .B(\data_in<9> ), .C(n1289), .D(\data_in<1> ), 
        .Y(n1290) );
  OAI21X1 U1790 ( .A(n3119), .B(n3252), .C(n277), .Y(n2274) );
  AOI22X1 U1791 ( .A(n1288), .B(\data_in<10> ), .C(n1289), .D(\data_in<2> ), 
        .Y(n1291) );
  OAI21X1 U1792 ( .A(n3119), .B(n3251), .C(n276), .Y(n2275) );
  AOI22X1 U1793 ( .A(n1288), .B(\data_in<11> ), .C(n1289), .D(\data_in<3> ), 
        .Y(n1292) );
  OAI21X1 U1794 ( .A(n3119), .B(n3250), .C(n275), .Y(n2276) );
  AOI22X1 U1795 ( .A(n1288), .B(\data_in<12> ), .C(n1289), .D(\data_in<4> ), 
        .Y(n1293) );
  OAI21X1 U1796 ( .A(n3119), .B(n3249), .C(n274), .Y(n2277) );
  AOI22X1 U1797 ( .A(n1288), .B(\data_in<13> ), .C(n1289), .D(\data_in<5> ), 
        .Y(n1294) );
  OAI21X1 U1798 ( .A(n3119), .B(n3248), .C(n273), .Y(n2278) );
  AOI22X1 U1799 ( .A(n1288), .B(\data_in<14> ), .C(n1289), .D(\data_in<6> ), 
        .Y(n1295) );
  OAI21X1 U1800 ( .A(n3119), .B(n3247), .C(n272), .Y(n2279) );
  AOI22X1 U1801 ( .A(n1288), .B(\data_in<15> ), .C(n1289), .D(\data_in<7> ), 
        .Y(n1296) );
  AOI21X1 U1802 ( .A(n2516), .B(n2518), .C(n3176), .Y(n1286) );
  OAI21X1 U1803 ( .A(n3118), .B(n3246), .C(n271), .Y(n2280) );
  AOI22X1 U1804 ( .A(n1300), .B(\data_in<8> ), .C(n1301), .D(\data_in<0> ), 
        .Y(n1299) );
  OAI21X1 U1805 ( .A(n3118), .B(n3245), .C(n270), .Y(n2281) );
  AOI22X1 U1806 ( .A(n1300), .B(\data_in<9> ), .C(n1301), .D(\data_in<1> ), 
        .Y(n1302) );
  OAI21X1 U1807 ( .A(n3118), .B(n3244), .C(n269), .Y(n2282) );
  AOI22X1 U1808 ( .A(n1300), .B(\data_in<10> ), .C(n1301), .D(\data_in<2> ), 
        .Y(n1303) );
  OAI21X1 U1809 ( .A(n3118), .B(n3243), .C(n268), .Y(n2283) );
  AOI22X1 U1810 ( .A(n1300), .B(\data_in<11> ), .C(n1301), .D(\data_in<3> ), 
        .Y(n1304) );
  OAI21X1 U1811 ( .A(n3118), .B(n3242), .C(n267), .Y(n2284) );
  AOI22X1 U1812 ( .A(n1300), .B(\data_in<12> ), .C(n1301), .D(\data_in<4> ), 
        .Y(n1305) );
  OAI21X1 U1813 ( .A(n3118), .B(n3241), .C(n266), .Y(n2285) );
  AOI22X1 U1814 ( .A(n1300), .B(\data_in<13> ), .C(n1301), .D(\data_in<5> ), 
        .Y(n1306) );
  OAI21X1 U1815 ( .A(n3118), .B(n3240), .C(n265), .Y(n2286) );
  AOI22X1 U1816 ( .A(n1300), .B(\data_in<14> ), .C(n1301), .D(\data_in<6> ), 
        .Y(n1307) );
  OAI21X1 U1817 ( .A(n3118), .B(n3239), .C(n264), .Y(n2287) );
  AOI22X1 U1818 ( .A(n1300), .B(\data_in<15> ), .C(n1301), .D(\data_in<7> ), 
        .Y(n1308) );
  AOI21X1 U1819 ( .A(n2518), .B(n2512), .C(n3176), .Y(n1298) );
  OAI21X1 U1820 ( .A(n3117), .B(n3238), .C(n263), .Y(n2288) );
  AOI22X1 U1821 ( .A(n1312), .B(\data_in<8> ), .C(n1313), .D(\data_in<0> ), 
        .Y(n1311) );
  OAI21X1 U1822 ( .A(n3117), .B(n3237), .C(n262), .Y(n2289) );
  AOI22X1 U1823 ( .A(n1312), .B(\data_in<9> ), .C(n1313), .D(\data_in<1> ), 
        .Y(n1314) );
  OAI21X1 U1824 ( .A(n3117), .B(n3236), .C(n261), .Y(n2290) );
  AOI22X1 U1825 ( .A(n1312), .B(\data_in<10> ), .C(n1313), .D(\data_in<2> ), 
        .Y(n1315) );
  OAI21X1 U1826 ( .A(n3117), .B(n3235), .C(n260), .Y(n2291) );
  AOI22X1 U1827 ( .A(n1312), .B(\data_in<11> ), .C(n1313), .D(\data_in<3> ), 
        .Y(n1316) );
  OAI21X1 U1828 ( .A(n3117), .B(n3234), .C(n259), .Y(n2292) );
  AOI22X1 U1829 ( .A(n1312), .B(\data_in<12> ), .C(n1313), .D(\data_in<4> ), 
        .Y(n1317) );
  OAI21X1 U1830 ( .A(n3117), .B(n3233), .C(n258), .Y(n2293) );
  AOI22X1 U1831 ( .A(n1312), .B(\data_in<13> ), .C(n1313), .D(\data_in<5> ), 
        .Y(n1318) );
  OAI21X1 U1832 ( .A(n3117), .B(n3232), .C(n257), .Y(n2294) );
  AOI22X1 U1833 ( .A(n1312), .B(\data_in<14> ), .C(n1313), .D(\data_in<6> ), 
        .Y(n1319) );
  OAI21X1 U1834 ( .A(n3117), .B(n3231), .C(n256), .Y(n2295) );
  AOI22X1 U1835 ( .A(n1312), .B(\data_in<15> ), .C(n1313), .D(\data_in<7> ), 
        .Y(n1320) );
  AOI21X1 U1836 ( .A(n2512), .B(n2514), .C(n3176), .Y(n1310) );
  OAI21X1 U1837 ( .A(n3116), .B(n3230), .C(n255), .Y(n2296) );
  AOI22X1 U1838 ( .A(n1324), .B(\data_in<8> ), .C(n1325), .D(\data_in<0> ), 
        .Y(n1323) );
  OAI21X1 U1839 ( .A(n3116), .B(n3229), .C(n254), .Y(n2297) );
  AOI22X1 U1840 ( .A(n1324), .B(\data_in<9> ), .C(n1325), .D(\data_in<1> ), 
        .Y(n1326) );
  OAI21X1 U1841 ( .A(n3116), .B(n3228), .C(n253), .Y(n2298) );
  AOI22X1 U1842 ( .A(n1324), .B(\data_in<10> ), .C(n1325), .D(\data_in<2> ), 
        .Y(n1327) );
  OAI21X1 U1843 ( .A(n3116), .B(n3227), .C(n252), .Y(n2299) );
  AOI22X1 U1844 ( .A(n1324), .B(\data_in<11> ), .C(n1325), .D(\data_in<3> ), 
        .Y(n1328) );
  OAI21X1 U1845 ( .A(n3116), .B(n3226), .C(n251), .Y(n2300) );
  AOI22X1 U1846 ( .A(n1324), .B(\data_in<12> ), .C(n1325), .D(\data_in<4> ), 
        .Y(n1329) );
  OAI21X1 U1847 ( .A(n3116), .B(n3225), .C(n250), .Y(n2301) );
  AOI22X1 U1848 ( .A(n1324), .B(\data_in<13> ), .C(n1325), .D(\data_in<5> ), 
        .Y(n1330) );
  OAI21X1 U1849 ( .A(n3116), .B(n3224), .C(n249), .Y(n2302) );
  AOI22X1 U1850 ( .A(n1324), .B(\data_in<14> ), .C(n1325), .D(\data_in<6> ), 
        .Y(n1331) );
  OAI21X1 U1851 ( .A(n3116), .B(n3223), .C(n248), .Y(n2303) );
  AOI22X1 U1852 ( .A(n1324), .B(\data_in<15> ), .C(n1325), .D(\data_in<7> ), 
        .Y(n1332) );
  AOI21X1 U1853 ( .A(n2514), .B(n2510), .C(n3176), .Y(n1322) );
  OAI21X1 U1854 ( .A(n3115), .B(n3222), .C(n247), .Y(n2304) );
  AOI22X1 U1855 ( .A(n1336), .B(\data_in<8> ), .C(n1337), .D(\data_in<0> ), 
        .Y(n1335) );
  OAI21X1 U1856 ( .A(n3115), .B(n3221), .C(n246), .Y(n2305) );
  AOI22X1 U1857 ( .A(n1336), .B(\data_in<9> ), .C(n1337), .D(\data_in<1> ), 
        .Y(n1338) );
  OAI21X1 U1858 ( .A(n3115), .B(n3220), .C(n245), .Y(n2306) );
  AOI22X1 U1859 ( .A(n1336), .B(\data_in<10> ), .C(n1337), .D(\data_in<2> ), 
        .Y(n1339) );
  OAI21X1 U1860 ( .A(n3115), .B(n3219), .C(n244), .Y(n2307) );
  AOI22X1 U1861 ( .A(n1336), .B(\data_in<11> ), .C(n1337), .D(\data_in<3> ), 
        .Y(n1340) );
  OAI21X1 U1862 ( .A(n3115), .B(n3218), .C(n243), .Y(n2308) );
  AOI22X1 U1863 ( .A(n1336), .B(\data_in<12> ), .C(n1337), .D(\data_in<4> ), 
        .Y(n1341) );
  OAI21X1 U1864 ( .A(n3115), .B(n3217), .C(n242), .Y(n2309) );
  AOI22X1 U1865 ( .A(n1336), .B(\data_in<13> ), .C(n1337), .D(\data_in<5> ), 
        .Y(n1342) );
  OAI21X1 U1866 ( .A(n3115), .B(n3216), .C(n241), .Y(n2310) );
  AOI22X1 U1867 ( .A(n1336), .B(\data_in<14> ), .C(n1337), .D(\data_in<6> ), 
        .Y(n1343) );
  OAI21X1 U1868 ( .A(n3115), .B(n3215), .C(n240), .Y(n2311) );
  AOI22X1 U1869 ( .A(n1336), .B(\data_in<15> ), .C(n1337), .D(\data_in<7> ), 
        .Y(n1344) );
  AOI21X1 U1870 ( .A(n2510), .B(n2582), .C(n3176), .Y(n1334) );
  OAI21X1 U1871 ( .A(n3114), .B(n3214), .C(n239), .Y(n2312) );
  AOI22X1 U1872 ( .A(n1348), .B(\data_in<8> ), .C(n1349), .D(\data_in<0> ), 
        .Y(n1347) );
  OAI21X1 U1873 ( .A(n3114), .B(n3213), .C(n238), .Y(n2313) );
  AOI22X1 U1874 ( .A(n1348), .B(\data_in<9> ), .C(n1349), .D(\data_in<1> ), 
        .Y(n1350) );
  OAI21X1 U1875 ( .A(n3114), .B(n3212), .C(n237), .Y(n2314) );
  AOI22X1 U1876 ( .A(n1348), .B(\data_in<10> ), .C(n1349), .D(\data_in<2> ), 
        .Y(n1351) );
  OAI21X1 U1877 ( .A(n3114), .B(n3211), .C(n236), .Y(n2315) );
  AOI22X1 U1878 ( .A(n1348), .B(\data_in<11> ), .C(n1349), .D(\data_in<3> ), 
        .Y(n1352) );
  OAI21X1 U1879 ( .A(n3114), .B(n3210), .C(n235), .Y(n2316) );
  AOI22X1 U1880 ( .A(n1348), .B(\data_in<12> ), .C(n1349), .D(\data_in<4> ), 
        .Y(n1353) );
  OAI21X1 U1881 ( .A(n3114), .B(n3209), .C(n234), .Y(n2317) );
  AOI22X1 U1882 ( .A(n1348), .B(\data_in<13> ), .C(n1349), .D(\data_in<5> ), 
        .Y(n1354) );
  OAI21X1 U1883 ( .A(n3114), .B(n3208), .C(n233), .Y(n2318) );
  AOI22X1 U1884 ( .A(n1348), .B(\data_in<14> ), .C(n1349), .D(\data_in<6> ), 
        .Y(n1355) );
  OAI21X1 U1885 ( .A(n3114), .B(n3207), .C(n232), .Y(n2319) );
  AOI22X1 U1886 ( .A(n1348), .B(\data_in<15> ), .C(n1349), .D(\data_in<7> ), 
        .Y(n1356) );
  OAI21X1 U1887 ( .A(n3176), .B(n2582), .C(n2458), .Y(n1346) );
  OAI21X1 U1888 ( .A(n3190), .B(n3206), .C(n2338), .Y(n2320) );
  OAI21X1 U1890 ( .A(n3190), .B(n3205), .C(n2336), .Y(n2321) );
  OAI21X1 U1892 ( .A(n3190), .B(n3204), .C(n2334), .Y(n2322) );
  OAI21X1 U1894 ( .A(n3190), .B(n3203), .C(n2332), .Y(n2323) );
  OAI21X1 U1896 ( .A(n3190), .B(n3202), .C(n2330), .Y(n2324) );
  OAI21X1 U1898 ( .A(n3190), .B(n3201), .C(n2328), .Y(n2325) );
  OAI21X1 U1900 ( .A(n3190), .B(n3200), .C(n1796), .Y(n2326) );
  OAI21X1 U1902 ( .A(n3190), .B(n3199), .C(n1794), .Y(n2327) );
  NAND3X1 U1905 ( .A(enable), .B(n3188), .C(wr), .Y(n625) );
  AOI21X1 U1906 ( .A(n1367), .B(n1368), .C(n2451), .Y(n3712) );
  NOR3X1 U1907 ( .A(n1370), .B(n180), .C(n188), .Y(n1368) );
  AOI22X1 U1909 ( .A(\mem<55><7> ), .B(n2577), .C(\mem<54><7> ), .D(n2580), 
        .Y(n1377) );
  AOI22X1 U1910 ( .A(\mem<53><7> ), .B(n2573), .C(\mem<52><7> ), .D(n2576), 
        .Y(n1376) );
  AOI22X1 U1911 ( .A(\mem<51><7> ), .B(n2569), .C(\mem<50><7> ), .D(n2572), 
        .Y(n1374) );
  AOI22X1 U1912 ( .A(\mem<49><7> ), .B(n2565), .C(\mem<48><7> ), .D(n2568), 
        .Y(n1373) );
  AOI22X1 U1914 ( .A(\mem<63><7> ), .B(n2459), .C(\mem<62><7> ), .D(n2564), 
        .Y(n1382) );
  AOI22X1 U1915 ( .A(\mem<61><7> ), .B(n2559), .C(\mem<60><7> ), .D(n2562), 
        .Y(n1381) );
  AOI22X1 U1916 ( .A(\mem<59><7> ), .B(n2555), .C(\mem<58><7> ), .D(n2558), 
        .Y(n1379) );
  AOI22X1 U1917 ( .A(\mem<57><7> ), .B(n2551), .C(\mem<56><7> ), .D(n2554), 
        .Y(n1378) );
  AOI22X1 U1919 ( .A(\mem<39><7> ), .B(n2547), .C(\mem<38><7> ), .D(n2550), 
        .Y(n1389) );
  AOI22X1 U1920 ( .A(\mem<37><7> ), .B(n2543), .C(\mem<36><7> ), .D(n2546), 
        .Y(n1388) );
  AOI22X1 U1921 ( .A(\mem<35><7> ), .B(n2539), .C(\mem<34><7> ), .D(n2542), 
        .Y(n1386) );
  AOI22X1 U1922 ( .A(\mem<33><7> ), .B(n2536), .C(\mem<32><7> ), .D(n2537), 
        .Y(n1385) );
  AOI22X1 U1924 ( .A(\mem<47><7> ), .B(n2531), .C(\mem<46><7> ), .D(n2534), 
        .Y(n1394) );
  AOI22X1 U1925 ( .A(\mem<45><7> ), .B(n2527), .C(\mem<44><7> ), .D(n2530), 
        .Y(n1393) );
  AOI22X1 U1926 ( .A(\mem<43><7> ), .B(n2523), .C(\mem<42><7> ), .D(n2526), 
        .Y(n1391) );
  AOI22X1 U1927 ( .A(\mem<41><7> ), .B(n2519), .C(\mem<40><7> ), .D(n2522), 
        .Y(n1390) );
  NOR3X1 U1928 ( .A(n1395), .B(n179), .C(n229), .Y(n1367) );
  AOI22X1 U1930 ( .A(\mem<7><7> ), .B(n2515), .C(\mem<6><7> ), .D(n2517), .Y(
        n1402) );
  AOI22X1 U1931 ( .A(\mem<5><7> ), .B(n2511), .C(\mem<4><7> ), .D(n2513), .Y(
        n1401) );
  AOI22X1 U1932 ( .A(\mem<3><7> ), .B(n2509), .C(\mem<2><7> ), .D(n2581), .Y(
        n1399) );
  AOI22X1 U1933 ( .A(\mem<1><7> ), .B(n2455), .C(n1403), .D(\mem<0><7> ), .Y(
        n1398) );
  AOI22X1 U1935 ( .A(\mem<15><7> ), .B(n2505), .C(\mem<14><7> ), .D(n2507), 
        .Y(n1408) );
  AOI22X1 U1936 ( .A(\mem<13><7> ), .B(n2501), .C(\mem<12><7> ), .D(n2503), 
        .Y(n1407) );
  AOI22X1 U1937 ( .A(\mem<11><7> ), .B(n2497), .C(\mem<10><7> ), .D(n2499), 
        .Y(n1405) );
  AOI22X1 U1938 ( .A(\mem<9><7> ), .B(n2493), .C(\mem<8><7> ), .D(n2495), .Y(
        n1404) );
  AOI22X1 U1940 ( .A(\mem<23><7> ), .B(n2489), .C(\mem<22><7> ), .D(n2492), 
        .Y(n1415) );
  AOI22X1 U1941 ( .A(\mem<21><7> ), .B(n2485), .C(\mem<20><7> ), .D(n2488), 
        .Y(n1414) );
  AOI22X1 U1942 ( .A(\mem<19><7> ), .B(n2481), .C(\mem<18><7> ), .D(n2484), 
        .Y(n1412) );
  AOI22X1 U1943 ( .A(\mem<17><7> ), .B(n2477), .C(\mem<16><7> ), .D(n2480), 
        .Y(n1411) );
  AOI22X1 U1945 ( .A(\mem<31><7> ), .B(n2473), .C(\mem<30><7> ), .D(n2476), 
        .Y(n1420) );
  AOI22X1 U1946 ( .A(\mem<29><7> ), .B(n2469), .C(\mem<28><7> ), .D(n2472), 
        .Y(n1419) );
  AOI22X1 U1947 ( .A(\mem<27><7> ), .B(n2465), .C(\mem<26><7> ), .D(n2468), 
        .Y(n1417) );
  AOI22X1 U1948 ( .A(\mem<25><7> ), .B(n2461), .C(\mem<24><7> ), .D(n2464), 
        .Y(n1416) );
  AOI21X1 U1949 ( .A(n1421), .B(n1422), .C(n2451), .Y(n3713) );
  NOR3X1 U1950 ( .A(n1423), .B(n178), .C(n187), .Y(n1422) );
  AOI22X1 U1952 ( .A(\mem<55><6> ), .B(n2577), .C(\mem<54><6> ), .D(n2580), 
        .Y(n1430) );
  AOI22X1 U1953 ( .A(\mem<53><6> ), .B(n2573), .C(\mem<52><6> ), .D(n2576), 
        .Y(n1429) );
  AOI22X1 U1954 ( .A(\mem<51><6> ), .B(n2569), .C(\mem<50><6> ), .D(n2572), 
        .Y(n1427) );
  AOI22X1 U1955 ( .A(\mem<49><6> ), .B(n2565), .C(\mem<48><6> ), .D(n2568), 
        .Y(n1426) );
  AOI22X1 U1957 ( .A(\mem<63><6> ), .B(n2459), .C(\mem<62><6> ), .D(n2564), 
        .Y(n1435) );
  AOI22X1 U1958 ( .A(\mem<61><6> ), .B(n2559), .C(\mem<60><6> ), .D(n2562), 
        .Y(n1434) );
  AOI22X1 U1959 ( .A(\mem<59><6> ), .B(n2555), .C(\mem<58><6> ), .D(n2558), 
        .Y(n1432) );
  AOI22X1 U1960 ( .A(\mem<57><6> ), .B(n2551), .C(\mem<56><6> ), .D(n2554), 
        .Y(n1431) );
  AOI22X1 U1962 ( .A(\mem<39><6> ), .B(n2547), .C(\mem<38><6> ), .D(n2550), 
        .Y(n1442) );
  AOI22X1 U1963 ( .A(\mem<37><6> ), .B(n2543), .C(\mem<36><6> ), .D(n2546), 
        .Y(n1441) );
  AOI22X1 U1964 ( .A(\mem<35><6> ), .B(n2539), .C(\mem<34><6> ), .D(n2542), 
        .Y(n1439) );
  AOI22X1 U1965 ( .A(\mem<33><6> ), .B(n2536), .C(\mem<32><6> ), .D(n2537), 
        .Y(n1438) );
  AOI22X1 U1967 ( .A(\mem<47><6> ), .B(n2531), .C(\mem<46><6> ), .D(n2534), 
        .Y(n1447) );
  AOI22X1 U1968 ( .A(\mem<45><6> ), .B(n2527), .C(\mem<44><6> ), .D(n2530), 
        .Y(n1446) );
  AOI22X1 U1969 ( .A(\mem<43><6> ), .B(n2523), .C(\mem<42><6> ), .D(n2526), 
        .Y(n1444) );
  AOI22X1 U1970 ( .A(\mem<41><6> ), .B(n2519), .C(\mem<40><6> ), .D(n2522), 
        .Y(n1443) );
  NOR3X1 U1971 ( .A(n1448), .B(n177), .C(n226), .Y(n1421) );
  AOI22X1 U1973 ( .A(\mem<7><6> ), .B(n2515), .C(\mem<6><6> ), .D(n2517), .Y(
        n1455) );
  AOI22X1 U1974 ( .A(\mem<5><6> ), .B(n2511), .C(\mem<4><6> ), .D(n2513), .Y(
        n1454) );
  AOI22X1 U1975 ( .A(\mem<3><6> ), .B(n2509), .C(\mem<2><6> ), .D(n2581), .Y(
        n1452) );
  AOI22X1 U1976 ( .A(\mem<1><6> ), .B(n2455), .C(n1403), .D(\mem<0><6> ), .Y(
        n1451) );
  AOI22X1 U1978 ( .A(\mem<15><6> ), .B(n2505), .C(\mem<14><6> ), .D(n2507), 
        .Y(n1460) );
  AOI22X1 U1979 ( .A(\mem<13><6> ), .B(n2501), .C(\mem<12><6> ), .D(n2503), 
        .Y(n1459) );
  AOI22X1 U1980 ( .A(\mem<11><6> ), .B(n2497), .C(\mem<10><6> ), .D(n2499), 
        .Y(n1457) );
  AOI22X1 U1981 ( .A(\mem<9><6> ), .B(n2493), .C(\mem<8><6> ), .D(n2495), .Y(
        n1456) );
  AOI22X1 U1983 ( .A(\mem<23><6> ), .B(n2489), .C(\mem<22><6> ), .D(n2492), 
        .Y(n1467) );
  AOI22X1 U1984 ( .A(\mem<21><6> ), .B(n2485), .C(\mem<20><6> ), .D(n2488), 
        .Y(n1466) );
  AOI22X1 U1985 ( .A(\mem<19><6> ), .B(n2481), .C(\mem<18><6> ), .D(n2484), 
        .Y(n1464) );
  AOI22X1 U1986 ( .A(\mem<17><6> ), .B(n2477), .C(\mem<16><6> ), .D(n2480), 
        .Y(n1463) );
  AOI22X1 U1988 ( .A(\mem<31><6> ), .B(n2473), .C(\mem<30><6> ), .D(n2476), 
        .Y(n1472) );
  AOI22X1 U1989 ( .A(\mem<29><6> ), .B(n2469), .C(\mem<28><6> ), .D(n2472), 
        .Y(n1471) );
  AOI22X1 U1990 ( .A(\mem<27><6> ), .B(n2465), .C(\mem<26><6> ), .D(n2468), 
        .Y(n1469) );
  AOI22X1 U1991 ( .A(\mem<25><6> ), .B(n2461), .C(\mem<24><6> ), .D(n2464), 
        .Y(n1468) );
  AOI21X1 U1992 ( .A(n1473), .B(n1474), .C(n2451), .Y(n3714) );
  NOR3X1 U1993 ( .A(n1475), .B(n176), .C(n186), .Y(n1474) );
  AOI22X1 U1995 ( .A(\mem<55><5> ), .B(n2577), .C(\mem<54><5> ), .D(n2580), 
        .Y(n1482) );
  AOI22X1 U1996 ( .A(\mem<53><5> ), .B(n2573), .C(\mem<52><5> ), .D(n2576), 
        .Y(n1481) );
  AOI22X1 U1997 ( .A(\mem<51><5> ), .B(n2569), .C(\mem<50><5> ), .D(n2572), 
        .Y(n1479) );
  AOI22X1 U1998 ( .A(\mem<49><5> ), .B(n2565), .C(\mem<48><5> ), .D(n2568), 
        .Y(n1478) );
  AOI22X1 U2000 ( .A(\mem<63><5> ), .B(n2459), .C(\mem<62><5> ), .D(n2564), 
        .Y(n1487) );
  AOI22X1 U2001 ( .A(\mem<61><5> ), .B(n2559), .C(\mem<60><5> ), .D(n2562), 
        .Y(n1486) );
  AOI22X1 U2002 ( .A(\mem<59><5> ), .B(n2555), .C(\mem<58><5> ), .D(n2558), 
        .Y(n1484) );
  AOI22X1 U2003 ( .A(\mem<57><5> ), .B(n2551), .C(\mem<56><5> ), .D(n2554), 
        .Y(n1483) );
  AOI22X1 U2005 ( .A(\mem<39><5> ), .B(n2547), .C(\mem<38><5> ), .D(n2550), 
        .Y(n1494) );
  AOI22X1 U2006 ( .A(\mem<37><5> ), .B(n2543), .C(\mem<36><5> ), .D(n2546), 
        .Y(n1493) );
  AOI22X1 U2007 ( .A(\mem<35><5> ), .B(n2539), .C(\mem<34><5> ), .D(n2542), 
        .Y(n1491) );
  AOI22X1 U2008 ( .A(\mem<33><5> ), .B(n2536), .C(\mem<32><5> ), .D(n2537), 
        .Y(n1490) );
  AOI22X1 U2010 ( .A(\mem<47><5> ), .B(n2531), .C(\mem<46><5> ), .D(n2534), 
        .Y(n1499) );
  AOI22X1 U2011 ( .A(\mem<45><5> ), .B(n2527), .C(\mem<44><5> ), .D(n2530), 
        .Y(n1498) );
  AOI22X1 U2012 ( .A(\mem<43><5> ), .B(n2523), .C(\mem<42><5> ), .D(n2526), 
        .Y(n1496) );
  AOI22X1 U2013 ( .A(\mem<41><5> ), .B(n2519), .C(\mem<40><5> ), .D(n2522), 
        .Y(n1495) );
  NOR3X1 U2014 ( .A(n1500), .B(n175), .C(n223), .Y(n1473) );
  AOI22X1 U2016 ( .A(\mem<7><5> ), .B(n2515), .C(\mem<6><5> ), .D(n2517), .Y(
        n1507) );
  AOI22X1 U2017 ( .A(\mem<5><5> ), .B(n2511), .C(\mem<4><5> ), .D(n2513), .Y(
        n1506) );
  AOI22X1 U2018 ( .A(\mem<3><5> ), .B(n2509), .C(\mem<2><5> ), .D(n2581), .Y(
        n1504) );
  AOI22X1 U2019 ( .A(\mem<1><5> ), .B(n2455), .C(n1403), .D(\mem<0><5> ), .Y(
        n1503) );
  AOI22X1 U2021 ( .A(\mem<15><5> ), .B(n2505), .C(\mem<14><5> ), .D(n2507), 
        .Y(n1512) );
  AOI22X1 U2022 ( .A(\mem<13><5> ), .B(n2501), .C(\mem<12><5> ), .D(n2503), 
        .Y(n1511) );
  AOI22X1 U2023 ( .A(\mem<11><5> ), .B(n2497), .C(\mem<10><5> ), .D(n2499), 
        .Y(n1509) );
  AOI22X1 U2024 ( .A(\mem<9><5> ), .B(n2493), .C(\mem<8><5> ), .D(n2495), .Y(
        n1508) );
  AOI22X1 U2026 ( .A(\mem<23><5> ), .B(n2489), .C(\mem<22><5> ), .D(n2492), 
        .Y(n1519) );
  AOI22X1 U2027 ( .A(\mem<21><5> ), .B(n2485), .C(\mem<20><5> ), .D(n2488), 
        .Y(n1518) );
  AOI22X1 U2028 ( .A(\mem<19><5> ), .B(n2481), .C(\mem<18><5> ), .D(n2484), 
        .Y(n1516) );
  AOI22X1 U2029 ( .A(\mem<17><5> ), .B(n2477), .C(\mem<16><5> ), .D(n2480), 
        .Y(n1515) );
  AOI22X1 U2031 ( .A(\mem<31><5> ), .B(n2473), .C(\mem<30><5> ), .D(n2476), 
        .Y(n1524) );
  AOI22X1 U2032 ( .A(\mem<29><5> ), .B(n2469), .C(\mem<28><5> ), .D(n2472), 
        .Y(n1523) );
  AOI22X1 U2033 ( .A(\mem<27><5> ), .B(n2465), .C(\mem<26><5> ), .D(n2468), 
        .Y(n1521) );
  AOI22X1 U2034 ( .A(\mem<25><5> ), .B(n2461), .C(\mem<24><5> ), .D(n2464), 
        .Y(n1520) );
  AOI21X1 U2035 ( .A(n1525), .B(n1526), .C(n2451), .Y(n3715) );
  NOR3X1 U2036 ( .A(n1527), .B(n174), .C(n185), .Y(n1526) );
  AOI22X1 U2038 ( .A(\mem<55><4> ), .B(n2577), .C(\mem<54><4> ), .D(n2580), 
        .Y(n1534) );
  AOI22X1 U2039 ( .A(\mem<53><4> ), .B(n2573), .C(\mem<52><4> ), .D(n2576), 
        .Y(n1533) );
  AOI22X1 U2040 ( .A(\mem<51><4> ), .B(n2569), .C(\mem<50><4> ), .D(n2572), 
        .Y(n1531) );
  AOI22X1 U2041 ( .A(\mem<49><4> ), .B(n2565), .C(\mem<48><4> ), .D(n2568), 
        .Y(n1530) );
  AOI22X1 U2043 ( .A(\mem<63><4> ), .B(n2459), .C(\mem<62><4> ), .D(n2564), 
        .Y(n1539) );
  AOI22X1 U2044 ( .A(\mem<61><4> ), .B(n2559), .C(\mem<60><4> ), .D(n2562), 
        .Y(n1538) );
  AOI22X1 U2045 ( .A(\mem<59><4> ), .B(n2555), .C(\mem<58><4> ), .D(n2558), 
        .Y(n1536) );
  AOI22X1 U2046 ( .A(\mem<57><4> ), .B(n2551), .C(\mem<56><4> ), .D(n2554), 
        .Y(n1535) );
  AOI22X1 U2048 ( .A(\mem<39><4> ), .B(n2547), .C(\mem<38><4> ), .D(n2550), 
        .Y(n1546) );
  AOI22X1 U2049 ( .A(\mem<37><4> ), .B(n2543), .C(\mem<36><4> ), .D(n2546), 
        .Y(n1545) );
  AOI22X1 U2050 ( .A(\mem<35><4> ), .B(n2539), .C(\mem<34><4> ), .D(n2542), 
        .Y(n1543) );
  AOI22X1 U2051 ( .A(\mem<33><4> ), .B(n2536), .C(\mem<32><4> ), .D(n2537), 
        .Y(n1542) );
  AOI22X1 U2053 ( .A(\mem<47><4> ), .B(n2531), .C(\mem<46><4> ), .D(n2534), 
        .Y(n1551) );
  AOI22X1 U2054 ( .A(\mem<45><4> ), .B(n2527), .C(\mem<44><4> ), .D(n2530), 
        .Y(n1550) );
  AOI22X1 U2055 ( .A(\mem<43><4> ), .B(n2523), .C(\mem<42><4> ), .D(n2526), 
        .Y(n1548) );
  AOI22X1 U2056 ( .A(\mem<41><4> ), .B(n2519), .C(\mem<40><4> ), .D(n2522), 
        .Y(n1547) );
  NOR3X1 U2057 ( .A(n1552), .B(n173), .C(n220), .Y(n1525) );
  AOI22X1 U2059 ( .A(\mem<7><4> ), .B(n2515), .C(\mem<6><4> ), .D(n2517), .Y(
        n1559) );
  AOI22X1 U2060 ( .A(\mem<5><4> ), .B(n2511), .C(\mem<4><4> ), .D(n2513), .Y(
        n1558) );
  AOI22X1 U2061 ( .A(\mem<3><4> ), .B(n2509), .C(\mem<2><4> ), .D(n2581), .Y(
        n1556) );
  AOI22X1 U2062 ( .A(\mem<1><4> ), .B(n2455), .C(n1403), .D(\mem<0><4> ), .Y(
        n1555) );
  AOI22X1 U2064 ( .A(\mem<15><4> ), .B(n2505), .C(\mem<14><4> ), .D(n2507), 
        .Y(n1564) );
  AOI22X1 U2065 ( .A(\mem<13><4> ), .B(n2501), .C(\mem<12><4> ), .D(n2503), 
        .Y(n1563) );
  AOI22X1 U2066 ( .A(\mem<11><4> ), .B(n2497), .C(\mem<10><4> ), .D(n2499), 
        .Y(n1561) );
  AOI22X1 U2067 ( .A(\mem<9><4> ), .B(n2493), .C(\mem<8><4> ), .D(n2495), .Y(
        n1560) );
  AOI22X1 U2069 ( .A(\mem<23><4> ), .B(n2489), .C(\mem<22><4> ), .D(n2492), 
        .Y(n1571) );
  AOI22X1 U2070 ( .A(\mem<21><4> ), .B(n2485), .C(\mem<20><4> ), .D(n2488), 
        .Y(n1570) );
  AOI22X1 U2071 ( .A(\mem<19><4> ), .B(n2481), .C(\mem<18><4> ), .D(n2484), 
        .Y(n1568) );
  AOI22X1 U2072 ( .A(\mem<17><4> ), .B(n2477), .C(\mem<16><4> ), .D(n2480), 
        .Y(n1567) );
  AOI22X1 U2074 ( .A(\mem<31><4> ), .B(n2473), .C(\mem<30><4> ), .D(n2476), 
        .Y(n1576) );
  AOI22X1 U2075 ( .A(\mem<29><4> ), .B(n2469), .C(\mem<28><4> ), .D(n2472), 
        .Y(n1575) );
  AOI22X1 U2076 ( .A(\mem<27><4> ), .B(n2465), .C(\mem<26><4> ), .D(n2468), 
        .Y(n1573) );
  AOI22X1 U2077 ( .A(\mem<25><4> ), .B(n2461), .C(\mem<24><4> ), .D(n2464), 
        .Y(n1572) );
  AOI21X1 U2078 ( .A(n1577), .B(n1578), .C(n2451), .Y(n3716) );
  NOR3X1 U2079 ( .A(n1579), .B(n172), .C(n184), .Y(n1578) );
  AOI22X1 U2081 ( .A(\mem<55><3> ), .B(n2577), .C(\mem<54><3> ), .D(n2580), 
        .Y(n1586) );
  AOI22X1 U2082 ( .A(\mem<53><3> ), .B(n2573), .C(\mem<52><3> ), .D(n2576), 
        .Y(n1585) );
  AOI22X1 U2083 ( .A(\mem<51><3> ), .B(n2569), .C(\mem<50><3> ), .D(n2572), 
        .Y(n1583) );
  AOI22X1 U2084 ( .A(\mem<49><3> ), .B(n2565), .C(\mem<48><3> ), .D(n2568), 
        .Y(n1582) );
  AOI22X1 U2086 ( .A(\mem<63><3> ), .B(n2459), .C(\mem<62><3> ), .D(n2564), 
        .Y(n1591) );
  AOI22X1 U2087 ( .A(\mem<61><3> ), .B(n2559), .C(\mem<60><3> ), .D(n2562), 
        .Y(n1590) );
  AOI22X1 U2088 ( .A(\mem<59><3> ), .B(n2555), .C(\mem<58><3> ), .D(n2558), 
        .Y(n1588) );
  AOI22X1 U2089 ( .A(\mem<57><3> ), .B(n2551), .C(\mem<56><3> ), .D(n2554), 
        .Y(n1587) );
  AOI22X1 U2091 ( .A(\mem<39><3> ), .B(n2547), .C(\mem<38><3> ), .D(n2550), 
        .Y(n1598) );
  AOI22X1 U2092 ( .A(\mem<37><3> ), .B(n2543), .C(\mem<36><3> ), .D(n2546), 
        .Y(n1597) );
  AOI22X1 U2093 ( .A(\mem<35><3> ), .B(n2539), .C(\mem<34><3> ), .D(n2542), 
        .Y(n1595) );
  AOI22X1 U2094 ( .A(\mem<33><3> ), .B(n2536), .C(\mem<32><3> ), .D(n2537), 
        .Y(n1594) );
  AOI22X1 U2096 ( .A(\mem<47><3> ), .B(n2531), .C(\mem<46><3> ), .D(n2534), 
        .Y(n1603) );
  AOI22X1 U2097 ( .A(\mem<45><3> ), .B(n2527), .C(\mem<44><3> ), .D(n2530), 
        .Y(n1602) );
  AOI22X1 U2098 ( .A(\mem<43><3> ), .B(n2523), .C(\mem<42><3> ), .D(n2526), 
        .Y(n1600) );
  AOI22X1 U2099 ( .A(\mem<41><3> ), .B(n2519), .C(\mem<40><3> ), .D(n2522), 
        .Y(n1599) );
  NOR3X1 U2100 ( .A(n1604), .B(n171), .C(n217), .Y(n1577) );
  AOI22X1 U2102 ( .A(\mem<7><3> ), .B(n2515), .C(\mem<6><3> ), .D(n2517), .Y(
        n1611) );
  AOI22X1 U2103 ( .A(\mem<5><3> ), .B(n2511), .C(\mem<4><3> ), .D(n2513), .Y(
        n1610) );
  AOI22X1 U2104 ( .A(\mem<3><3> ), .B(n2509), .C(\mem<2><3> ), .D(n2581), .Y(
        n1608) );
  AOI22X1 U2105 ( .A(\mem<1><3> ), .B(n2455), .C(n1403), .D(\mem<0><3> ), .Y(
        n1607) );
  AOI22X1 U2107 ( .A(\mem<15><3> ), .B(n2505), .C(\mem<14><3> ), .D(n2507), 
        .Y(n1616) );
  AOI22X1 U2108 ( .A(\mem<13><3> ), .B(n2501), .C(\mem<12><3> ), .D(n2503), 
        .Y(n1615) );
  AOI22X1 U2109 ( .A(\mem<11><3> ), .B(n2497), .C(\mem<10><3> ), .D(n2499), 
        .Y(n1613) );
  AOI22X1 U2110 ( .A(\mem<9><3> ), .B(n2493), .C(\mem<8><3> ), .D(n2495), .Y(
        n1612) );
  AOI22X1 U2112 ( .A(\mem<23><3> ), .B(n2489), .C(\mem<22><3> ), .D(n2492), 
        .Y(n1623) );
  AOI22X1 U2113 ( .A(\mem<21><3> ), .B(n2485), .C(\mem<20><3> ), .D(n2488), 
        .Y(n1622) );
  AOI22X1 U2114 ( .A(\mem<19><3> ), .B(n2481), .C(\mem<18><3> ), .D(n2484), 
        .Y(n1620) );
  AOI22X1 U2115 ( .A(\mem<17><3> ), .B(n2477), .C(\mem<16><3> ), .D(n2480), 
        .Y(n1619) );
  AOI22X1 U2117 ( .A(\mem<31><3> ), .B(n2473), .C(\mem<30><3> ), .D(n2476), 
        .Y(n1628) );
  AOI22X1 U2118 ( .A(\mem<29><3> ), .B(n2469), .C(\mem<28><3> ), .D(n2472), 
        .Y(n1627) );
  AOI22X1 U2119 ( .A(\mem<27><3> ), .B(n2465), .C(\mem<26><3> ), .D(n2468), 
        .Y(n1625) );
  AOI22X1 U2120 ( .A(\mem<25><3> ), .B(n2461), .C(\mem<24><3> ), .D(n2464), 
        .Y(n1624) );
  AOI21X1 U2121 ( .A(n1629), .B(n1630), .C(n2451), .Y(n3717) );
  NOR3X1 U2122 ( .A(n1631), .B(n170), .C(n183), .Y(n1630) );
  AOI22X1 U2124 ( .A(\mem<55><2> ), .B(n2577), .C(\mem<54><2> ), .D(n2580), 
        .Y(n1638) );
  AOI22X1 U2125 ( .A(\mem<53><2> ), .B(n2573), .C(\mem<52><2> ), .D(n2576), 
        .Y(n1637) );
  AOI22X1 U2126 ( .A(\mem<51><2> ), .B(n2569), .C(\mem<50><2> ), .D(n2572), 
        .Y(n1635) );
  AOI22X1 U2127 ( .A(\mem<49><2> ), .B(n2565), .C(\mem<48><2> ), .D(n2568), 
        .Y(n1634) );
  AOI22X1 U2129 ( .A(\mem<63><2> ), .B(n2459), .C(\mem<62><2> ), .D(n2564), 
        .Y(n1643) );
  AOI22X1 U2130 ( .A(\mem<61><2> ), .B(n2559), .C(\mem<60><2> ), .D(n2562), 
        .Y(n1642) );
  AOI22X1 U2131 ( .A(\mem<59><2> ), .B(n2555), .C(\mem<58><2> ), .D(n2558), 
        .Y(n1640) );
  AOI22X1 U2132 ( .A(\mem<57><2> ), .B(n2551), .C(\mem<56><2> ), .D(n2554), 
        .Y(n1639) );
  AOI22X1 U2134 ( .A(\mem<39><2> ), .B(n2547), .C(\mem<38><2> ), .D(n2550), 
        .Y(n1650) );
  AOI22X1 U2135 ( .A(\mem<37><2> ), .B(n2543), .C(\mem<36><2> ), .D(n2546), 
        .Y(n1649) );
  AOI22X1 U2136 ( .A(\mem<35><2> ), .B(n2539), .C(\mem<34><2> ), .D(n2542), 
        .Y(n1647) );
  AOI22X1 U2137 ( .A(\mem<33><2> ), .B(n2536), .C(\mem<32><2> ), .D(n2537), 
        .Y(n1646) );
  AOI22X1 U2139 ( .A(\mem<47><2> ), .B(n2531), .C(\mem<46><2> ), .D(n2534), 
        .Y(n1655) );
  AOI22X1 U2140 ( .A(\mem<45><2> ), .B(n2527), .C(\mem<44><2> ), .D(n2530), 
        .Y(n1654) );
  AOI22X1 U2141 ( .A(\mem<43><2> ), .B(n2523), .C(\mem<42><2> ), .D(n2526), 
        .Y(n1652) );
  AOI22X1 U2142 ( .A(\mem<41><2> ), .B(n2519), .C(\mem<40><2> ), .D(n2522), 
        .Y(n1651) );
  NOR3X1 U2143 ( .A(n1656), .B(n169), .C(n214), .Y(n1629) );
  AOI22X1 U2145 ( .A(\mem<7><2> ), .B(n2515), .C(\mem<6><2> ), .D(n2517), .Y(
        n1663) );
  AOI22X1 U2146 ( .A(\mem<5><2> ), .B(n2511), .C(\mem<4><2> ), .D(n2513), .Y(
        n1662) );
  AOI22X1 U2147 ( .A(\mem<3><2> ), .B(n2509), .C(\mem<2><2> ), .D(n2581), .Y(
        n1660) );
  AOI22X1 U2148 ( .A(\mem<1><2> ), .B(n2455), .C(n1403), .D(\mem<0><2> ), .Y(
        n1659) );
  AOI22X1 U2150 ( .A(\mem<15><2> ), .B(n2505), .C(\mem<14><2> ), .D(n2507), 
        .Y(n1668) );
  AOI22X1 U2151 ( .A(\mem<13><2> ), .B(n2501), .C(\mem<12><2> ), .D(n2503), 
        .Y(n1667) );
  AOI22X1 U2152 ( .A(\mem<11><2> ), .B(n2497), .C(\mem<10><2> ), .D(n2499), 
        .Y(n1665) );
  AOI22X1 U2153 ( .A(\mem<9><2> ), .B(n2493), .C(\mem<8><2> ), .D(n2495), .Y(
        n1664) );
  AOI22X1 U2155 ( .A(\mem<23><2> ), .B(n2489), .C(\mem<22><2> ), .D(n2492), 
        .Y(n1675) );
  AOI22X1 U2156 ( .A(\mem<21><2> ), .B(n2485), .C(\mem<20><2> ), .D(n2488), 
        .Y(n1674) );
  AOI22X1 U2157 ( .A(\mem<19><2> ), .B(n2481), .C(\mem<18><2> ), .D(n2484), 
        .Y(n1672) );
  AOI22X1 U2158 ( .A(\mem<17><2> ), .B(n2477), .C(\mem<16><2> ), .D(n2480), 
        .Y(n1671) );
  AOI22X1 U2160 ( .A(\mem<31><2> ), .B(n2473), .C(\mem<30><2> ), .D(n2476), 
        .Y(n1680) );
  AOI22X1 U2161 ( .A(\mem<29><2> ), .B(n2469), .C(\mem<28><2> ), .D(n2472), 
        .Y(n1679) );
  AOI22X1 U2162 ( .A(\mem<27><2> ), .B(n2465), .C(\mem<26><2> ), .D(n2468), 
        .Y(n1677) );
  AOI22X1 U2163 ( .A(\mem<25><2> ), .B(n2461), .C(\mem<24><2> ), .D(n2464), 
        .Y(n1676) );
  AOI21X1 U2164 ( .A(n1681), .B(n1682), .C(n2451), .Y(n3718) );
  NOR3X1 U2165 ( .A(n1683), .B(n168), .C(n182), .Y(n1682) );
  AOI22X1 U2167 ( .A(\mem<55><1> ), .B(n2577), .C(\mem<54><1> ), .D(n2580), 
        .Y(n1690) );
  AOI22X1 U2168 ( .A(\mem<53><1> ), .B(n2573), .C(\mem<52><1> ), .D(n2576), 
        .Y(n1689) );
  AOI22X1 U2169 ( .A(\mem<51><1> ), .B(n2569), .C(\mem<50><1> ), .D(n2572), 
        .Y(n1687) );
  AOI22X1 U2170 ( .A(\mem<49><1> ), .B(n2565), .C(\mem<48><1> ), .D(n2568), 
        .Y(n1686) );
  AOI22X1 U2172 ( .A(\mem<63><1> ), .B(n2459), .C(\mem<62><1> ), .D(n2564), 
        .Y(n1695) );
  AOI22X1 U2173 ( .A(\mem<61><1> ), .B(n2559), .C(\mem<60><1> ), .D(n2562), 
        .Y(n1694) );
  AOI22X1 U2174 ( .A(\mem<59><1> ), .B(n2555), .C(\mem<58><1> ), .D(n2558), 
        .Y(n1692) );
  AOI22X1 U2175 ( .A(\mem<57><1> ), .B(n2551), .C(\mem<56><1> ), .D(n2554), 
        .Y(n1691) );
  AOI22X1 U2177 ( .A(\mem<39><1> ), .B(n2547), .C(\mem<38><1> ), .D(n2550), 
        .Y(n1702) );
  AOI22X1 U2178 ( .A(\mem<37><1> ), .B(n2543), .C(\mem<36><1> ), .D(n2546), 
        .Y(n1701) );
  AOI22X1 U2179 ( .A(\mem<35><1> ), .B(n2539), .C(\mem<34><1> ), .D(n2542), 
        .Y(n1699) );
  AOI22X1 U2180 ( .A(\mem<33><1> ), .B(n2536), .C(\mem<32><1> ), .D(n2537), 
        .Y(n1698) );
  AOI22X1 U2182 ( .A(\mem<47><1> ), .B(n2531), .C(\mem<46><1> ), .D(n2534), 
        .Y(n1707) );
  AOI22X1 U2183 ( .A(\mem<45><1> ), .B(n2527), .C(\mem<44><1> ), .D(n2530), 
        .Y(n1706) );
  AOI22X1 U2184 ( .A(\mem<43><1> ), .B(n2523), .C(\mem<42><1> ), .D(n2526), 
        .Y(n1704) );
  AOI22X1 U2185 ( .A(\mem<41><1> ), .B(n2519), .C(\mem<40><1> ), .D(n2522), 
        .Y(n1703) );
  NOR3X1 U2186 ( .A(n1708), .B(n167), .C(n211), .Y(n1681) );
  AOI22X1 U2188 ( .A(\mem<7><1> ), .B(n2515), .C(\mem<6><1> ), .D(n2517), .Y(
        n1715) );
  AOI22X1 U2189 ( .A(\mem<5><1> ), .B(n2511), .C(\mem<4><1> ), .D(n2513), .Y(
        n1714) );
  AOI22X1 U2190 ( .A(\mem<3><1> ), .B(n2509), .C(\mem<2><1> ), .D(n2581), .Y(
        n1712) );
  AOI22X1 U2191 ( .A(\mem<1><1> ), .B(n2455), .C(n1403), .D(\mem<0><1> ), .Y(
        n1711) );
  AOI22X1 U2193 ( .A(\mem<15><1> ), .B(n2505), .C(\mem<14><1> ), .D(n2507), 
        .Y(n1720) );
  AOI22X1 U2194 ( .A(\mem<13><1> ), .B(n2501), .C(\mem<12><1> ), .D(n2503), 
        .Y(n1719) );
  AOI22X1 U2195 ( .A(\mem<11><1> ), .B(n2497), .C(\mem<10><1> ), .D(n2499), 
        .Y(n1717) );
  AOI22X1 U2196 ( .A(\mem<9><1> ), .B(n2493), .C(\mem<8><1> ), .D(n2495), .Y(
        n1716) );
  AOI22X1 U2198 ( .A(\mem<23><1> ), .B(n2489), .C(\mem<22><1> ), .D(n2492), 
        .Y(n1727) );
  AOI22X1 U2199 ( .A(\mem<21><1> ), .B(n2485), .C(\mem<20><1> ), .D(n2488), 
        .Y(n1726) );
  AOI22X1 U2200 ( .A(\mem<19><1> ), .B(n2481), .C(\mem<18><1> ), .D(n2484), 
        .Y(n1724) );
  AOI22X1 U2201 ( .A(\mem<17><1> ), .B(n2477), .C(\mem<16><1> ), .D(n2480), 
        .Y(n1723) );
  AOI22X1 U2203 ( .A(\mem<31><1> ), .B(n2473), .C(\mem<30><1> ), .D(n2476), 
        .Y(n1732) );
  AOI22X1 U2204 ( .A(\mem<29><1> ), .B(n2469), .C(\mem<28><1> ), .D(n2472), 
        .Y(n1731) );
  AOI22X1 U2205 ( .A(\mem<27><1> ), .B(n2465), .C(\mem<26><1> ), .D(n2468), 
        .Y(n1729) );
  AOI22X1 U2206 ( .A(\mem<25><1> ), .B(n2461), .C(\mem<24><1> ), .D(n2464), 
        .Y(n1728) );
  AOI21X1 U2207 ( .A(n1733), .B(n1734), .C(n2451), .Y(n3719) );
  NOR3X1 U2209 ( .A(n1735), .B(n166), .C(n181), .Y(n1734) );
  AOI22X1 U2211 ( .A(\mem<55><0> ), .B(n2577), .C(\mem<54><0> ), .D(n2580), 
        .Y(n1742) );
  AOI22X1 U2214 ( .A(\mem<53><0> ), .B(n2573), .C(\mem<52><0> ), .D(n2576), 
        .Y(n1741) );
  AOI22X1 U2217 ( .A(\mem<51><0> ), .B(n2569), .C(\mem<50><0> ), .D(n2572), 
        .Y(n1739) );
  AOI22X1 U2220 ( .A(\mem<49><0> ), .B(n2565), .C(\mem<48><0> ), .D(n2568), 
        .Y(n1738) );
  AOI22X1 U2224 ( .A(\mem<63><0> ), .B(n2459), .C(\mem<62><0> ), .D(n2564), 
        .Y(n1754) );
  AOI22X1 U2227 ( .A(\mem<61><0> ), .B(n2559), .C(\mem<60><0> ), .D(n2562), 
        .Y(n1753) );
  AOI22X1 U2230 ( .A(\mem<59><0> ), .B(n2555), .C(\mem<58><0> ), .D(n2558), 
        .Y(n1751) );
  AOI22X1 U2233 ( .A(\mem<57><0> ), .B(n2551), .C(\mem<56><0> ), .D(n2554), 
        .Y(n1750) );
  NAND3X1 U2235 ( .A(n1756), .B(N182), .C(n1757), .Y(n1755) );
  AOI22X1 U2239 ( .A(\mem<39><0> ), .B(n2547), .C(\mem<38><0> ), .D(n2550), 
        .Y(n1764) );
  AOI22X1 U2242 ( .A(\mem<37><0> ), .B(n2543), .C(\mem<36><0> ), .D(n2546), 
        .Y(n1763) );
  AOI22X1 U2245 ( .A(\mem<35><0> ), .B(n2539), .C(\mem<34><0> ), .D(n2542), 
        .Y(n1761) );
  AOI22X1 U2248 ( .A(\mem<33><0> ), .B(n2536), .C(\mem<32><0> ), .D(n2537), 
        .Y(n1760) );
  AOI22X1 U2252 ( .A(\mem<47><0> ), .B(n2531), .C(\mem<46><0> ), .D(n2534), 
        .Y(n1769) );
  AOI22X1 U2255 ( .A(\mem<45><0> ), .B(n2527), .C(\mem<44><0> ), .D(n2530), 
        .Y(n1768) );
  AOI22X1 U2258 ( .A(\mem<43><0> ), .B(n2523), .C(\mem<42><0> ), .D(n2526), 
        .Y(n1766) );
  AOI22X1 U2261 ( .A(\mem<41><0> ), .B(n2519), .C(\mem<40><0> ), .D(n2522), 
        .Y(n1765) );
  NAND3X1 U2263 ( .A(n1756), .B(N182), .C(n2353), .Y(n1770) );
  NAND3X1 U2266 ( .A(n1756), .B(N182), .C(n2351), .Y(n1772) );
  NOR3X1 U2268 ( .A(n1774), .B(n165), .C(n208), .Y(n1733) );
  AOI22X1 U2270 ( .A(\mem<7><0> ), .B(n2515), .C(\mem<6><0> ), .D(n2517), .Y(
        n1781) );
  AOI22X1 U2273 ( .A(\mem<5><0> ), .B(n2511), .C(\mem<4><0> ), .D(n2513), .Y(
        n1780) );
  AOI22X1 U2276 ( .A(\mem<3><0> ), .B(n2509), .C(\mem<2><0> ), .D(n2581), .Y(
        n1778) );
  AOI22X1 U2279 ( .A(\mem<1><0> ), .B(n2455), .C(n1403), .D(\mem<0><0> ), .Y(
        n1777) );
  NOR3X1 U2280 ( .A(n1782), .B(n1783), .C(n1784), .Y(n1403) );
  NAND3X1 U2281 ( .A(\addr<8> ), .B(\addr<7> ), .C(\addr<9> ), .Y(n1786) );
  NAND3X1 U2282 ( .A(\addr<15> ), .B(\addr<14> ), .C(\addr<6> ), .Y(n1785) );
  NAND3X1 U2283 ( .A(\addr<10> ), .B(n3195), .C(n3189), .Y(n1783) );
  NAND3X1 U2284 ( .A(N181), .B(N180), .C(N182), .Y(n1787) );
  NAND3X1 U2285 ( .A(\addr<13> ), .B(\addr<11> ), .C(\addr<12> ), .Y(n1782) );
  AOI22X1 U2288 ( .A(\mem<15><0> ), .B(n2505), .C(\mem<14><0> ), .D(n2507), 
        .Y(n1792) );
  AOI22X1 U2291 ( .A(\mem<13><0> ), .B(n2501), .C(\mem<12><0> ), .D(n2503), 
        .Y(n1791) );
  AOI22X1 U2294 ( .A(\mem<11><0> ), .B(n2497), .C(\mem<10><0> ), .D(n2499), 
        .Y(n1789) );
  AOI22X1 U2297 ( .A(\mem<9><0> ), .B(n2493), .C(\mem<8><0> ), .D(n2495), .Y(
        n1788) );
  AOI22X1 U2302 ( .A(\mem<23><0> ), .B(n2489), .C(\mem<22><0> ), .D(n2492), 
        .Y(n1801) );
  AOI22X1 U2305 ( .A(\mem<21><0> ), .B(n2485), .C(\mem<20><0> ), .D(n2488), 
        .Y(n1800) );
  AOI22X1 U2308 ( .A(\mem<19><0> ), .B(n2481), .C(\mem<18><0> ), .D(n2484), 
        .Y(n1798) );
  AOI22X1 U2311 ( .A(\mem<17><0> ), .B(n2477), .C(\mem<16><0> ), .D(n2480), 
        .Y(n1797) );
  AOI22X1 U2317 ( .A(\mem<31><0> ), .B(n2473), .C(\mem<30><0> ), .D(n2476), 
        .Y(n1807) );
  NOR3X1 U2319 ( .A(n3079), .B(n3185), .C(n3184), .Y(n1743) );
  NOR3X1 U2321 ( .A(n3186), .B(N177), .C(n3079), .Y(n1744) );
  AOI22X1 U2322 ( .A(\mem<29><0> ), .B(n2469), .C(\mem<28><0> ), .D(n2472), 
        .Y(n1806) );
  NOR3X1 U2324 ( .A(n3186), .B(N179), .C(n3184), .Y(n1745) );
  NOR3X1 U2326 ( .A(N177), .B(n3185), .C(n3079), .Y(n1746) );
  AOI22X1 U2327 ( .A(\mem<27><0> ), .B(n2465), .C(\mem<26><0> ), .D(n2468), 
        .Y(n1804) );
  NOR3X1 U2329 ( .A(n3185), .B(N179), .C(n3184), .Y(n1747) );
  NOR3X1 U2331 ( .A(N177), .B(N179), .C(n3186), .Y(n1748) );
  AOI22X1 U2332 ( .A(\mem<25><0> ), .B(n2461), .C(\mem<24><0> ), .D(n2464), 
        .Y(n1803) );
  NAND3X1 U2334 ( .A(N179), .B(n3185), .C(N177), .Y(n612) );
  NAND3X1 U2335 ( .A(n1756), .B(N181), .C(n1809), .Y(n1808) );
  NOR2X1 U2336 ( .A(N182), .B(N180), .Y(n1809) );
  NOR3X1 U2338 ( .A(n3185), .B(N179), .C(N177), .Y(n1749) );
  NAND3X1 U2339 ( .A(n1811), .B(N181), .C(n1756), .Y(n1810) );
  NOR2X1 U2340 ( .A(N182), .B(n3187), .Y(n1811) );
  NOR3X1 U2341 ( .A(n3197), .B(\addr<6> ), .C(\addr<15> ), .Y(n1813) );
  NOR3X1 U2342 ( .A(\addr<8> ), .B(\addr<9> ), .C(\addr<7> ), .Y(n1814) );
  NOR3X1 U2343 ( .A(n3198), .B(\addr<11> ), .C(\addr<10> ), .Y(n1812) );
  NOR3X1 U2344 ( .A(\addr<13> ), .B(\addr<14> ), .C(\addr<12> ), .Y(n1815) );
  AND2X1 U3 ( .A(n1812), .B(n1813), .Y(n1756) );
  INVX1 U4 ( .A(n1815), .Y(n3198) );
  BUFX2 U5 ( .A(n1346), .Y(n3114) );
  OR2X1 U6 ( .A(n8), .B(n9), .Y(n7) );
  OR2X1 U7 ( .A(n18), .B(n19), .Y(n17) );
  OR2X1 U8 ( .A(n28), .B(n29), .Y(n27) );
  OR2X1 U9 ( .A(n38), .B(n39), .Y(n37) );
  OR2X1 U10 ( .A(n48), .B(n49), .Y(n47) );
  OR2X1 U11 ( .A(n58), .B(n59), .Y(n57) );
  OR2X1 U12 ( .A(n68), .B(n69), .Y(n67) );
  OR2X1 U13 ( .A(n78), .B(n79), .Y(n77) );
  OR2X1 U14 ( .A(n88), .B(n89), .Y(n87) );
  OR2X1 U15 ( .A(n98), .B(n99), .Y(n97) );
  OR2X1 U16 ( .A(n108), .B(n109), .Y(n107) );
  OR2X1 U17 ( .A(n118), .B(n119), .Y(n117) );
  OR2X1 U18 ( .A(n128), .B(n129), .Y(n127) );
  OR2X1 U19 ( .A(n138), .B(n139), .Y(n137) );
  OR2X1 U20 ( .A(n148), .B(n149), .Y(n147) );
  OR2X1 U21 ( .A(n158), .B(n159), .Y(n157) );
  AND2X1 U22 ( .A(N189), .B(n2450), .Y(\data_out<11> ) );
  AND2X1 U23 ( .A(n3183), .B(n610), .Y(n598) );
  AND2X1 U24 ( .A(n598), .B(n2460), .Y(n600) );
  AND2X1 U25 ( .A(n2459), .B(n598), .Y(n601) );
  AND2X1 U26 ( .A(n3175), .B(n2563), .Y(n615) );
  AND2X1 U27 ( .A(n2564), .B(n3175), .Y(n616) );
  AND2X1 U28 ( .A(n3174), .B(n2560), .Y(n628) );
  AND2X1 U29 ( .A(n2559), .B(n3174), .Y(n629) );
  AND2X1 U30 ( .A(n3173), .B(n2561), .Y(n640) );
  AND2X1 U31 ( .A(n2562), .B(n3173), .Y(n641) );
  AND2X1 U32 ( .A(n3172), .B(n2556), .Y(n652) );
  AND2X1 U33 ( .A(n2555), .B(n3172), .Y(n653) );
  AND2X1 U34 ( .A(n3171), .B(n2557), .Y(n664) );
  AND2X1 U35 ( .A(n2558), .B(n3171), .Y(n665) );
  AND2X1 U36 ( .A(n3170), .B(n2552), .Y(n676) );
  AND2X1 U37 ( .A(n2551), .B(n3170), .Y(n677) );
  AND2X1 U38 ( .A(n3169), .B(n2553), .Y(n688) );
  AND2X1 U39 ( .A(n2554), .B(n3169), .Y(n689) );
  AND2X1 U40 ( .A(n3168), .B(n2578), .Y(n700) );
  AND2X1 U41 ( .A(n2577), .B(n3168), .Y(n701) );
  AND2X1 U42 ( .A(n3167), .B(n2579), .Y(n712) );
  AND2X1 U43 ( .A(n2580), .B(n3167), .Y(n713) );
  AND2X1 U44 ( .A(n3166), .B(n2574), .Y(n724) );
  AND2X1 U45 ( .A(n2573), .B(n3166), .Y(n725) );
  AND2X1 U46 ( .A(n3165), .B(n2575), .Y(n736) );
  AND2X1 U47 ( .A(n2576), .B(n3165), .Y(n737) );
  AND2X1 U48 ( .A(n3164), .B(n2570), .Y(n748) );
  AND2X1 U49 ( .A(n2569), .B(n3164), .Y(n749) );
  AND2X1 U50 ( .A(n3163), .B(n2571), .Y(n760) );
  AND2X1 U51 ( .A(n2572), .B(n3163), .Y(n761) );
  AND2X1 U52 ( .A(n3162), .B(n2566), .Y(n772) );
  AND2X1 U53 ( .A(n2565), .B(n3162), .Y(n773) );
  AND2X1 U54 ( .A(n3161), .B(n2567), .Y(n784) );
  AND2X1 U55 ( .A(n2568), .B(n3161), .Y(n785) );
  AND2X1 U56 ( .A(n3160), .B(n2532), .Y(n796) );
  AND2X1 U57 ( .A(n2531), .B(n3160), .Y(n797) );
  AND2X1 U58 ( .A(n3159), .B(n2533), .Y(n808) );
  AND2X1 U59 ( .A(n2534), .B(n3159), .Y(n809) );
  AND2X1 U60 ( .A(n3158), .B(n2528), .Y(n820) );
  AND2X1 U61 ( .A(n2527), .B(n3158), .Y(n821) );
  AND2X1 U62 ( .A(n3157), .B(n2529), .Y(n832) );
  AND2X1 U63 ( .A(n2530), .B(n3157), .Y(n833) );
  AND2X1 U64 ( .A(n3156), .B(n2524), .Y(n844) );
  AND2X1 U65 ( .A(n2523), .B(n3156), .Y(n845) );
  AND2X1 U66 ( .A(n3155), .B(n2525), .Y(n856) );
  AND2X1 U67 ( .A(n2526), .B(n3155), .Y(n857) );
  AND2X1 U68 ( .A(n3154), .B(n2520), .Y(n868) );
  AND2X1 U69 ( .A(n2519), .B(n3154), .Y(n869) );
  AND2X1 U70 ( .A(n3153), .B(n2521), .Y(n880) );
  AND2X1 U71 ( .A(n2522), .B(n3153), .Y(n881) );
  AND2X1 U72 ( .A(n3152), .B(n2548), .Y(n892) );
  AND2X1 U73 ( .A(n2547), .B(n3152), .Y(n893) );
  AND2X1 U74 ( .A(n3151), .B(n2549), .Y(n904) );
  AND2X1 U75 ( .A(n2550), .B(n3151), .Y(n905) );
  AND2X1 U76 ( .A(n3150), .B(n2544), .Y(n916) );
  AND2X1 U77 ( .A(n2543), .B(n3150), .Y(n917) );
  AND2X1 U78 ( .A(n3149), .B(n2545), .Y(n928) );
  AND2X1 U79 ( .A(n2546), .B(n3149), .Y(n929) );
  AND2X1 U80 ( .A(n3148), .B(n2540), .Y(n940) );
  AND2X1 U81 ( .A(n2539), .B(n3148), .Y(n941) );
  AND2X1 U82 ( .A(n3147), .B(n2541), .Y(n952) );
  AND2X1 U83 ( .A(n2542), .B(n3147), .Y(n953) );
  AND2X1 U84 ( .A(n3146), .B(n2535), .Y(n964) );
  AND2X1 U85 ( .A(n2536), .B(n3146), .Y(n965) );
  AND2X1 U86 ( .A(n3145), .B(n2538), .Y(n976) );
  AND2X1 U87 ( .A(n2537), .B(n3145), .Y(n977) );
  AND2X1 U88 ( .A(n3144), .B(n2474), .Y(n988) );
  AND2X1 U89 ( .A(n2473), .B(n3144), .Y(n989) );
  AND2X1 U90 ( .A(n3143), .B(n2475), .Y(n1000) );
  AND2X1 U91 ( .A(n2476), .B(n3143), .Y(n1001) );
  AND2X1 U92 ( .A(n3142), .B(n2470), .Y(n1012) );
  AND2X1 U93 ( .A(n2469), .B(n3142), .Y(n1013) );
  AND2X1 U94 ( .A(n3141), .B(n2471), .Y(n1024) );
  AND2X1 U95 ( .A(n2472), .B(n3141), .Y(n1025) );
  AND2X1 U96 ( .A(n3140), .B(n2466), .Y(n1036) );
  AND2X1 U97 ( .A(n2465), .B(n3140), .Y(n1037) );
  AND2X1 U98 ( .A(n3139), .B(n2467), .Y(n1048) );
  AND2X1 U99 ( .A(n2468), .B(n3139), .Y(n1049) );
  AND2X1 U100 ( .A(n3138), .B(n2462), .Y(n1060) );
  AND2X1 U101 ( .A(n2461), .B(n3138), .Y(n1061) );
  AND2X1 U102 ( .A(n3137), .B(n2463), .Y(n1072) );
  AND2X1 U103 ( .A(n2464), .B(n3137), .Y(n1073) );
  AND2X1 U104 ( .A(n3136), .B(n2490), .Y(n1084) );
  AND2X1 U105 ( .A(n2489), .B(n3136), .Y(n1085) );
  AND2X1 U106 ( .A(n3135), .B(n2491), .Y(n1096) );
  AND2X1 U107 ( .A(n2492), .B(n3135), .Y(n1097) );
  AND2X1 U108 ( .A(n3134), .B(n2486), .Y(n1108) );
  AND2X1 U109 ( .A(n2485), .B(n3134), .Y(n1109) );
  AND2X1 U110 ( .A(n3133), .B(n2487), .Y(n1120) );
  AND2X1 U111 ( .A(n2488), .B(n3133), .Y(n1121) );
  AND2X1 U112 ( .A(n3132), .B(n2482), .Y(n1132) );
  AND2X1 U113 ( .A(n2481), .B(n3132), .Y(n1133) );
  AND2X1 U114 ( .A(n3131), .B(n2483), .Y(n1144) );
  AND2X1 U115 ( .A(n2484), .B(n3131), .Y(n1145) );
  AND2X1 U116 ( .A(n3130), .B(n2478), .Y(n1156) );
  AND2X1 U117 ( .A(n2477), .B(n3130), .Y(n1157) );
  AND2X1 U118 ( .A(n3129), .B(n2479), .Y(n1168) );
  AND2X1 U119 ( .A(n2480), .B(n3129), .Y(n1169) );
  AND2X1 U120 ( .A(n3128), .B(n2506), .Y(n1180) );
  AND2X1 U121 ( .A(n2505), .B(n3128), .Y(n1181) );
  AND2X1 U122 ( .A(n3127), .B(n2508), .Y(n1192) );
  AND2X1 U123 ( .A(n2507), .B(n3127), .Y(n1193) );
  AND2X1 U124 ( .A(n3126), .B(n2502), .Y(n1204) );
  AND2X1 U125 ( .A(n2501), .B(n3126), .Y(n1205) );
  AND2X1 U126 ( .A(n3125), .B(n2504), .Y(n1216) );
  AND2X1 U127 ( .A(n2503), .B(n3125), .Y(n1217) );
  AND2X1 U128 ( .A(n3124), .B(n2498), .Y(n1228) );
  AND2X1 U129 ( .A(n2497), .B(n3124), .Y(n1229) );
  AND2X1 U130 ( .A(n3123), .B(n2500), .Y(n1240) );
  AND2X1 U131 ( .A(n2499), .B(n3123), .Y(n1241) );
  AND2X1 U134 ( .A(n3122), .B(n2494), .Y(n1252) );
  AND2X1 U139 ( .A(n2493), .B(n3122), .Y(n1253) );
  AND2X1 U144 ( .A(n3121), .B(n2496), .Y(n1264) );
  AND2X1 U149 ( .A(n2495), .B(n3121), .Y(n1265) );
  AND2X1 U154 ( .A(n3120), .B(n2516), .Y(n1276) );
  AND2X1 U159 ( .A(n2515), .B(n3120), .Y(n1277) );
  AND2X1 U164 ( .A(n3119), .B(n2518), .Y(n1288) );
  AND2X1 U169 ( .A(n2517), .B(n3119), .Y(n1289) );
  AND2X1 U174 ( .A(n3118), .B(n2512), .Y(n1300) );
  AND2X1 U179 ( .A(n2511), .B(n3118), .Y(n1301) );
  AND2X1 U184 ( .A(n3117), .B(n2514), .Y(n1312) );
  AND2X1 U189 ( .A(n2513), .B(n3117), .Y(n1313) );
  AND2X1 U194 ( .A(n3116), .B(n2510), .Y(n1324) );
  AND2X1 U199 ( .A(n2509), .B(n3116), .Y(n1325) );
  AND2X1 U202 ( .A(n3115), .B(n2582), .Y(n1336) );
  AND2X1 U203 ( .A(n2581), .B(n3115), .Y(n1337) );
  AND2X1 U204 ( .A(n3114), .B(n2456), .Y(n1348) );
  AND2X1 U205 ( .A(n2455), .B(n3114), .Y(n1349) );
  INVX1 U206 ( .A(n2458), .Y(n3190) );
  INVX1 U207 ( .A(n3094), .Y(n3102) );
  INVX1 U210 ( .A(n3094), .Y(n3103) );
  INVX1 U211 ( .A(n3093), .Y(n3104) );
  INVX1 U217 ( .A(n3093), .Y(n3105) );
  INVX1 U220 ( .A(n3093), .Y(n3106) );
  INVX1 U221 ( .A(n3092), .Y(n3107) );
  INVX1 U222 ( .A(n3092), .Y(n3108) );
  INVX1 U223 ( .A(n3092), .Y(n3109) );
  INVX1 U224 ( .A(n3091), .Y(n3110) );
  INVX1 U225 ( .A(n3091), .Y(n3112) );
  INVX1 U226 ( .A(n3091), .Y(n3111) );
  INVX1 U227 ( .A(n1814), .Y(n3197) );
  AND2X1 U228 ( .A(n3187), .B(N181), .Y(n1757) );
  OR2X1 U229 ( .A(n2341), .B(n190), .Y(n161) );
  OR2X1 U230 ( .A(n2341), .B(n191), .Y(n163) );
  OR2X1 U231 ( .A(n1), .B(n6), .Y(n1774) );
  OR2X1 U232 ( .A(n11), .B(n16), .Y(n1735) );
  OR2X1 U233 ( .A(n21), .B(n26), .Y(n1708) );
  OR2X1 U234 ( .A(n31), .B(n36), .Y(n1683) );
  OR2X1 U235 ( .A(n41), .B(n46), .Y(n1656) );
  OR2X1 U236 ( .A(n51), .B(n56), .Y(n1631) );
  OR2X1 U237 ( .A(n61), .B(n66), .Y(n1604) );
  OR2X1 U238 ( .A(n71), .B(n76), .Y(n1579) );
  OR2X1 U239 ( .A(n81), .B(n86), .Y(n1552) );
  OR2X1 U240 ( .A(n91), .B(n96), .Y(n1527) );
  OR2X1 U241 ( .A(n101), .B(n106), .Y(n1500) );
  OR2X1 U242 ( .A(n111), .B(n116), .Y(n1475) );
  OR2X1 U243 ( .A(n121), .B(n126), .Y(n1448) );
  OR2X1 U244 ( .A(n131), .B(n136), .Y(n1423) );
  OR2X1 U245 ( .A(n141), .B(n146), .Y(n1395) );
  OR2X1 U246 ( .A(n151), .B(n156), .Y(n1370) );
  INVX1 U247 ( .A(wr), .Y(n3711) );
  INVX2 U248 ( .A(n2452), .Y(n3182) );
  INVX2 U249 ( .A(n2452), .Y(n3181) );
  AND2X1 U250 ( .A(N192), .B(n2450), .Y(\data_out<8> ) );
  AND2X1 U251 ( .A(N191), .B(n2450), .Y(\data_out<9> ) );
  AND2X1 U252 ( .A(N190), .B(n2450), .Y(\data_out<10> ) );
  AND2X1 U253 ( .A(N188), .B(n2450), .Y(\data_out<12> ) );
  AND2X1 U254 ( .A(N187), .B(n2450), .Y(\data_out<13> ) );
  AND2X1 U255 ( .A(N186), .B(n2450), .Y(\data_out<14> ) );
  AND2X1 U256 ( .A(N185), .B(n2450), .Y(\data_out<15> ) );
  INVX1 U257 ( .A(\mem<63><0> ), .Y(n3710) );
  INVX1 U258 ( .A(\mem<63><1> ), .Y(n3709) );
  INVX1 U259 ( .A(\mem<63><2> ), .Y(n3708) );
  INVX1 U260 ( .A(\mem<63><3> ), .Y(n3707) );
  INVX1 U261 ( .A(\mem<63><4> ), .Y(n3706) );
  INVX1 U262 ( .A(\mem<63><5> ), .Y(n3705) );
  INVX1 U263 ( .A(\mem<63><6> ), .Y(n3704) );
  INVX1 U264 ( .A(\mem<63><7> ), .Y(n3703) );
  INVX1 U265 ( .A(\mem<62><0> ), .Y(n3702) );
  INVX1 U266 ( .A(\mem<62><1> ), .Y(n3701) );
  INVX1 U267 ( .A(\mem<62><2> ), .Y(n3700) );
  INVX1 U268 ( .A(\mem<62><3> ), .Y(n3699) );
  INVX1 U269 ( .A(\mem<62><4> ), .Y(n3698) );
  INVX1 U270 ( .A(\mem<62><5> ), .Y(n3697) );
  INVX1 U271 ( .A(\mem<62><6> ), .Y(n3696) );
  INVX1 U272 ( .A(\mem<62><7> ), .Y(n3695) );
  INVX1 U273 ( .A(\mem<61><0> ), .Y(n3694) );
  INVX1 U274 ( .A(\mem<61><1> ), .Y(n3693) );
  INVX1 U275 ( .A(\mem<61><2> ), .Y(n3692) );
  INVX1 U276 ( .A(\mem<61><3> ), .Y(n3691) );
  INVX1 U277 ( .A(\mem<61><4> ), .Y(n3690) );
  INVX1 U278 ( .A(\mem<61><5> ), .Y(n3689) );
  INVX1 U279 ( .A(\mem<61><6> ), .Y(n3688) );
  INVX1 U280 ( .A(\mem<61><7> ), .Y(n3687) );
  INVX1 U281 ( .A(\mem<60><0> ), .Y(n3686) );
  INVX1 U282 ( .A(\mem<60><1> ), .Y(n3685) );
  INVX1 U283 ( .A(\mem<60><2> ), .Y(n3684) );
  INVX1 U284 ( .A(\mem<60><3> ), .Y(n3683) );
  INVX1 U285 ( .A(\mem<60><4> ), .Y(n3682) );
  INVX1 U286 ( .A(\mem<60><5> ), .Y(n3681) );
  INVX1 U287 ( .A(\mem<60><6> ), .Y(n3680) );
  INVX1 U288 ( .A(\mem<60><7> ), .Y(n3679) );
  INVX1 U289 ( .A(\mem<59><0> ), .Y(n3678) );
  INVX1 U290 ( .A(\mem<59><1> ), .Y(n3677) );
  INVX1 U291 ( .A(\mem<59><2> ), .Y(n3676) );
  INVX1 U292 ( .A(\mem<59><3> ), .Y(n3675) );
  INVX1 U293 ( .A(\mem<59><4> ), .Y(n3674) );
  INVX1 U294 ( .A(\mem<59><5> ), .Y(n3673) );
  INVX1 U295 ( .A(\mem<59><6> ), .Y(n3672) );
  INVX1 U296 ( .A(\mem<59><7> ), .Y(n3671) );
  INVX1 U297 ( .A(\mem<58><0> ), .Y(n3670) );
  INVX1 U298 ( .A(\mem<58><1> ), .Y(n3669) );
  INVX1 U299 ( .A(\mem<58><2> ), .Y(n3668) );
  INVX1 U300 ( .A(\mem<58><3> ), .Y(n3667) );
  INVX1 U301 ( .A(\mem<58><4> ), .Y(n3666) );
  INVX1 U302 ( .A(\mem<58><5> ), .Y(n3665) );
  INVX1 U303 ( .A(\mem<58><6> ), .Y(n3664) );
  INVX1 U304 ( .A(\mem<58><7> ), .Y(n3663) );
  INVX1 U305 ( .A(\mem<57><0> ), .Y(n3662) );
  INVX1 U306 ( .A(\mem<57><1> ), .Y(n3661) );
  INVX1 U307 ( .A(\mem<57><2> ), .Y(n3660) );
  INVX1 U308 ( .A(\mem<57><3> ), .Y(n3659) );
  INVX1 U309 ( .A(\mem<57><4> ), .Y(n3658) );
  INVX1 U310 ( .A(\mem<57><5> ), .Y(n3657) );
  INVX1 U311 ( .A(\mem<57><6> ), .Y(n3656) );
  INVX1 U312 ( .A(\mem<57><7> ), .Y(n3655) );
  INVX1 U313 ( .A(\mem<56><0> ), .Y(n3654) );
  INVX1 U314 ( .A(\mem<56><1> ), .Y(n3653) );
  INVX1 U315 ( .A(\mem<56><2> ), .Y(n3652) );
  INVX1 U316 ( .A(\mem<56><3> ), .Y(n3651) );
  INVX1 U317 ( .A(\mem<56><4> ), .Y(n3650) );
  INVX1 U318 ( .A(\mem<56><5> ), .Y(n3649) );
  INVX1 U319 ( .A(\mem<56><6> ), .Y(n3648) );
  INVX1 U320 ( .A(\mem<56><7> ), .Y(n3647) );
  INVX1 U321 ( .A(\mem<55><0> ), .Y(n3646) );
  INVX1 U322 ( .A(\mem<55><1> ), .Y(n3645) );
  INVX1 U323 ( .A(\mem<55><2> ), .Y(n3644) );
  INVX1 U324 ( .A(\mem<55><3> ), .Y(n3643) );
  INVX1 U325 ( .A(\mem<55><4> ), .Y(n3642) );
  INVX1 U326 ( .A(\mem<55><5> ), .Y(n3641) );
  INVX1 U327 ( .A(\mem<55><6> ), .Y(n3640) );
  INVX1 U328 ( .A(\mem<55><7> ), .Y(n3639) );
  INVX1 U329 ( .A(\mem<54><0> ), .Y(n3638) );
  INVX1 U330 ( .A(\mem<54><1> ), .Y(n3637) );
  INVX1 U331 ( .A(\mem<54><2> ), .Y(n3636) );
  INVX1 U332 ( .A(\mem<54><3> ), .Y(n3635) );
  INVX1 U333 ( .A(\mem<54><4> ), .Y(n3634) );
  INVX1 U334 ( .A(\mem<54><5> ), .Y(n3633) );
  INVX1 U335 ( .A(\mem<54><6> ), .Y(n3632) );
  INVX1 U336 ( .A(\mem<54><7> ), .Y(n3631) );
  INVX1 U337 ( .A(\mem<53><0> ), .Y(n3630) );
  INVX1 U338 ( .A(\mem<53><1> ), .Y(n3629) );
  INVX1 U339 ( .A(\mem<53><2> ), .Y(n3628) );
  INVX1 U340 ( .A(\mem<53><3> ), .Y(n3627) );
  INVX1 U341 ( .A(\mem<53><4> ), .Y(n3626) );
  INVX1 U342 ( .A(\mem<53><5> ), .Y(n3625) );
  INVX1 U343 ( .A(\mem<53><6> ), .Y(n3624) );
  INVX1 U344 ( .A(\mem<53><7> ), .Y(n3623) );
  INVX1 U345 ( .A(\mem<52><0> ), .Y(n3622) );
  INVX1 U346 ( .A(\mem<52><1> ), .Y(n3621) );
  INVX1 U347 ( .A(\mem<52><2> ), .Y(n3620) );
  INVX1 U348 ( .A(\mem<52><3> ), .Y(n3619) );
  INVX1 U349 ( .A(\mem<52><4> ), .Y(n3618) );
  INVX1 U350 ( .A(\mem<52><5> ), .Y(n3617) );
  INVX1 U351 ( .A(\mem<52><6> ), .Y(n3616) );
  INVX1 U352 ( .A(\mem<52><7> ), .Y(n3615) );
  INVX1 U353 ( .A(\mem<51><0> ), .Y(n3614) );
  INVX1 U354 ( .A(\mem<51><1> ), .Y(n3613) );
  INVX1 U355 ( .A(\mem<51><2> ), .Y(n3612) );
  INVX1 U356 ( .A(\mem<51><3> ), .Y(n3611) );
  INVX1 U357 ( .A(\mem<51><4> ), .Y(n3610) );
  INVX1 U358 ( .A(\mem<51><5> ), .Y(n3609) );
  INVX1 U359 ( .A(\mem<51><6> ), .Y(n3608) );
  INVX1 U360 ( .A(\mem<51><7> ), .Y(n3607) );
  INVX1 U361 ( .A(\mem<50><0> ), .Y(n3606) );
  INVX1 U362 ( .A(\mem<50><1> ), .Y(n3605) );
  INVX1 U363 ( .A(\mem<50><2> ), .Y(n3604) );
  INVX1 U364 ( .A(\mem<50><3> ), .Y(n3603) );
  INVX1 U365 ( .A(\mem<50><4> ), .Y(n3602) );
  INVX1 U366 ( .A(\mem<50><5> ), .Y(n3601) );
  INVX1 U367 ( .A(\mem<50><6> ), .Y(n3600) );
  INVX1 U368 ( .A(\mem<50><7> ), .Y(n3599) );
  INVX1 U369 ( .A(\mem<49><0> ), .Y(n3598) );
  INVX1 U370 ( .A(\mem<49><1> ), .Y(n3597) );
  INVX1 U371 ( .A(\mem<49><2> ), .Y(n3596) );
  INVX1 U372 ( .A(\mem<49><3> ), .Y(n3595) );
  INVX1 U373 ( .A(\mem<49><4> ), .Y(n3594) );
  INVX1 U374 ( .A(\mem<49><5> ), .Y(n3593) );
  INVX1 U375 ( .A(\mem<49><6> ), .Y(n3592) );
  INVX1 U376 ( .A(\mem<49><7> ), .Y(n3591) );
  INVX1 U377 ( .A(\mem<48><0> ), .Y(n3590) );
  INVX1 U378 ( .A(\mem<48><1> ), .Y(n3589) );
  INVX1 U379 ( .A(\mem<48><2> ), .Y(n3588) );
  INVX1 U380 ( .A(\mem<48><3> ), .Y(n3587) );
  INVX1 U381 ( .A(\mem<48><4> ), .Y(n3586) );
  INVX1 U382 ( .A(\mem<48><5> ), .Y(n3585) );
  INVX1 U383 ( .A(\mem<48><6> ), .Y(n3584) );
  INVX1 U384 ( .A(\mem<48><7> ), .Y(n3583) );
  INVX1 U385 ( .A(\mem<47><0> ), .Y(n3582) );
  INVX1 U386 ( .A(\mem<47><1> ), .Y(n3581) );
  INVX1 U387 ( .A(\mem<47><2> ), .Y(n3580) );
  INVX1 U388 ( .A(\mem<47><3> ), .Y(n3579) );
  INVX1 U389 ( .A(\mem<47><4> ), .Y(n3578) );
  INVX1 U390 ( .A(\mem<47><5> ), .Y(n3577) );
  INVX1 U391 ( .A(\mem<47><6> ), .Y(n3576) );
  INVX1 U392 ( .A(\mem<47><7> ), .Y(n3575) );
  INVX1 U393 ( .A(\mem<46><0> ), .Y(n3574) );
  INVX1 U394 ( .A(\mem<46><1> ), .Y(n3573) );
  INVX1 U395 ( .A(\mem<46><2> ), .Y(n3572) );
  INVX1 U396 ( .A(\mem<46><3> ), .Y(n3571) );
  INVX1 U397 ( .A(\mem<46><4> ), .Y(n3570) );
  INVX1 U398 ( .A(\mem<46><5> ), .Y(n3569) );
  INVX1 U399 ( .A(\mem<46><6> ), .Y(n3568) );
  INVX1 U400 ( .A(\mem<46><7> ), .Y(n3567) );
  INVX1 U401 ( .A(\mem<45><0> ), .Y(n3566) );
  INVX1 U402 ( .A(\mem<45><1> ), .Y(n3565) );
  INVX1 U403 ( .A(\mem<45><2> ), .Y(n3564) );
  INVX1 U404 ( .A(\mem<45><3> ), .Y(n3563) );
  INVX1 U405 ( .A(\mem<45><4> ), .Y(n3562) );
  INVX1 U406 ( .A(\mem<45><5> ), .Y(n3561) );
  INVX1 U407 ( .A(\mem<45><6> ), .Y(n3560) );
  INVX1 U408 ( .A(\mem<45><7> ), .Y(n3559) );
  INVX1 U409 ( .A(\mem<44><0> ), .Y(n3558) );
  INVX1 U410 ( .A(\mem<44><1> ), .Y(n3557) );
  INVX1 U411 ( .A(\mem<44><2> ), .Y(n3556) );
  INVX1 U412 ( .A(\mem<44><3> ), .Y(n3555) );
  INVX1 U413 ( .A(\mem<44><4> ), .Y(n3554) );
  INVX1 U414 ( .A(\mem<44><5> ), .Y(n3553) );
  INVX1 U415 ( .A(\mem<44><6> ), .Y(n3552) );
  INVX1 U416 ( .A(\mem<44><7> ), .Y(n3551) );
  INVX1 U417 ( .A(\mem<43><0> ), .Y(n3550) );
  INVX1 U418 ( .A(\mem<43><1> ), .Y(n3549) );
  INVX1 U419 ( .A(\mem<43><2> ), .Y(n3548) );
  INVX1 U420 ( .A(\mem<43><3> ), .Y(n3547) );
  INVX1 U421 ( .A(\mem<43><4> ), .Y(n3546) );
  INVX1 U422 ( .A(\mem<43><5> ), .Y(n3545) );
  INVX1 U423 ( .A(\mem<43><6> ), .Y(n3544) );
  INVX1 U424 ( .A(\mem<43><7> ), .Y(n3543) );
  INVX1 U425 ( .A(\mem<42><0> ), .Y(n3542) );
  INVX1 U426 ( .A(\mem<42><1> ), .Y(n3541) );
  INVX1 U427 ( .A(\mem<42><2> ), .Y(n3540) );
  INVX1 U428 ( .A(\mem<42><3> ), .Y(n3539) );
  INVX1 U429 ( .A(\mem<42><4> ), .Y(n3538) );
  INVX1 U430 ( .A(\mem<42><5> ), .Y(n3537) );
  INVX1 U431 ( .A(\mem<42><6> ), .Y(n3536) );
  INVX1 U432 ( .A(\mem<42><7> ), .Y(n3535) );
  INVX1 U433 ( .A(\mem<41><0> ), .Y(n3534) );
  INVX1 U434 ( .A(\mem<41><1> ), .Y(n3533) );
  INVX1 U435 ( .A(\mem<41><2> ), .Y(n3532) );
  INVX1 U436 ( .A(\mem<41><3> ), .Y(n3531) );
  INVX1 U437 ( .A(\mem<41><4> ), .Y(n3530) );
  INVX1 U438 ( .A(\mem<41><5> ), .Y(n3529) );
  INVX1 U439 ( .A(\mem<41><6> ), .Y(n3528) );
  INVX1 U440 ( .A(\mem<41><7> ), .Y(n3527) );
  INVX1 U441 ( .A(\mem<40><0> ), .Y(n3526) );
  INVX1 U442 ( .A(\mem<40><1> ), .Y(n3525) );
  INVX1 U443 ( .A(\mem<40><2> ), .Y(n3524) );
  INVX1 U444 ( .A(\mem<40><3> ), .Y(n3523) );
  INVX1 U445 ( .A(\mem<40><4> ), .Y(n3522) );
  INVX1 U446 ( .A(\mem<40><5> ), .Y(n3521) );
  INVX1 U447 ( .A(\mem<40><6> ), .Y(n3520) );
  INVX1 U448 ( .A(\mem<40><7> ), .Y(n3519) );
  INVX1 U449 ( .A(\mem<39><0> ), .Y(n3518) );
  INVX1 U450 ( .A(\mem<39><1> ), .Y(n3517) );
  INVX1 U451 ( .A(\mem<39><2> ), .Y(n3516) );
  INVX1 U452 ( .A(\mem<39><3> ), .Y(n3515) );
  INVX1 U453 ( .A(\mem<39><4> ), .Y(n3514) );
  INVX1 U454 ( .A(\mem<39><5> ), .Y(n3513) );
  INVX1 U455 ( .A(\mem<39><6> ), .Y(n3512) );
  INVX1 U456 ( .A(\mem<39><7> ), .Y(n3511) );
  INVX1 U457 ( .A(\mem<38><0> ), .Y(n3510) );
  INVX1 U458 ( .A(\mem<38><1> ), .Y(n3509) );
  INVX1 U459 ( .A(\mem<38><2> ), .Y(n3508) );
  INVX1 U460 ( .A(\mem<38><3> ), .Y(n3507) );
  INVX1 U461 ( .A(\mem<38><4> ), .Y(n3506) );
  INVX1 U462 ( .A(\mem<38><5> ), .Y(n3505) );
  INVX1 U463 ( .A(\mem<38><6> ), .Y(n3504) );
  INVX1 U464 ( .A(\mem<38><7> ), .Y(n3503) );
  INVX1 U465 ( .A(\mem<37><0> ), .Y(n3502) );
  INVX1 U466 ( .A(\mem<37><1> ), .Y(n3501) );
  INVX1 U467 ( .A(\mem<37><2> ), .Y(n3500) );
  INVX1 U468 ( .A(\mem<37><3> ), .Y(n3499) );
  INVX1 U469 ( .A(\mem<37><4> ), .Y(n3498) );
  INVX1 U470 ( .A(\mem<37><5> ), .Y(n3497) );
  INVX1 U471 ( .A(\mem<37><6> ), .Y(n3496) );
  INVX1 U472 ( .A(\mem<37><7> ), .Y(n3495) );
  INVX1 U473 ( .A(\mem<36><0> ), .Y(n3494) );
  INVX1 U474 ( .A(\mem<36><1> ), .Y(n3493) );
  INVX1 U475 ( .A(\mem<36><2> ), .Y(n3492) );
  INVX1 U476 ( .A(\mem<36><3> ), .Y(n3491) );
  INVX1 U477 ( .A(\mem<36><4> ), .Y(n3490) );
  INVX1 U478 ( .A(\mem<36><5> ), .Y(n3489) );
  INVX1 U479 ( .A(\mem<36><6> ), .Y(n3488) );
  INVX1 U480 ( .A(\mem<36><7> ), .Y(n3487) );
  INVX1 U481 ( .A(\mem<35><0> ), .Y(n3486) );
  INVX1 U482 ( .A(\mem<35><1> ), .Y(n3485) );
  INVX1 U483 ( .A(\mem<35><2> ), .Y(n3484) );
  INVX1 U484 ( .A(\mem<35><3> ), .Y(n3483) );
  INVX1 U485 ( .A(\mem<35><4> ), .Y(n3482) );
  INVX1 U486 ( .A(\mem<35><5> ), .Y(n3481) );
  INVX1 U487 ( .A(\mem<35><6> ), .Y(n3480) );
  INVX1 U488 ( .A(\mem<35><7> ), .Y(n3479) );
  INVX1 U489 ( .A(\mem<34><0> ), .Y(n3478) );
  INVX1 U490 ( .A(\mem<34><1> ), .Y(n3477) );
  INVX1 U491 ( .A(\mem<34><2> ), .Y(n3476) );
  INVX1 U492 ( .A(\mem<34><3> ), .Y(n3475) );
  INVX1 U493 ( .A(\mem<34><4> ), .Y(n3474) );
  INVX1 U494 ( .A(\mem<34><5> ), .Y(n3473) );
  INVX1 U495 ( .A(\mem<34><6> ), .Y(n3472) );
  INVX1 U496 ( .A(\mem<34><7> ), .Y(n3471) );
  INVX1 U497 ( .A(\mem<33><0> ), .Y(n3470) );
  INVX1 U498 ( .A(\mem<33><1> ), .Y(n3469) );
  INVX1 U499 ( .A(\mem<33><2> ), .Y(n3468) );
  INVX1 U500 ( .A(\mem<33><3> ), .Y(n3467) );
  INVX1 U501 ( .A(\mem<33><4> ), .Y(n3466) );
  INVX1 U502 ( .A(\mem<33><5> ), .Y(n3465) );
  INVX1 U503 ( .A(\mem<33><6> ), .Y(n3464) );
  INVX1 U504 ( .A(\mem<33><7> ), .Y(n3463) );
  INVX1 U505 ( .A(\mem<32><0> ), .Y(n3462) );
  INVX1 U506 ( .A(\mem<32><1> ), .Y(n3461) );
  INVX1 U507 ( .A(\mem<32><2> ), .Y(n3460) );
  INVX1 U508 ( .A(\mem<32><3> ), .Y(n3459) );
  INVX1 U509 ( .A(\mem<32><4> ), .Y(n3458) );
  INVX1 U510 ( .A(\mem<32><5> ), .Y(n3457) );
  INVX1 U511 ( .A(\mem<32><6> ), .Y(n3456) );
  INVX1 U512 ( .A(\mem<32><7> ), .Y(n3455) );
  INVX1 U513 ( .A(\mem<31><0> ), .Y(n3454) );
  INVX1 U514 ( .A(\mem<31><1> ), .Y(n3453) );
  INVX1 U515 ( .A(\mem<31><2> ), .Y(n3452) );
  INVX1 U516 ( .A(\mem<31><3> ), .Y(n3451) );
  INVX1 U517 ( .A(\mem<31><4> ), .Y(n3450) );
  INVX1 U518 ( .A(\mem<31><5> ), .Y(n3449) );
  INVX1 U519 ( .A(\mem<31><6> ), .Y(n3448) );
  INVX1 U520 ( .A(\mem<31><7> ), .Y(n3447) );
  INVX1 U521 ( .A(\mem<30><0> ), .Y(n3446) );
  INVX1 U522 ( .A(\mem<30><1> ), .Y(n3445) );
  INVX1 U523 ( .A(\mem<30><2> ), .Y(n3444) );
  INVX1 U524 ( .A(\mem<30><3> ), .Y(n3443) );
  INVX1 U525 ( .A(\mem<30><4> ), .Y(n3442) );
  INVX1 U526 ( .A(\mem<30><5> ), .Y(n3441) );
  INVX1 U527 ( .A(\mem<30><6> ), .Y(n3440) );
  INVX1 U528 ( .A(\mem<30><7> ), .Y(n3439) );
  INVX1 U529 ( .A(\mem<29><0> ), .Y(n3438) );
  INVX1 U530 ( .A(\mem<29><1> ), .Y(n3437) );
  INVX1 U531 ( .A(\mem<29><2> ), .Y(n3436) );
  INVX1 U532 ( .A(\mem<29><3> ), .Y(n3435) );
  INVX1 U533 ( .A(\mem<29><4> ), .Y(n3434) );
  INVX1 U534 ( .A(\mem<29><5> ), .Y(n3433) );
  INVX1 U535 ( .A(\mem<29><6> ), .Y(n3432) );
  INVX1 U536 ( .A(\mem<29><7> ), .Y(n3431) );
  INVX1 U537 ( .A(\mem<28><0> ), .Y(n3430) );
  INVX1 U538 ( .A(\mem<28><1> ), .Y(n3429) );
  INVX1 U539 ( .A(\mem<28><2> ), .Y(n3428) );
  INVX1 U540 ( .A(\mem<28><3> ), .Y(n3427) );
  INVX1 U541 ( .A(\mem<28><4> ), .Y(n3426) );
  INVX1 U542 ( .A(\mem<28><5> ), .Y(n3425) );
  INVX1 U543 ( .A(\mem<28><6> ), .Y(n3424) );
  INVX1 U544 ( .A(\mem<28><7> ), .Y(n3423) );
  INVX1 U545 ( .A(\mem<27><0> ), .Y(n3422) );
  INVX1 U546 ( .A(\mem<27><1> ), .Y(n3421) );
  INVX1 U547 ( .A(\mem<27><2> ), .Y(n3420) );
  INVX1 U548 ( .A(\mem<27><3> ), .Y(n3419) );
  INVX1 U549 ( .A(\mem<27><4> ), .Y(n3418) );
  INVX1 U550 ( .A(\mem<27><5> ), .Y(n3417) );
  INVX1 U551 ( .A(\mem<27><6> ), .Y(n3416) );
  INVX1 U552 ( .A(\mem<27><7> ), .Y(n3415) );
  INVX1 U553 ( .A(\mem<26><0> ), .Y(n3414) );
  INVX1 U554 ( .A(\mem<26><1> ), .Y(n3413) );
  INVX1 U555 ( .A(\mem<26><2> ), .Y(n3412) );
  INVX1 U556 ( .A(\mem<26><3> ), .Y(n3411) );
  INVX1 U557 ( .A(\mem<26><4> ), .Y(n3410) );
  INVX1 U558 ( .A(\mem<26><5> ), .Y(n3409) );
  INVX1 U559 ( .A(\mem<26><6> ), .Y(n3408) );
  INVX1 U560 ( .A(\mem<26><7> ), .Y(n3407) );
  INVX1 U561 ( .A(\mem<25><0> ), .Y(n3406) );
  INVX1 U562 ( .A(\mem<25><1> ), .Y(n3405) );
  INVX1 U563 ( .A(\mem<25><2> ), .Y(n3404) );
  INVX1 U564 ( .A(\mem<25><3> ), .Y(n3403) );
  INVX1 U565 ( .A(\mem<25><4> ), .Y(n3402) );
  INVX1 U566 ( .A(\mem<25><5> ), .Y(n3401) );
  INVX1 U567 ( .A(\mem<25><6> ), .Y(n3400) );
  INVX1 U568 ( .A(\mem<25><7> ), .Y(n3399) );
  INVX1 U569 ( .A(\mem<24><0> ), .Y(n3398) );
  INVX1 U570 ( .A(\mem<24><1> ), .Y(n3397) );
  INVX1 U571 ( .A(\mem<24><2> ), .Y(n3396) );
  INVX1 U572 ( .A(\mem<24><3> ), .Y(n3395) );
  INVX1 U573 ( .A(\mem<24><4> ), .Y(n3394) );
  INVX1 U574 ( .A(\mem<24><5> ), .Y(n3393) );
  INVX1 U575 ( .A(\mem<24><6> ), .Y(n3392) );
  INVX1 U576 ( .A(\mem<24><7> ), .Y(n3391) );
  INVX1 U577 ( .A(\mem<23><0> ), .Y(n3390) );
  INVX1 U578 ( .A(\mem<23><1> ), .Y(n3389) );
  INVX1 U579 ( .A(\mem<23><2> ), .Y(n3388) );
  INVX1 U580 ( .A(\mem<23><3> ), .Y(n3387) );
  INVX1 U581 ( .A(\mem<23><4> ), .Y(n3386) );
  INVX1 U582 ( .A(\mem<23><5> ), .Y(n3385) );
  INVX1 U583 ( .A(\mem<23><6> ), .Y(n3384) );
  INVX1 U584 ( .A(\mem<23><7> ), .Y(n3383) );
  INVX1 U585 ( .A(\mem<22><0> ), .Y(n3382) );
  INVX1 U586 ( .A(\mem<22><1> ), .Y(n3381) );
  INVX1 U587 ( .A(\mem<22><2> ), .Y(n3380) );
  INVX1 U588 ( .A(\mem<22><3> ), .Y(n3379) );
  INVX1 U589 ( .A(\mem<22><4> ), .Y(n3378) );
  INVX1 U590 ( .A(\mem<22><5> ), .Y(n3377) );
  INVX1 U591 ( .A(\mem<22><6> ), .Y(n3376) );
  INVX1 U592 ( .A(\mem<22><7> ), .Y(n3375) );
  INVX1 U593 ( .A(\mem<21><0> ), .Y(n3374) );
  INVX1 U594 ( .A(\mem<21><1> ), .Y(n3373) );
  INVX1 U595 ( .A(\mem<21><2> ), .Y(n3372) );
  INVX1 U596 ( .A(\mem<21><3> ), .Y(n3371) );
  INVX1 U597 ( .A(\mem<21><4> ), .Y(n3370) );
  INVX1 U598 ( .A(\mem<21><5> ), .Y(n3369) );
  INVX1 U599 ( .A(\mem<21><6> ), .Y(n3368) );
  INVX1 U600 ( .A(\mem<21><7> ), .Y(n3367) );
  INVX1 U601 ( .A(\mem<20><0> ), .Y(n3366) );
  INVX1 U602 ( .A(\mem<20><1> ), .Y(n3365) );
  INVX1 U603 ( .A(\mem<20><2> ), .Y(n3364) );
  INVX1 U604 ( .A(\mem<20><3> ), .Y(n3363) );
  INVX1 U605 ( .A(\mem<20><4> ), .Y(n3362) );
  INVX1 U606 ( .A(\mem<20><5> ), .Y(n3361) );
  INVX1 U607 ( .A(\mem<20><6> ), .Y(n3360) );
  INVX1 U608 ( .A(\mem<20><7> ), .Y(n3359) );
  INVX1 U609 ( .A(\mem<19><0> ), .Y(n3358) );
  INVX1 U610 ( .A(\mem<19><1> ), .Y(n3357) );
  INVX1 U611 ( .A(\mem<19><2> ), .Y(n3356) );
  INVX1 U612 ( .A(\mem<19><3> ), .Y(n3355) );
  INVX1 U613 ( .A(\mem<19><4> ), .Y(n3354) );
  INVX1 U614 ( .A(\mem<19><5> ), .Y(n3353) );
  INVX1 U615 ( .A(\mem<19><6> ), .Y(n3352) );
  INVX1 U616 ( .A(\mem<19><7> ), .Y(n3351) );
  INVX1 U617 ( .A(\mem<18><0> ), .Y(n3350) );
  INVX1 U618 ( .A(\mem<18><1> ), .Y(n3349) );
  INVX1 U619 ( .A(\mem<18><2> ), .Y(n3348) );
  INVX1 U620 ( .A(\mem<18><3> ), .Y(n3347) );
  INVX1 U621 ( .A(\mem<18><4> ), .Y(n3346) );
  INVX1 U622 ( .A(\mem<18><5> ), .Y(n3345) );
  INVX1 U623 ( .A(\mem<18><6> ), .Y(n3344) );
  INVX1 U624 ( .A(\mem<18><7> ), .Y(n3343) );
  INVX1 U625 ( .A(\mem<17><0> ), .Y(n3342) );
  INVX1 U626 ( .A(\mem<17><1> ), .Y(n3341) );
  INVX1 U627 ( .A(\mem<17><2> ), .Y(n3340) );
  INVX1 U628 ( .A(\mem<17><3> ), .Y(n3339) );
  INVX1 U629 ( .A(\mem<17><4> ), .Y(n3338) );
  INVX1 U630 ( .A(\mem<17><5> ), .Y(n3337) );
  INVX1 U631 ( .A(\mem<17><6> ), .Y(n3336) );
  INVX1 U632 ( .A(\mem<17><7> ), .Y(n3335) );
  INVX1 U633 ( .A(\mem<16><0> ), .Y(n3334) );
  INVX1 U634 ( .A(\mem<16><1> ), .Y(n3333) );
  INVX1 U635 ( .A(\mem<16><2> ), .Y(n3332) );
  INVX1 U636 ( .A(\mem<16><3> ), .Y(n3331) );
  INVX1 U637 ( .A(\mem<16><4> ), .Y(n3330) );
  INVX1 U638 ( .A(\mem<16><5> ), .Y(n3329) );
  INVX1 U639 ( .A(\mem<16><6> ), .Y(n3328) );
  INVX1 U640 ( .A(\mem<16><7> ), .Y(n3327) );
  INVX1 U641 ( .A(\mem<15><0> ), .Y(n3326) );
  INVX1 U642 ( .A(\mem<15><1> ), .Y(n3325) );
  INVX1 U643 ( .A(\mem<15><2> ), .Y(n3324) );
  INVX1 U644 ( .A(\mem<15><3> ), .Y(n3323) );
  INVX1 U645 ( .A(\mem<15><4> ), .Y(n3322) );
  INVX1 U646 ( .A(\mem<15><5> ), .Y(n3321) );
  INVX1 U647 ( .A(\mem<15><6> ), .Y(n3320) );
  INVX1 U648 ( .A(\mem<15><7> ), .Y(n3319) );
  INVX1 U649 ( .A(\mem<14><0> ), .Y(n3318) );
  INVX1 U650 ( .A(\mem<14><1> ), .Y(n3317) );
  INVX1 U651 ( .A(\mem<14><2> ), .Y(n3316) );
  INVX1 U652 ( .A(\mem<14><3> ), .Y(n3315) );
  INVX1 U653 ( .A(\mem<14><4> ), .Y(n3314) );
  INVX1 U654 ( .A(\mem<14><5> ), .Y(n3313) );
  INVX1 U655 ( .A(\mem<14><6> ), .Y(n3312) );
  INVX1 U656 ( .A(\mem<14><7> ), .Y(n3311) );
  INVX1 U657 ( .A(\mem<13><0> ), .Y(n3310) );
  INVX1 U658 ( .A(\mem<13><1> ), .Y(n3309) );
  INVX1 U659 ( .A(\mem<13><2> ), .Y(n3308) );
  INVX1 U660 ( .A(\mem<13><3> ), .Y(n3307) );
  INVX1 U661 ( .A(\mem<13><4> ), .Y(n3306) );
  INVX1 U662 ( .A(\mem<13><5> ), .Y(n3305) );
  INVX1 U663 ( .A(\mem<13><6> ), .Y(n3304) );
  INVX1 U664 ( .A(\mem<13><7> ), .Y(n3303) );
  INVX1 U665 ( .A(\mem<12><0> ), .Y(n3302) );
  INVX1 U666 ( .A(\mem<12><1> ), .Y(n3301) );
  INVX1 U667 ( .A(\mem<12><2> ), .Y(n3300) );
  INVX1 U668 ( .A(\mem<12><3> ), .Y(n3299) );
  INVX1 U669 ( .A(\mem<12><4> ), .Y(n3298) );
  INVX1 U670 ( .A(\mem<12><5> ), .Y(n3297) );
  INVX1 U671 ( .A(\mem<12><6> ), .Y(n3296) );
  INVX1 U672 ( .A(\mem<12><7> ), .Y(n3295) );
  INVX1 U673 ( .A(\mem<11><0> ), .Y(n3294) );
  INVX1 U674 ( .A(\mem<11><1> ), .Y(n3293) );
  INVX1 U675 ( .A(\mem<11><2> ), .Y(n3292) );
  INVX1 U676 ( .A(\mem<11><3> ), .Y(n3291) );
  INVX1 U677 ( .A(\mem<11><4> ), .Y(n3290) );
  INVX1 U678 ( .A(\mem<11><5> ), .Y(n3289) );
  INVX1 U679 ( .A(\mem<11><6> ), .Y(n3288) );
  INVX1 U680 ( .A(\mem<11><7> ), .Y(n3287) );
  INVX1 U681 ( .A(\mem<10><0> ), .Y(n3286) );
  INVX1 U682 ( .A(\mem<10><1> ), .Y(n3285) );
  INVX1 U683 ( .A(\mem<10><2> ), .Y(n3284) );
  INVX1 U684 ( .A(\mem<10><3> ), .Y(n3283) );
  INVX1 U685 ( .A(\mem<10><4> ), .Y(n3282) );
  INVX1 U686 ( .A(\mem<10><5> ), .Y(n3281) );
  INVX1 U687 ( .A(\mem<10><6> ), .Y(n3280) );
  INVX1 U688 ( .A(\mem<10><7> ), .Y(n3279) );
  INVX1 U689 ( .A(\mem<9><0> ), .Y(n3278) );
  INVX1 U690 ( .A(\mem<9><1> ), .Y(n3277) );
  INVX1 U691 ( .A(\mem<9><2> ), .Y(n3276) );
  INVX1 U692 ( .A(\mem<9><3> ), .Y(n3275) );
  INVX1 U693 ( .A(\mem<9><4> ), .Y(n3274) );
  INVX1 U694 ( .A(\mem<9><5> ), .Y(n3273) );
  INVX1 U695 ( .A(\mem<9><6> ), .Y(n3272) );
  INVX1 U696 ( .A(\mem<9><7> ), .Y(n3271) );
  INVX1 U697 ( .A(\mem<8><0> ), .Y(n3270) );
  INVX1 U698 ( .A(\mem<8><1> ), .Y(n3269) );
  INVX1 U699 ( .A(\mem<8><2> ), .Y(n3268) );
  INVX1 U700 ( .A(\mem<8><3> ), .Y(n3267) );
  INVX1 U701 ( .A(\mem<8><4> ), .Y(n3266) );
  INVX1 U702 ( .A(\mem<8><5> ), .Y(n3265) );
  INVX1 U703 ( .A(\mem<8><6> ), .Y(n3264) );
  INVX1 U704 ( .A(\mem<8><7> ), .Y(n3263) );
  INVX1 U705 ( .A(\mem<7><0> ), .Y(n3262) );
  INVX1 U706 ( .A(\mem<7><1> ), .Y(n3261) );
  INVX1 U707 ( .A(\mem<7><2> ), .Y(n3260) );
  INVX1 U708 ( .A(\mem<7><3> ), .Y(n3259) );
  INVX1 U709 ( .A(\mem<7><4> ), .Y(n3258) );
  INVX1 U710 ( .A(\mem<7><5> ), .Y(n3257) );
  INVX1 U711 ( .A(\mem<7><6> ), .Y(n3256) );
  INVX1 U712 ( .A(\mem<7><7> ), .Y(n3255) );
  INVX1 U713 ( .A(\mem<6><0> ), .Y(n3254) );
  INVX1 U714 ( .A(\mem<6><1> ), .Y(n3253) );
  INVX1 U715 ( .A(\mem<6><2> ), .Y(n3252) );
  INVX1 U716 ( .A(\mem<6><3> ), .Y(n3251) );
  INVX1 U717 ( .A(\mem<6><4> ), .Y(n3250) );
  INVX1 U718 ( .A(\mem<6><5> ), .Y(n3249) );
  INVX1 U719 ( .A(\mem<6><6> ), .Y(n3248) );
  INVX1 U720 ( .A(\mem<6><7> ), .Y(n3247) );
  INVX1 U721 ( .A(\mem<5><0> ), .Y(n3246) );
  INVX1 U722 ( .A(\mem<5><1> ), .Y(n3245) );
  INVX1 U723 ( .A(\mem<5><2> ), .Y(n3244) );
  INVX1 U724 ( .A(\mem<5><3> ), .Y(n3243) );
  INVX1 U725 ( .A(\mem<5><4> ), .Y(n3242) );
  INVX1 U726 ( .A(\mem<5><5> ), .Y(n3241) );
  INVX1 U727 ( .A(\mem<5><6> ), .Y(n3240) );
  INVX1 U728 ( .A(\mem<5><7> ), .Y(n3239) );
  INVX1 U729 ( .A(\mem<4><0> ), .Y(n3238) );
  INVX1 U730 ( .A(\mem<4><1> ), .Y(n3237) );
  INVX1 U731 ( .A(\mem<4><2> ), .Y(n3236) );
  INVX1 U732 ( .A(\mem<4><3> ), .Y(n3235) );
  INVX1 U733 ( .A(\mem<4><4> ), .Y(n3234) );
  INVX1 U734 ( .A(\mem<4><5> ), .Y(n3233) );
  INVX1 U735 ( .A(\mem<4><6> ), .Y(n3232) );
  INVX1 U736 ( .A(\mem<4><7> ), .Y(n3231) );
  INVX1 U737 ( .A(\mem<3><0> ), .Y(n3230) );
  INVX1 U738 ( .A(\mem<3><1> ), .Y(n3229) );
  INVX1 U739 ( .A(\mem<3><2> ), .Y(n3228) );
  INVX1 U740 ( .A(\mem<3><3> ), .Y(n3227) );
  INVX1 U741 ( .A(\mem<3><4> ), .Y(n3226) );
  INVX1 U742 ( .A(\mem<3><5> ), .Y(n3225) );
  INVX1 U743 ( .A(\mem<3><6> ), .Y(n3224) );
  INVX1 U744 ( .A(\mem<3><7> ), .Y(n3223) );
  INVX1 U745 ( .A(\mem<2><0> ), .Y(n3222) );
  INVX1 U746 ( .A(\mem<2><1> ), .Y(n3221) );
  INVX1 U747 ( .A(\mem<2><2> ), .Y(n3220) );
  INVX1 U748 ( .A(\mem<2><3> ), .Y(n3219) );
  INVX1 U749 ( .A(\mem<2><4> ), .Y(n3218) );
  INVX1 U750 ( .A(\mem<2><5> ), .Y(n3217) );
  INVX1 U751 ( .A(\mem<2><6> ), .Y(n3216) );
  INVX1 U752 ( .A(\mem<2><7> ), .Y(n3215) );
  INVX1 U753 ( .A(\mem<1><0> ), .Y(n3214) );
  INVX1 U754 ( .A(\mem<1><1> ), .Y(n3213) );
  INVX1 U755 ( .A(\mem<1><2> ), .Y(n3212) );
  INVX1 U756 ( .A(\mem<1><3> ), .Y(n3211) );
  INVX1 U757 ( .A(\mem<1><4> ), .Y(n3210) );
  INVX1 U758 ( .A(\mem<1><5> ), .Y(n3209) );
  INVX1 U759 ( .A(\mem<1><6> ), .Y(n3208) );
  INVX1 U760 ( .A(\mem<1><7> ), .Y(n3207) );
  INVX1 U761 ( .A(\mem<0><0> ), .Y(n3206) );
  INVX1 U762 ( .A(\mem<0><1> ), .Y(n3205) );
  INVX1 U763 ( .A(\mem<0><2> ), .Y(n3204) );
  INVX1 U764 ( .A(\mem<0><3> ), .Y(n3203) );
  INVX1 U765 ( .A(\mem<0><4> ), .Y(n3202) );
  INVX1 U766 ( .A(\mem<0><5> ), .Y(n3201) );
  INVX1 U767 ( .A(\mem<0><6> ), .Y(n3200) );
  INVX1 U768 ( .A(\mem<0><7> ), .Y(n3199) );
  INVX1 U769 ( .A(n3113), .Y(n3091) );
  INVX1 U770 ( .A(n3113), .Y(n3093) );
  INVX1 U771 ( .A(n3113), .Y(n3092) );
  INVX1 U772 ( .A(n3113), .Y(n3094) );
  INVX1 U773 ( .A(n3184), .Y(n3099) );
  INVX1 U774 ( .A(n3184), .Y(n3097) );
  INVX1 U775 ( .A(n3186), .Y(n3088) );
  INVX1 U776 ( .A(n3186), .Y(n3087) );
  INVX1 U777 ( .A(n3186), .Y(n3089) );
  INVX1 U778 ( .A(n3184), .Y(n3095) );
  INVX1 U779 ( .A(n3184), .Y(n3096) );
  INVX1 U780 ( .A(n3079), .Y(n3083) );
  INVX1 U781 ( .A(n3079), .Y(n3082) );
  INVX1 U782 ( .A(n3186), .Y(n3084) );
  INVX1 U783 ( .A(n3186), .Y(n3090) );
  INVX1 U784 ( .A(n3091), .Y(n3100) );
  INVX1 U785 ( .A(n3093), .Y(n3101) );
  INVX1 U786 ( .A(n3092), .Y(n3098) );
  INVX1 U787 ( .A(N178), .Y(n3186) );
  INVX1 U788 ( .A(n3186), .Y(n3085) );
  INVX1 U789 ( .A(n3186), .Y(n3086) );
  OR2X1 U790 ( .A(n2407), .B(n210), .Y(n181) );
  OR2X1 U791 ( .A(n2413), .B(n213), .Y(n182) );
  OR2X1 U792 ( .A(n2419), .B(n216), .Y(n183) );
  OR2X1 U793 ( .A(n2425), .B(n219), .Y(n184) );
  OR2X1 U794 ( .A(n2431), .B(n222), .Y(n185) );
  OR2X1 U795 ( .A(n2437), .B(n225), .Y(n186) );
  OR2X1 U796 ( .A(n2443), .B(n228), .Y(n187) );
  OR2X1 U797 ( .A(n2449), .B(n231), .Y(n188) );
  INVX1 U798 ( .A(N180), .Y(n3187) );
  INVX1 U799 ( .A(N177), .Y(n3184) );
  OR2X1 U800 ( .A(n2356), .B(n192), .Y(n165) );
  OR2X1 U801 ( .A(n2359), .B(n193), .Y(n166) );
  OR2X1 U802 ( .A(n2362), .B(n194), .Y(n167) );
  OR2X1 U803 ( .A(n2365), .B(n195), .Y(n168) );
  OR2X1 U804 ( .A(n2368), .B(n196), .Y(n169) );
  OR2X1 U805 ( .A(n2371), .B(n197), .Y(n170) );
  OR2X1 U806 ( .A(n2374), .B(n198), .Y(n171) );
  OR2X1 U807 ( .A(n2377), .B(n199), .Y(n172) );
  OR2X1 U808 ( .A(n2380), .B(n200), .Y(n173) );
  OR2X1 U809 ( .A(n2383), .B(n201), .Y(n174) );
  OR2X1 U810 ( .A(n2386), .B(n202), .Y(n175) );
  OR2X1 U811 ( .A(n2389), .B(n203), .Y(n176) );
  OR2X1 U812 ( .A(n2392), .B(n204), .Y(n177) );
  OR2X1 U813 ( .A(n2395), .B(n205), .Y(n178) );
  OR2X1 U814 ( .A(n2398), .B(n206), .Y(n179) );
  OR2X1 U815 ( .A(n2401), .B(n207), .Y(n180) );
  OR2X1 U816 ( .A(n189), .B(n3187), .Y(n190) );
  OR2X1 U1889 ( .A(n10), .B(n7), .Y(n6) );
  OR2X1 U1891 ( .A(n20), .B(n17), .Y(n16) );
  OR2X1 U1893 ( .A(n30), .B(n27), .Y(n26) );
  OR2X1 U1895 ( .A(n40), .B(n37), .Y(n36) );
  OR2X1 U1897 ( .A(n50), .B(n47), .Y(n46) );
  OR2X1 U1899 ( .A(n60), .B(n57), .Y(n56) );
  OR2X1 U1901 ( .A(n70), .B(n67), .Y(n66) );
  OR2X1 U1903 ( .A(n80), .B(n77), .Y(n76) );
  OR2X1 U1904 ( .A(n90), .B(n87), .Y(n86) );
  OR2X1 U1908 ( .A(n100), .B(n97), .Y(n96) );
  OR2X1 U1913 ( .A(n110), .B(n107), .Y(n106) );
  OR2X1 U1918 ( .A(n120), .B(n117), .Y(n116) );
  OR2X1 U1923 ( .A(n130), .B(n127), .Y(n126) );
  OR2X1 U1929 ( .A(n140), .B(n137), .Y(n136) );
  OR2X1 U1934 ( .A(n150), .B(n147), .Y(n146) );
  OR2X1 U1939 ( .A(n160), .B(n157), .Y(n156) );
  INVX1 U1944 ( .A(n3184), .Y(n3113) );
  INVX1 U1951 ( .A(n3186), .Y(n3185) );
  OR2X1 U1956 ( .A(n3), .B(n4), .Y(n2) );
  OR2X1 U1961 ( .A(n13), .B(n14), .Y(n12) );
  OR2X1 U1966 ( .A(n23), .B(n24), .Y(n22) );
  OR2X1 U1972 ( .A(n33), .B(n34), .Y(n32) );
  OR2X1 U1977 ( .A(n43), .B(n44), .Y(n42) );
  OR2X1 U1982 ( .A(n53), .B(n54), .Y(n52) );
  OR2X1 U1987 ( .A(n63), .B(n64), .Y(n62) );
  OR2X1 U1994 ( .A(n73), .B(n74), .Y(n72) );
  OR2X1 U1999 ( .A(n83), .B(n84), .Y(n82) );
  OR2X1 U2004 ( .A(n93), .B(n94), .Y(n92) );
  OR2X1 U2009 ( .A(n103), .B(n104), .Y(n102) );
  OR2X1 U2015 ( .A(n113), .B(n114), .Y(n112) );
  OR2X1 U2020 ( .A(n123), .B(n124), .Y(n122) );
  OR2X1 U2025 ( .A(n133), .B(n134), .Y(n132) );
  OR2X1 U2030 ( .A(n143), .B(n144), .Y(n142) );
  OR2X1 U2037 ( .A(n153), .B(n154), .Y(n152) );
  OR2X1 U2042 ( .A(n5), .B(n2), .Y(n1) );
  OR2X1 U2047 ( .A(n15), .B(n12), .Y(n11) );
  OR2X1 U2052 ( .A(n25), .B(n22), .Y(n21) );
  OR2X1 U2058 ( .A(n35), .B(n32), .Y(n31) );
  OR2X1 U2063 ( .A(n45), .B(n42), .Y(n41) );
  OR2X1 U2068 ( .A(n55), .B(n52), .Y(n51) );
  OR2X1 U2073 ( .A(n65), .B(n62), .Y(n61) );
  OR2X1 U2080 ( .A(n75), .B(n72), .Y(n71) );
  OR2X1 U2085 ( .A(n85), .B(n82), .Y(n81) );
  OR2X1 U2090 ( .A(n95), .B(n92), .Y(n91) );
  OR2X1 U2095 ( .A(n105), .B(n102), .Y(n101) );
  OR2X1 U2101 ( .A(n115), .B(n112), .Y(n111) );
  OR2X1 U2106 ( .A(n125), .B(n122), .Y(n121) );
  OR2X1 U2111 ( .A(n135), .B(n132), .Y(n131) );
  OR2X1 U2116 ( .A(n145), .B(n142), .Y(n141) );
  OR2X1 U2123 ( .A(n155), .B(n152), .Y(n151) );
  INVX1 U2128 ( .A(N179), .Y(n3079) );
  INVX1 U2133 ( .A(n3079), .Y(n3081) );
  INVX1 U2138 ( .A(n3079), .Y(n3080) );
  INVX1 U2144 ( .A(n3181), .Y(n3178) );
  INVX1 U2149 ( .A(n3182), .Y(n3179) );
  INVX1 U2154 ( .A(n1805), .Y(n3) );
  INVX1 U2159 ( .A(n1804), .Y(n4) );
  INVX1 U2166 ( .A(n1803), .Y(n5) );
  INVX1 U2171 ( .A(n1799), .Y(n8) );
  INVX1 U2176 ( .A(n1798), .Y(n9) );
  INVX1 U2181 ( .A(n1797), .Y(n10) );
  INVX1 U2187 ( .A(n1767), .Y(n13) );
  INVX1 U2192 ( .A(n1766), .Y(n14) );
  INVX1 U2197 ( .A(n1765), .Y(n15) );
  INVX1 U2202 ( .A(n1762), .Y(n18) );
  INVX1 U2208 ( .A(n1761), .Y(n19) );
  INVX1 U2210 ( .A(n1760), .Y(n20) );
  INVX1 U2212 ( .A(n1730), .Y(n23) );
  INVX1 U2213 ( .A(n1729), .Y(n24) );
  INVX1 U2215 ( .A(n1728), .Y(n25) );
  INVX1 U2216 ( .A(n1725), .Y(n28) );
  INVX1 U2218 ( .A(n1724), .Y(n29) );
  INVX1 U2219 ( .A(n1723), .Y(n30) );
  INVX1 U2221 ( .A(n1705), .Y(n33) );
  INVX1 U2222 ( .A(n1704), .Y(n34) );
  INVX1 U2223 ( .A(n1703), .Y(n35) );
  INVX1 U2225 ( .A(n1700), .Y(n38) );
  INVX1 U2226 ( .A(n1699), .Y(n39) );
  INVX1 U2228 ( .A(n1698), .Y(n40) );
  INVX1 U2229 ( .A(n1678), .Y(n43) );
  INVX1 U2231 ( .A(n1677), .Y(n44) );
  INVX1 U2232 ( .A(n1676), .Y(n45) );
  INVX1 U2234 ( .A(n1673), .Y(n48) );
  INVX1 U2236 ( .A(n1672), .Y(n49) );
  INVX1 U2237 ( .A(n1671), .Y(n50) );
  INVX1 U2238 ( .A(n1653), .Y(n53) );
  INVX1 U2240 ( .A(n1652), .Y(n54) );
  INVX1 U2241 ( .A(n1651), .Y(n55) );
  INVX1 U2243 ( .A(n1648), .Y(n58) );
  INVX1 U2244 ( .A(n1647), .Y(n59) );
  INVX1 U2246 ( .A(n1646), .Y(n60) );
  INVX1 U2247 ( .A(n1626), .Y(n63) );
  INVX1 U2249 ( .A(n1625), .Y(n64) );
  INVX1 U2250 ( .A(n1624), .Y(n65) );
  INVX1 U2251 ( .A(n1621), .Y(n68) );
  INVX1 U2253 ( .A(n1620), .Y(n69) );
  INVX1 U2254 ( .A(n1619), .Y(n70) );
  INVX1 U2256 ( .A(n1601), .Y(n73) );
  INVX1 U2257 ( .A(n1600), .Y(n74) );
  INVX1 U2259 ( .A(n1599), .Y(n75) );
  INVX1 U2260 ( .A(n1596), .Y(n78) );
  INVX1 U2262 ( .A(n1595), .Y(n79) );
  INVX1 U2264 ( .A(n1594), .Y(n80) );
  INVX1 U2265 ( .A(n1574), .Y(n83) );
  INVX1 U2267 ( .A(n1573), .Y(n84) );
  INVX1 U2269 ( .A(n1572), .Y(n85) );
  INVX1 U2271 ( .A(n1569), .Y(n88) );
  INVX1 U2272 ( .A(n1568), .Y(n89) );
  INVX1 U2274 ( .A(n1567), .Y(n90) );
  INVX1 U2275 ( .A(n1549), .Y(n93) );
  INVX1 U2277 ( .A(n1548), .Y(n94) );
  INVX1 U2278 ( .A(n1547), .Y(n95) );
  INVX1 U2286 ( .A(n1544), .Y(n98) );
  INVX1 U2287 ( .A(n1543), .Y(n99) );
  INVX1 U2289 ( .A(n1542), .Y(n100) );
  INVX1 U2290 ( .A(n1522), .Y(n103) );
  INVX1 U2292 ( .A(n1521), .Y(n104) );
  INVX1 U2293 ( .A(n1520), .Y(n105) );
  INVX1 U2295 ( .A(n1517), .Y(n108) );
  INVX1 U2296 ( .A(n1516), .Y(n109) );
  INVX1 U2298 ( .A(n1515), .Y(n110) );
  INVX1 U2299 ( .A(n1497), .Y(n113) );
  INVX1 U2300 ( .A(n1496), .Y(n114) );
  INVX1 U2301 ( .A(n1495), .Y(n115) );
  INVX1 U2303 ( .A(n1492), .Y(n118) );
  INVX1 U2304 ( .A(n1491), .Y(n119) );
  INVX1 U2306 ( .A(n1490), .Y(n120) );
  INVX1 U2307 ( .A(n1470), .Y(n123) );
  INVX1 U2309 ( .A(n1469), .Y(n124) );
  INVX1 U2310 ( .A(n1468), .Y(n125) );
  INVX1 U2312 ( .A(n1465), .Y(n128) );
  INVX1 U2313 ( .A(n1464), .Y(n129) );
  INVX1 U2314 ( .A(n1463), .Y(n130) );
  INVX1 U2315 ( .A(n1445), .Y(n133) );
  INVX1 U2316 ( .A(n1444), .Y(n134) );
  INVX1 U2318 ( .A(n1443), .Y(n135) );
  INVX1 U2320 ( .A(n1440), .Y(n138) );
  INVX1 U2323 ( .A(n1439), .Y(n139) );
  INVX1 U2325 ( .A(n1438), .Y(n140) );
  INVX1 U2328 ( .A(n1418), .Y(n143) );
  INVX1 U2330 ( .A(n1417), .Y(n144) );
  INVX1 U2333 ( .A(n1416), .Y(n145) );
  INVX1 U2337 ( .A(n1413), .Y(n148) );
  INVX1 U2345 ( .A(n1412), .Y(n149) );
  INVX1 U2346 ( .A(n1411), .Y(n150) );
  INVX1 U2347 ( .A(n1392), .Y(n153) );
  INVX1 U2348 ( .A(n1391), .Y(n154) );
  INVX1 U2349 ( .A(n1390), .Y(n155) );
  INVX1 U2350 ( .A(n1387), .Y(n158) );
  INVX1 U2351 ( .A(n1386), .Y(n159) );
  INVX1 U2352 ( .A(n1385), .Y(n160) );
  INVX1 U2353 ( .A(n161), .Y(n162) );
  INVX1 U2354 ( .A(n163), .Y(n164) );
  OR2X1 U2355 ( .A(N182), .B(N181), .Y(n189) );
  INVX1 U2356 ( .A(rst), .Y(n3188) );
  OR2X1 U2357 ( .A(n189), .B(N180), .Y(n191) );
  OR2X1 U2358 ( .A(n2354), .B(n2355), .Y(n192) );
  OR2X1 U2359 ( .A(n2357), .B(n2358), .Y(n193) );
  OR2X1 U2360 ( .A(n2360), .B(n2361), .Y(n194) );
  OR2X1 U2361 ( .A(n2363), .B(n2364), .Y(n195) );
  OR2X1 U2362 ( .A(n2366), .B(n2367), .Y(n196) );
  OR2X1 U2363 ( .A(n2369), .B(n2370), .Y(n197) );
  OR2X1 U2364 ( .A(n2372), .B(n2373), .Y(n198) );
  OR2X1 U2365 ( .A(n2375), .B(n2376), .Y(n199) );
  OR2X1 U2366 ( .A(n2378), .B(n2379), .Y(n200) );
  OR2X1 U2367 ( .A(n2381), .B(n2382), .Y(n201) );
  OR2X1 U2368 ( .A(n2384), .B(n2385), .Y(n202) );
  OR2X1 U2369 ( .A(n2387), .B(n2388), .Y(n203) );
  OR2X1 U2370 ( .A(n2390), .B(n2391), .Y(n204) );
  OR2X1 U2371 ( .A(n2393), .B(n2394), .Y(n205) );
  OR2X1 U2372 ( .A(n2396), .B(n2397), .Y(n206) );
  OR2X1 U2373 ( .A(n2399), .B(n2400), .Y(n207) );
  OR2X1 U2374 ( .A(n2404), .B(n209), .Y(n208) );
  OR2X1 U2375 ( .A(n2402), .B(n2403), .Y(n209) );
  OR2X1 U2376 ( .A(n2405), .B(n2406), .Y(n210) );
  OR2X1 U2377 ( .A(n2410), .B(n212), .Y(n211) );
  OR2X1 U2378 ( .A(n2408), .B(n2409), .Y(n212) );
  OR2X1 U2379 ( .A(n2411), .B(n2412), .Y(n213) );
  OR2X1 U2380 ( .A(n2416), .B(n215), .Y(n214) );
  OR2X1 U2381 ( .A(n2414), .B(n2415), .Y(n215) );
  OR2X1 U2382 ( .A(n2417), .B(n2418), .Y(n216) );
  OR2X1 U2383 ( .A(n2422), .B(n218), .Y(n217) );
  OR2X1 U2384 ( .A(n2420), .B(n2421), .Y(n218) );
  OR2X1 U2385 ( .A(n2423), .B(n2424), .Y(n219) );
  OR2X1 U2386 ( .A(n2428), .B(n221), .Y(n220) );
  OR2X1 U2387 ( .A(n2426), .B(n2427), .Y(n221) );
  OR2X1 U2388 ( .A(n2429), .B(n2430), .Y(n222) );
  OR2X1 U2389 ( .A(n2434), .B(n224), .Y(n223) );
  OR2X1 U2390 ( .A(n2432), .B(n2433), .Y(n224) );
  OR2X1 U2391 ( .A(n2435), .B(n2436), .Y(n225) );
  OR2X1 U2392 ( .A(n2440), .B(n227), .Y(n226) );
  OR2X1 U2393 ( .A(n2438), .B(n2439), .Y(n227) );
  OR2X1 U2394 ( .A(n2441), .B(n2442), .Y(n228) );
  OR2X1 U2395 ( .A(n2446), .B(n230), .Y(n229) );
  OR2X1 U2396 ( .A(n2444), .B(n2445), .Y(n230) );
  OR2X1 U2397 ( .A(n2447), .B(n2448), .Y(n231) );
  BUFX2 U2398 ( .A(n1356), .Y(n232) );
  BUFX2 U2399 ( .A(n1355), .Y(n233) );
  BUFX2 U2400 ( .A(n1354), .Y(n234) );
  BUFX2 U2401 ( .A(n1353), .Y(n235) );
  BUFX2 U2402 ( .A(n1352), .Y(n236) );
  BUFX2 U2403 ( .A(n1351), .Y(n237) );
  BUFX2 U2404 ( .A(n1350), .Y(n238) );
  BUFX2 U2405 ( .A(n1347), .Y(n239) );
  BUFX2 U2406 ( .A(n1344), .Y(n240) );
  BUFX2 U2407 ( .A(n1343), .Y(n241) );
  BUFX2 U2408 ( .A(n1342), .Y(n242) );
  BUFX2 U2409 ( .A(n1341), .Y(n243) );
  BUFX2 U2410 ( .A(n1340), .Y(n244) );
  BUFX2 U2411 ( .A(n1339), .Y(n245) );
  BUFX2 U2412 ( .A(n1338), .Y(n246) );
  BUFX2 U2413 ( .A(n1335), .Y(n247) );
  BUFX2 U2414 ( .A(n1332), .Y(n248) );
  BUFX2 U2415 ( .A(n1331), .Y(n249) );
  BUFX2 U2416 ( .A(n1330), .Y(n250) );
  BUFX2 U2417 ( .A(n1329), .Y(n251) );
  BUFX2 U2418 ( .A(n1328), .Y(n252) );
  BUFX2 U2419 ( .A(n1327), .Y(n253) );
  BUFX2 U2420 ( .A(n1326), .Y(n254) );
  BUFX2 U2421 ( .A(n1323), .Y(n255) );
  BUFX2 U2422 ( .A(n1320), .Y(n256) );
  BUFX2 U2423 ( .A(n1319), .Y(n257) );
  BUFX2 U2424 ( .A(n1318), .Y(n258) );
  BUFX2 U2425 ( .A(n1317), .Y(n259) );
  BUFX2 U2426 ( .A(n1316), .Y(n260) );
  BUFX2 U2427 ( .A(n1315), .Y(n261) );
  BUFX2 U2428 ( .A(n1314), .Y(n262) );
  BUFX2 U2429 ( .A(n1311), .Y(n263) );
  BUFX2 U2430 ( .A(n1308), .Y(n264) );
  BUFX2 U2431 ( .A(n1307), .Y(n265) );
  BUFX2 U2432 ( .A(n1306), .Y(n266) );
  BUFX2 U2433 ( .A(n1305), .Y(n267) );
  BUFX2 U2434 ( .A(n1304), .Y(n268) );
  BUFX2 U2435 ( .A(n1303), .Y(n269) );
  BUFX2 U2436 ( .A(n1302), .Y(n270) );
  BUFX2 U2437 ( .A(n1299), .Y(n271) );
  BUFX2 U2438 ( .A(n1296), .Y(n272) );
  BUFX2 U2439 ( .A(n1295), .Y(n273) );
  BUFX2 U2440 ( .A(n1294), .Y(n274) );
  BUFX2 U2441 ( .A(n1293), .Y(n275) );
  BUFX2 U2442 ( .A(n1292), .Y(n276) );
  BUFX2 U2443 ( .A(n1291), .Y(n277) );
  BUFX2 U2444 ( .A(n1290), .Y(n278) );
  BUFX2 U2445 ( .A(n1287), .Y(n279) );
  BUFX2 U2446 ( .A(n1284), .Y(n280) );
  BUFX2 U2447 ( .A(n1283), .Y(n281) );
  BUFX2 U2448 ( .A(n1282), .Y(n282) );
  BUFX2 U2449 ( .A(n1281), .Y(n283) );
  BUFX2 U2450 ( .A(n1280), .Y(n284) );
  BUFX2 U2451 ( .A(n1279), .Y(n285) );
  BUFX2 U2452 ( .A(n1278), .Y(n286) );
  BUFX2 U2453 ( .A(n1275), .Y(n287) );
  BUFX2 U2454 ( .A(n1272), .Y(n288) );
  BUFX2 U2455 ( .A(n1271), .Y(n289) );
  BUFX2 U2456 ( .A(n1270), .Y(n290) );
  BUFX2 U2457 ( .A(n1269), .Y(n291) );
  BUFX2 U2458 ( .A(n1268), .Y(n292) );
  BUFX2 U2459 ( .A(n1267), .Y(n293) );
  BUFX2 U2460 ( .A(n1266), .Y(n294) );
  BUFX2 U2461 ( .A(n1263), .Y(n295) );
  BUFX2 U2462 ( .A(n1260), .Y(n296) );
  BUFX2 U2463 ( .A(n1259), .Y(n297) );
  BUFX2 U2464 ( .A(n1258), .Y(n298) );
  BUFX2 U2465 ( .A(n1257), .Y(n299) );
  BUFX2 U2466 ( .A(n1256), .Y(n300) );
  BUFX2 U2467 ( .A(n1255), .Y(n301) );
  BUFX2 U2468 ( .A(n1254), .Y(n302) );
  BUFX2 U2469 ( .A(n1251), .Y(n303) );
  BUFX2 U2470 ( .A(n1248), .Y(n304) );
  BUFX2 U2471 ( .A(n1247), .Y(n305) );
  BUFX2 U2472 ( .A(n1246), .Y(n306) );
  BUFX2 U2473 ( .A(n1245), .Y(n307) );
  BUFX2 U2474 ( .A(n1244), .Y(n308) );
  BUFX2 U2475 ( .A(n1243), .Y(n309) );
  BUFX2 U2476 ( .A(n1242), .Y(n310) );
  BUFX2 U2477 ( .A(n1239), .Y(n311) );
  BUFX2 U2478 ( .A(n1236), .Y(n312) );
  BUFX2 U2479 ( .A(n1235), .Y(n313) );
  BUFX2 U2480 ( .A(n1234), .Y(n314) );
  BUFX2 U2481 ( .A(n1233), .Y(n315) );
  BUFX2 U2482 ( .A(n1232), .Y(n316) );
  BUFX2 U2483 ( .A(n1231), .Y(n317) );
  BUFX2 U2484 ( .A(n1230), .Y(n318) );
  BUFX2 U2485 ( .A(n1227), .Y(n319) );
  BUFX2 U2486 ( .A(n1224), .Y(n320) );
  BUFX2 U2487 ( .A(n1223), .Y(n321) );
  BUFX2 U2488 ( .A(n1222), .Y(n322) );
  BUFX2 U2489 ( .A(n1221), .Y(n323) );
  BUFX2 U2490 ( .A(n1220), .Y(n324) );
  BUFX2 U2491 ( .A(n1219), .Y(n325) );
  BUFX2 U2492 ( .A(n1218), .Y(n326) );
  BUFX2 U2493 ( .A(n1215), .Y(n327) );
  BUFX2 U2494 ( .A(n1212), .Y(n328) );
  BUFX2 U2495 ( .A(n1211), .Y(n329) );
  BUFX2 U2496 ( .A(n1210), .Y(n330) );
  BUFX2 U2497 ( .A(n1209), .Y(n331) );
  BUFX2 U2498 ( .A(n1208), .Y(n332) );
  BUFX2 U2499 ( .A(n1207), .Y(n333) );
  BUFX2 U2500 ( .A(n1206), .Y(n334) );
  BUFX2 U2501 ( .A(n1203), .Y(n335) );
  BUFX2 U2502 ( .A(n1200), .Y(n336) );
  BUFX2 U2503 ( .A(n1199), .Y(n337) );
  BUFX2 U2504 ( .A(n1198), .Y(n338) );
  BUFX2 U2505 ( .A(n1197), .Y(n339) );
  BUFX2 U2506 ( .A(n1196), .Y(n340) );
  BUFX2 U2507 ( .A(n1195), .Y(n341) );
  BUFX2 U2508 ( .A(n1194), .Y(n342) );
  BUFX2 U2509 ( .A(n1191), .Y(n343) );
  BUFX2 U2510 ( .A(n1188), .Y(n344) );
  BUFX2 U2511 ( .A(n1187), .Y(n345) );
  BUFX2 U2512 ( .A(n1186), .Y(n346) );
  BUFX2 U2513 ( .A(n1185), .Y(n347) );
  BUFX2 U2514 ( .A(n1184), .Y(n348) );
  BUFX2 U2515 ( .A(n1183), .Y(n349) );
  BUFX2 U2516 ( .A(n1182), .Y(n350) );
  BUFX2 U2517 ( .A(n1179), .Y(n351) );
  BUFX2 U2518 ( .A(n1176), .Y(n352) );
  BUFX2 U2519 ( .A(n1175), .Y(n353) );
  BUFX2 U2520 ( .A(n1174), .Y(n354) );
  BUFX2 U2521 ( .A(n1173), .Y(n355) );
  BUFX2 U2522 ( .A(n1172), .Y(n356) );
  BUFX2 U2523 ( .A(n1171), .Y(n357) );
  BUFX2 U2524 ( .A(n1170), .Y(n358) );
  BUFX2 U2525 ( .A(n1167), .Y(n359) );
  BUFX2 U2526 ( .A(n1164), .Y(n360) );
  BUFX2 U2527 ( .A(n1163), .Y(n361) );
  BUFX2 U2528 ( .A(n1162), .Y(n362) );
  BUFX2 U2529 ( .A(n1161), .Y(n363) );
  BUFX2 U2530 ( .A(n1160), .Y(n364) );
  BUFX2 U2531 ( .A(n1159), .Y(n365) );
  BUFX2 U2532 ( .A(n1158), .Y(n366) );
  BUFX2 U2533 ( .A(n1155), .Y(n367) );
  BUFX2 U2534 ( .A(n1152), .Y(n368) );
  BUFX2 U2535 ( .A(n1151), .Y(n369) );
  BUFX2 U2536 ( .A(n1150), .Y(n370) );
  BUFX2 U2537 ( .A(n1149), .Y(n371) );
  BUFX2 U2538 ( .A(n1148), .Y(n372) );
  BUFX2 U2539 ( .A(n1147), .Y(n373) );
  BUFX2 U2540 ( .A(n1146), .Y(n374) );
  BUFX2 U2541 ( .A(n1143), .Y(n375) );
  BUFX2 U2542 ( .A(n1140), .Y(n376) );
  BUFX2 U2543 ( .A(n1139), .Y(n377) );
  BUFX2 U2544 ( .A(n1138), .Y(n378) );
  BUFX2 U2545 ( .A(n1137), .Y(n379) );
  BUFX2 U2546 ( .A(n1136), .Y(n380) );
  BUFX2 U2547 ( .A(n1135), .Y(n381) );
  BUFX2 U2548 ( .A(n1134), .Y(n382) );
  BUFX2 U2549 ( .A(n1131), .Y(n383) );
  BUFX2 U2550 ( .A(n1128), .Y(n384) );
  BUFX2 U2551 ( .A(n1127), .Y(n385) );
  BUFX2 U2552 ( .A(n1126), .Y(n386) );
  BUFX2 U2553 ( .A(n1125), .Y(n387) );
  BUFX2 U2554 ( .A(n1124), .Y(n388) );
  BUFX2 U2555 ( .A(n1123), .Y(n389) );
  BUFX2 U2556 ( .A(n1122), .Y(n390) );
  BUFX2 U2557 ( .A(n1119), .Y(n391) );
  BUFX2 U2558 ( .A(n1116), .Y(n392) );
  BUFX2 U2559 ( .A(n1115), .Y(n393) );
  BUFX2 U2560 ( .A(n1114), .Y(n394) );
  BUFX2 U2561 ( .A(n1113), .Y(n395) );
  BUFX2 U2562 ( .A(n1112), .Y(n396) );
  BUFX2 U2563 ( .A(n1111), .Y(n397) );
  BUFX2 U2564 ( .A(n1110), .Y(n398) );
  BUFX2 U2565 ( .A(n1107), .Y(n399) );
  BUFX2 U2566 ( .A(n1104), .Y(n400) );
  BUFX2 U2567 ( .A(n1103), .Y(n401) );
  BUFX2 U2568 ( .A(n1102), .Y(n402) );
  BUFX2 U2569 ( .A(n1101), .Y(n403) );
  BUFX2 U2570 ( .A(n1100), .Y(n404) );
  BUFX2 U2571 ( .A(n1099), .Y(n405) );
  BUFX2 U2572 ( .A(n1098), .Y(n406) );
  BUFX2 U2573 ( .A(n1095), .Y(n407) );
  BUFX2 U2574 ( .A(n1092), .Y(n408) );
  BUFX2 U2575 ( .A(n1091), .Y(n409) );
  BUFX2 U2576 ( .A(n1090), .Y(n410) );
  BUFX2 U2577 ( .A(n1089), .Y(n411) );
  BUFX2 U2578 ( .A(n1088), .Y(n412) );
  BUFX2 U2579 ( .A(n1087), .Y(n413) );
  BUFX2 U2580 ( .A(n1086), .Y(n414) );
  BUFX2 U2581 ( .A(n1083), .Y(n415) );
  BUFX2 U2582 ( .A(n1080), .Y(n416) );
  BUFX2 U2583 ( .A(n1079), .Y(n417) );
  BUFX2 U2584 ( .A(n1078), .Y(n418) );
  BUFX2 U2585 ( .A(n1077), .Y(n419) );
  BUFX2 U2586 ( .A(n1076), .Y(n420) );
  BUFX2 U2587 ( .A(n1075), .Y(n421) );
  BUFX2 U2588 ( .A(n1074), .Y(n422) );
  BUFX2 U2589 ( .A(n1071), .Y(n423) );
  BUFX2 U2590 ( .A(n1068), .Y(n424) );
  BUFX2 U2591 ( .A(n1067), .Y(n425) );
  BUFX2 U2592 ( .A(n1066), .Y(n426) );
  BUFX2 U2593 ( .A(n1065), .Y(n427) );
  BUFX2 U2594 ( .A(n1064), .Y(n428) );
  BUFX2 U2595 ( .A(n1063), .Y(n429) );
  BUFX2 U2596 ( .A(n1062), .Y(n430) );
  BUFX2 U2597 ( .A(n1059), .Y(n431) );
  BUFX2 U2598 ( .A(n1056), .Y(n432) );
  BUFX2 U2599 ( .A(n1055), .Y(n433) );
  BUFX2 U2600 ( .A(n1054), .Y(n434) );
  BUFX2 U2601 ( .A(n1053), .Y(n435) );
  BUFX2 U2602 ( .A(n1052), .Y(n436) );
  BUFX2 U2603 ( .A(n1051), .Y(n437) );
  BUFX2 U2604 ( .A(n1050), .Y(n438) );
  BUFX2 U2605 ( .A(n1047), .Y(n439) );
  BUFX2 U2606 ( .A(n1044), .Y(n440) );
  BUFX2 U2607 ( .A(n1043), .Y(n441) );
  BUFX2 U2608 ( .A(n1042), .Y(n442) );
  BUFX2 U2609 ( .A(n1041), .Y(n443) );
  BUFX2 U2610 ( .A(n1040), .Y(n444) );
  BUFX2 U2611 ( .A(n1039), .Y(n445) );
  BUFX2 U2612 ( .A(n1038), .Y(n446) );
  BUFX2 U2613 ( .A(n1035), .Y(n447) );
  BUFX2 U2614 ( .A(n1032), .Y(n448) );
  BUFX2 U2615 ( .A(n1031), .Y(n449) );
  BUFX2 U2616 ( .A(n1030), .Y(n450) );
  BUFX2 U2617 ( .A(n1029), .Y(n451) );
  BUFX2 U2618 ( .A(n1028), .Y(n452) );
  BUFX2 U2619 ( .A(n1027), .Y(n453) );
  BUFX2 U2620 ( .A(n1026), .Y(n454) );
  BUFX2 U2621 ( .A(n1023), .Y(n455) );
  BUFX2 U2622 ( .A(n1020), .Y(n456) );
  BUFX2 U2623 ( .A(n1019), .Y(n457) );
  BUFX2 U2624 ( .A(n1018), .Y(n458) );
  BUFX2 U2625 ( .A(n1017), .Y(n459) );
  BUFX2 U2626 ( .A(n1016), .Y(n460) );
  BUFX2 U2627 ( .A(n1015), .Y(n461) );
  BUFX2 U2628 ( .A(n1014), .Y(n462) );
  BUFX2 U2629 ( .A(n1011), .Y(n463) );
  BUFX2 U2630 ( .A(n1008), .Y(n464) );
  BUFX2 U2631 ( .A(n1007), .Y(n465) );
  BUFX2 U2632 ( .A(n1006), .Y(n466) );
  BUFX2 U2633 ( .A(n1005), .Y(n467) );
  BUFX2 U2634 ( .A(n1004), .Y(n468) );
  BUFX2 U2635 ( .A(n1003), .Y(n469) );
  BUFX2 U2636 ( .A(n1002), .Y(n470) );
  BUFX2 U2637 ( .A(n999), .Y(n471) );
  BUFX2 U2638 ( .A(n996), .Y(n472) );
  BUFX2 U2639 ( .A(n995), .Y(n473) );
  BUFX2 U2640 ( .A(n994), .Y(n474) );
  BUFX2 U2641 ( .A(n993), .Y(n475) );
  BUFX2 U2642 ( .A(n992), .Y(n476) );
  BUFX2 U2643 ( .A(n991), .Y(n477) );
  BUFX2 U2644 ( .A(n990), .Y(n478) );
  BUFX2 U2645 ( .A(n987), .Y(n479) );
  BUFX2 U2646 ( .A(n984), .Y(n480) );
  BUFX2 U2647 ( .A(n983), .Y(n481) );
  BUFX2 U2648 ( .A(n982), .Y(n482) );
  BUFX2 U2649 ( .A(n981), .Y(n483) );
  BUFX2 U2650 ( .A(n980), .Y(n484) );
  BUFX2 U2651 ( .A(n979), .Y(n485) );
  BUFX2 U2652 ( .A(n978), .Y(n486) );
  BUFX2 U2653 ( .A(n975), .Y(n487) );
  BUFX2 U2654 ( .A(n972), .Y(n488) );
  BUFX2 U2655 ( .A(n971), .Y(n489) );
  BUFX2 U2656 ( .A(n970), .Y(n490) );
  BUFX2 U2657 ( .A(n969), .Y(n491) );
  BUFX2 U2658 ( .A(n968), .Y(n492) );
  BUFX2 U2659 ( .A(n967), .Y(n493) );
  BUFX2 U2660 ( .A(n966), .Y(n494) );
  BUFX2 U2661 ( .A(n963), .Y(n495) );
  BUFX2 U2662 ( .A(n960), .Y(n496) );
  BUFX2 U2663 ( .A(n959), .Y(n497) );
  BUFX2 U2664 ( .A(n958), .Y(n498) );
  BUFX2 U2665 ( .A(n957), .Y(n499) );
  BUFX2 U2666 ( .A(n956), .Y(n500) );
  BUFX2 U2667 ( .A(n955), .Y(n501) );
  BUFX2 U2668 ( .A(n954), .Y(n502) );
  BUFX2 U2669 ( .A(n951), .Y(n503) );
  BUFX2 U2670 ( .A(n948), .Y(n504) );
  BUFX2 U2671 ( .A(n947), .Y(n505) );
  BUFX2 U2672 ( .A(n946), .Y(n506) );
  BUFX2 U2673 ( .A(n945), .Y(n507) );
  BUFX2 U2674 ( .A(n944), .Y(n508) );
  BUFX2 U2675 ( .A(n943), .Y(n509) );
  BUFX2 U2676 ( .A(n942), .Y(n510) );
  BUFX2 U2677 ( .A(n939), .Y(n511) );
  BUFX2 U2678 ( .A(n936), .Y(n512) );
  BUFX2 U2679 ( .A(n935), .Y(n513) );
  BUFX2 U2680 ( .A(n934), .Y(n514) );
  BUFX2 U2681 ( .A(n933), .Y(n515) );
  BUFX2 U2682 ( .A(n932), .Y(n516) );
  BUFX2 U2683 ( .A(n931), .Y(n517) );
  BUFX2 U2684 ( .A(n930), .Y(n518) );
  BUFX2 U2685 ( .A(n927), .Y(n519) );
  BUFX2 U2686 ( .A(n924), .Y(n520) );
  BUFX2 U2687 ( .A(n923), .Y(n521) );
  BUFX2 U2688 ( .A(n922), .Y(n522) );
  BUFX2 U2689 ( .A(n921), .Y(n523) );
  BUFX2 U2690 ( .A(n920), .Y(n524) );
  BUFX2 U2691 ( .A(n919), .Y(n525) );
  BUFX2 U2692 ( .A(n918), .Y(n526) );
  BUFX2 U2693 ( .A(n915), .Y(n527) );
  BUFX2 U2694 ( .A(n912), .Y(n528) );
  BUFX2 U2695 ( .A(n911), .Y(n529) );
  BUFX2 U2696 ( .A(n910), .Y(n530) );
  BUFX2 U2697 ( .A(n909), .Y(n531) );
  BUFX2 U2698 ( .A(n908), .Y(n532) );
  BUFX2 U2699 ( .A(n907), .Y(n533) );
  BUFX2 U2700 ( .A(n906), .Y(n534) );
  BUFX2 U2701 ( .A(n903), .Y(n535) );
  BUFX2 U2702 ( .A(n900), .Y(n536) );
  BUFX2 U2703 ( .A(n899), .Y(n537) );
  BUFX2 U2704 ( .A(n898), .Y(n538) );
  BUFX2 U2705 ( .A(n897), .Y(n539) );
  BUFX2 U2706 ( .A(n896), .Y(n540) );
  BUFX2 U2707 ( .A(n895), .Y(n541) );
  BUFX2 U2708 ( .A(n894), .Y(n542) );
  BUFX2 U2709 ( .A(n891), .Y(n543) );
  BUFX2 U2710 ( .A(n888), .Y(n544) );
  BUFX2 U2711 ( .A(n887), .Y(n545) );
  BUFX2 U2712 ( .A(n886), .Y(n546) );
  BUFX2 U2713 ( .A(n885), .Y(n547) );
  BUFX2 U2714 ( .A(n884), .Y(n548) );
  BUFX2 U2715 ( .A(n883), .Y(n549) );
  BUFX2 U2716 ( .A(n882), .Y(n550) );
  BUFX2 U2717 ( .A(n879), .Y(n551) );
  BUFX2 U2718 ( .A(n876), .Y(n552) );
  BUFX2 U2719 ( .A(n875), .Y(n553) );
  BUFX2 U2720 ( .A(n874), .Y(n554) );
  BUFX2 U2721 ( .A(n873), .Y(n555) );
  BUFX2 U2722 ( .A(n872), .Y(n556) );
  BUFX2 U2723 ( .A(n871), .Y(n557) );
  BUFX2 U2724 ( .A(n870), .Y(n558) );
  BUFX2 U2725 ( .A(n867), .Y(n559) );
  BUFX2 U2726 ( .A(n864), .Y(n560) );
  BUFX2 U2727 ( .A(n863), .Y(n561) );
  BUFX2 U2728 ( .A(n862), .Y(n562) );
  BUFX2 U2729 ( .A(n861), .Y(n563) );
  BUFX2 U2730 ( .A(n860), .Y(n564) );
  BUFX2 U2731 ( .A(n859), .Y(n565) );
  BUFX2 U2732 ( .A(n858), .Y(n566) );
  BUFX2 U2733 ( .A(n855), .Y(n567) );
  BUFX2 U2734 ( .A(n852), .Y(n568) );
  BUFX2 U2735 ( .A(n851), .Y(n569) );
  BUFX2 U2736 ( .A(n850), .Y(n570) );
  BUFX2 U2737 ( .A(n849), .Y(n571) );
  BUFX2 U2738 ( .A(n848), .Y(n572) );
  BUFX2 U2739 ( .A(n847), .Y(n573) );
  BUFX2 U2740 ( .A(n846), .Y(n574) );
  BUFX2 U2741 ( .A(n843), .Y(n575) );
  BUFX2 U2742 ( .A(n840), .Y(n576) );
  BUFX2 U2743 ( .A(n839), .Y(n577) );
  BUFX2 U2744 ( .A(n838), .Y(n578) );
  BUFX2 U2745 ( .A(n837), .Y(n579) );
  BUFX2 U2746 ( .A(n836), .Y(n580) );
  BUFX2 U2747 ( .A(n835), .Y(n581) );
  BUFX2 U2748 ( .A(n834), .Y(n582) );
  BUFX2 U2749 ( .A(n831), .Y(n583) );
  BUFX2 U2750 ( .A(n828), .Y(n584) );
  BUFX2 U2751 ( .A(n827), .Y(n585) );
  BUFX2 U2752 ( .A(n826), .Y(n586) );
  BUFX2 U2753 ( .A(n825), .Y(n587) );
  BUFX2 U2754 ( .A(n824), .Y(n588) );
  BUFX2 U2755 ( .A(n823), .Y(n589) );
  BUFX2 U2756 ( .A(n822), .Y(n590) );
  BUFX2 U2757 ( .A(n819), .Y(n591) );
  BUFX2 U2758 ( .A(n816), .Y(n592) );
  BUFX2 U2759 ( .A(n815), .Y(n593) );
  BUFX2 U2760 ( .A(n814), .Y(n594) );
  BUFX2 U2761 ( .A(n813), .Y(n595) );
  BUFX2 U2762 ( .A(n812), .Y(n596) );
  BUFX2 U2763 ( .A(n811), .Y(n597) );
  BUFX2 U2764 ( .A(n810), .Y(n609) );
  BUFX2 U2765 ( .A(n807), .Y(n611) );
  BUFX2 U2766 ( .A(n804), .Y(n624) );
  BUFX2 U2767 ( .A(n803), .Y(n637) );
  BUFX2 U2768 ( .A(n802), .Y(n649) );
  BUFX2 U2769 ( .A(n801), .Y(n661) );
  BUFX2 U2770 ( .A(n800), .Y(n673) );
  BUFX2 U2771 ( .A(n799), .Y(n685) );
  BUFX2 U2772 ( .A(n798), .Y(n697) );
  BUFX2 U2773 ( .A(n795), .Y(n709) );
  BUFX2 U2774 ( .A(n792), .Y(n721) );
  BUFX2 U2775 ( .A(n791), .Y(n733) );
  BUFX2 U2776 ( .A(n790), .Y(n745) );
  BUFX2 U2777 ( .A(n789), .Y(n757) );
  BUFX2 U2778 ( .A(n788), .Y(n769) );
  BUFX2 U2779 ( .A(n787), .Y(n781) );
  BUFX2 U2780 ( .A(n786), .Y(n793) );
  BUFX2 U2781 ( .A(n783), .Y(n805) );
  BUFX2 U2782 ( .A(n780), .Y(n817) );
  BUFX2 U2783 ( .A(n779), .Y(n829) );
  BUFX2 U2784 ( .A(n778), .Y(n841) );
  BUFX2 U2785 ( .A(n777), .Y(n853) );
  BUFX2 U2786 ( .A(n776), .Y(n865) );
  BUFX2 U2787 ( .A(n775), .Y(n877) );
  BUFX2 U2788 ( .A(n774), .Y(n889) );
  BUFX2 U2789 ( .A(n771), .Y(n901) );
  BUFX2 U2790 ( .A(n768), .Y(n913) );
  BUFX2 U2791 ( .A(n767), .Y(n925) );
  BUFX2 U2792 ( .A(n766), .Y(n937) );
  BUFX2 U2793 ( .A(n765), .Y(n949) );
  BUFX2 U2794 ( .A(n764), .Y(n961) );
  BUFX2 U2795 ( .A(n763), .Y(n973) );
  BUFX2 U2796 ( .A(n762), .Y(n985) );
  BUFX2 U2797 ( .A(n759), .Y(n997) );
  BUFX2 U2798 ( .A(n756), .Y(n1009) );
  BUFX2 U2799 ( .A(n755), .Y(n1021) );
  BUFX2 U2800 ( .A(n754), .Y(n1033) );
  BUFX2 U2801 ( .A(n753), .Y(n1045) );
  BUFX2 U2802 ( .A(n752), .Y(n1057) );
  BUFX2 U2803 ( .A(n751), .Y(n1069) );
  BUFX2 U2804 ( .A(n750), .Y(n1081) );
  BUFX2 U2805 ( .A(n747), .Y(n1093) );
  BUFX2 U2806 ( .A(n744), .Y(n1105) );
  BUFX2 U2807 ( .A(n743), .Y(n1117) );
  BUFX2 U2808 ( .A(n742), .Y(n1129) );
  BUFX2 U2809 ( .A(n741), .Y(n1141) );
  BUFX2 U2810 ( .A(n740), .Y(n1153) );
  BUFX2 U2811 ( .A(n739), .Y(n1165) );
  BUFX2 U2812 ( .A(n738), .Y(n1177) );
  BUFX2 U2813 ( .A(n735), .Y(n1189) );
  BUFX2 U2814 ( .A(n732), .Y(n1201) );
  BUFX2 U2815 ( .A(n731), .Y(n1213) );
  BUFX2 U2816 ( .A(n730), .Y(n1225) );
  BUFX2 U2817 ( .A(n729), .Y(n1237) );
  BUFX2 U2818 ( .A(n728), .Y(n1249) );
  BUFX2 U2819 ( .A(n727), .Y(n1261) );
  BUFX2 U2820 ( .A(n726), .Y(n1273) );
  BUFX2 U2821 ( .A(n723), .Y(n1285) );
  BUFX2 U2822 ( .A(n720), .Y(n1297) );
  BUFX2 U2823 ( .A(n719), .Y(n1309) );
  BUFX2 U2824 ( .A(n718), .Y(n1321) );
  BUFX2 U2825 ( .A(n717), .Y(n1333) );
  BUFX2 U2826 ( .A(n716), .Y(n1345) );
  BUFX2 U2827 ( .A(n715), .Y(n1357) );
  BUFX2 U2828 ( .A(n714), .Y(n1358) );
  BUFX2 U2829 ( .A(n711), .Y(n1359) );
  BUFX2 U2830 ( .A(n708), .Y(n1360) );
  BUFX2 U2831 ( .A(n707), .Y(n1361) );
  BUFX2 U2832 ( .A(n706), .Y(n1362) );
  BUFX2 U2833 ( .A(n705), .Y(n1363) );
  BUFX2 U2834 ( .A(n704), .Y(n1364) );
  BUFX2 U2835 ( .A(n703), .Y(n1365) );
  BUFX2 U2836 ( .A(n702), .Y(n1366) );
  BUFX2 U2837 ( .A(n699), .Y(n1369) );
  BUFX2 U2838 ( .A(n696), .Y(n1371) );
  BUFX2 U2839 ( .A(n695), .Y(n1372) );
  BUFX2 U2840 ( .A(n694), .Y(n1383) );
  BUFX2 U2841 ( .A(n693), .Y(n1384) );
  BUFX2 U2842 ( .A(n692), .Y(n1396) );
  BUFX2 U2843 ( .A(n691), .Y(n1397) );
  BUFX2 U2844 ( .A(n690), .Y(n1409) );
  BUFX2 U2845 ( .A(n687), .Y(n1410) );
  BUFX2 U2846 ( .A(n684), .Y(n1424) );
  BUFX2 U2847 ( .A(n683), .Y(n1425) );
  BUFX2 U2848 ( .A(n682), .Y(n1436) );
  BUFX2 U2849 ( .A(n681), .Y(n1437) );
  BUFX2 U2850 ( .A(n680), .Y(n1449) );
  BUFX2 U2851 ( .A(n679), .Y(n1450) );
  BUFX2 U2852 ( .A(n678), .Y(n1461) );
  BUFX2 U2853 ( .A(n675), .Y(n1462) );
  BUFX2 U2854 ( .A(n672), .Y(n1476) );
  BUFX2 U2855 ( .A(n671), .Y(n1477) );
  BUFX2 U2856 ( .A(n670), .Y(n1488) );
  BUFX2 U2857 ( .A(n669), .Y(n1489) );
  BUFX2 U2858 ( .A(n668), .Y(n1501) );
  BUFX2 U2859 ( .A(n667), .Y(n1502) );
  BUFX2 U2860 ( .A(n666), .Y(n1513) );
  BUFX2 U2861 ( .A(n663), .Y(n1514) );
  BUFX2 U2862 ( .A(n660), .Y(n1528) );
  BUFX2 U2863 ( .A(n659), .Y(n1529) );
  BUFX2 U2864 ( .A(n658), .Y(n1540) );
  BUFX2 U2865 ( .A(n657), .Y(n1541) );
  BUFX2 U2866 ( .A(n656), .Y(n1553) );
  BUFX2 U2867 ( .A(n655), .Y(n1554) );
  BUFX2 U2868 ( .A(n654), .Y(n1565) );
  BUFX2 U2869 ( .A(n651), .Y(n1566) );
  BUFX2 U2870 ( .A(n648), .Y(n1580) );
  BUFX2 U2871 ( .A(n647), .Y(n1581) );
  BUFX2 U2872 ( .A(n646), .Y(n1592) );
  BUFX2 U2873 ( .A(n645), .Y(n1593) );
  BUFX2 U2874 ( .A(n644), .Y(n1605) );
  BUFX2 U2875 ( .A(n643), .Y(n1606) );
  BUFX2 U2876 ( .A(n642), .Y(n1617) );
  BUFX2 U2877 ( .A(n639), .Y(n1618) );
  BUFX2 U2878 ( .A(n636), .Y(n1632) );
  BUFX2 U2879 ( .A(n635), .Y(n1633) );
  BUFX2 U2880 ( .A(n634), .Y(n1644) );
  BUFX2 U2881 ( .A(n633), .Y(n1645) );
  BUFX2 U2882 ( .A(n632), .Y(n1657) );
  BUFX2 U2883 ( .A(n631), .Y(n1658) );
  BUFX2 U2884 ( .A(n630), .Y(n1669) );
  BUFX2 U2885 ( .A(n627), .Y(n1670) );
  BUFX2 U2886 ( .A(n623), .Y(n1684) );
  BUFX2 U2887 ( .A(n622), .Y(n1685) );
  BUFX2 U2888 ( .A(n621), .Y(n1696) );
  BUFX2 U2889 ( .A(n620), .Y(n1697) );
  BUFX2 U2890 ( .A(n619), .Y(n1709) );
  BUFX2 U2891 ( .A(n618), .Y(n1710) );
  BUFX2 U2892 ( .A(n617), .Y(n1721) );
  BUFX2 U2893 ( .A(n614), .Y(n1722) );
  BUFX2 U2894 ( .A(n608), .Y(n1736) );
  BUFX2 U2895 ( .A(n607), .Y(n1737) );
  BUFX2 U2896 ( .A(n606), .Y(n1758) );
  BUFX2 U2897 ( .A(n605), .Y(n1759) );
  BUFX2 U2898 ( .A(n604), .Y(n1771) );
  BUFX2 U2899 ( .A(n603), .Y(n1773) );
  BUFX2 U2900 ( .A(n602), .Y(n1775) );
  BUFX2 U2901 ( .A(n599), .Y(n1776) );
  AND2X1 U2902 ( .A(n3190), .B(\data_in<15> ), .Y(n1793) );
  INVX1 U2903 ( .A(n1793), .Y(n1794) );
  AND2X1 U2904 ( .A(n3190), .B(\data_in<14> ), .Y(n1795) );
  INVX1 U2905 ( .A(n1795), .Y(n1796) );
  AND2X1 U2906 ( .A(n3190), .B(\data_in<13> ), .Y(n1802) );
  INVX1 U2907 ( .A(n1802), .Y(n2328) );
  AND2X1 U2908 ( .A(n3190), .B(\data_in<12> ), .Y(n2329) );
  INVX1 U2909 ( .A(n2329), .Y(n2330) );
  AND2X1 U2910 ( .A(n3190), .B(\data_in<11> ), .Y(n2331) );
  INVX1 U2911 ( .A(n2331), .Y(n2332) );
  AND2X1 U2912 ( .A(n3190), .B(\data_in<10> ), .Y(n2333) );
  INVX1 U2913 ( .A(n2333), .Y(n2334) );
  AND2X1 U2914 ( .A(n3190), .B(\data_in<9> ), .Y(n2335) );
  INVX1 U2915 ( .A(n2335), .Y(n2336) );
  AND2X1 U2916 ( .A(n3190), .B(\data_in<8> ), .Y(n2337) );
  INVX1 U2917 ( .A(n2337), .Y(n2338) );
  BUFX2 U2918 ( .A(n1810), .Y(n2339) );
  INVX1 U2919 ( .A(n2339), .Y(n3191) );
  BUFX2 U2920 ( .A(n1808), .Y(n2340) );
  INVX1 U2921 ( .A(n2340), .Y(n3196) );
  INVX1 U2922 ( .A(n1756), .Y(n2341) );
  INVX1 U2923 ( .A(n1787), .Y(n3195) );
  INVX1 U2924 ( .A(n1772), .Y(n3192) );
  INVX1 U2925 ( .A(n1770), .Y(n3194) );
  INVX1 U2926 ( .A(n1755), .Y(n3193) );
  BUFX2 U2927 ( .A(n3719), .Y(\data_out<0> ) );
  BUFX2 U2928 ( .A(n3718), .Y(\data_out<1> ) );
  BUFX2 U2929 ( .A(n3717), .Y(\data_out<2> ) );
  BUFX2 U2930 ( .A(n3716), .Y(\data_out<3> ) );
  BUFX2 U2931 ( .A(n3715), .Y(\data_out<4> ) );
  BUFX2 U2932 ( .A(n3714), .Y(\data_out<5> ) );
  BUFX2 U2933 ( .A(n3713), .Y(\data_out<6> ) );
  BUFX2 U2934 ( .A(n3712), .Y(\data_out<7> ) );
  OR2X1 U2935 ( .A(N181), .B(n3187), .Y(n2350) );
  INVX1 U2936 ( .A(n2350), .Y(n2351) );
  OR2X1 U2937 ( .A(N181), .B(N180), .Y(n2352) );
  INVX1 U2938 ( .A(n2352), .Y(n2353) );
  INVX1 U2939 ( .A(n1790), .Y(n2354) );
  INVX1 U2940 ( .A(n1789), .Y(n2355) );
  INVX1 U2941 ( .A(n1788), .Y(n2356) );
  INVX1 U2942 ( .A(n612), .Y(n3189) );
  INVX1 U2943 ( .A(n1752), .Y(n2357) );
  INVX1 U2944 ( .A(n1751), .Y(n2358) );
  INVX1 U2945 ( .A(n1750), .Y(n2359) );
  INVX1 U2946 ( .A(n1718), .Y(n2360) );
  INVX1 U2947 ( .A(n1717), .Y(n2361) );
  INVX1 U2948 ( .A(n1716), .Y(n2362) );
  INVX1 U2949 ( .A(n1693), .Y(n2363) );
  INVX1 U2950 ( .A(n1692), .Y(n2364) );
  INVX1 U2951 ( .A(n1691), .Y(n2365) );
  INVX1 U2952 ( .A(n1666), .Y(n2366) );
  INVX1 U2953 ( .A(n1665), .Y(n2367) );
  INVX1 U2954 ( .A(n1664), .Y(n2368) );
  INVX1 U2955 ( .A(n1641), .Y(n2369) );
  INVX1 U2956 ( .A(n1640), .Y(n2370) );
  INVX1 U2957 ( .A(n1639), .Y(n2371) );
  INVX1 U2958 ( .A(n1614), .Y(n2372) );
  INVX1 U2959 ( .A(n1613), .Y(n2373) );
  INVX1 U2960 ( .A(n1612), .Y(n2374) );
  INVX1 U2961 ( .A(n1589), .Y(n2375) );
  INVX1 U2962 ( .A(n1588), .Y(n2376) );
  INVX1 U2963 ( .A(n1587), .Y(n2377) );
  INVX1 U2964 ( .A(n1562), .Y(n2378) );
  INVX1 U2965 ( .A(n1561), .Y(n2379) );
  INVX1 U2966 ( .A(n1560), .Y(n2380) );
  INVX1 U2967 ( .A(n1537), .Y(n2381) );
  INVX1 U2968 ( .A(n1536), .Y(n2382) );
  INVX1 U2969 ( .A(n1535), .Y(n2383) );
  INVX1 U2970 ( .A(n1510), .Y(n2384) );
  INVX1 U2971 ( .A(n1509), .Y(n2385) );
  INVX1 U2972 ( .A(n1508), .Y(n2386) );
  INVX1 U2973 ( .A(n1485), .Y(n2387) );
  INVX1 U2974 ( .A(n1484), .Y(n2388) );
  INVX1 U2975 ( .A(n1483), .Y(n2389) );
  INVX1 U2976 ( .A(n1458), .Y(n2390) );
  INVX1 U2977 ( .A(n1457), .Y(n2391) );
  INVX1 U2978 ( .A(n1456), .Y(n2392) );
  INVX1 U2979 ( .A(n1433), .Y(n2393) );
  INVX1 U2980 ( .A(n1432), .Y(n2394) );
  INVX1 U2981 ( .A(n1431), .Y(n2395) );
  INVX1 U2982 ( .A(n1406), .Y(n2396) );
  INVX1 U2983 ( .A(n1405), .Y(n2397) );
  INVX1 U2984 ( .A(n1404), .Y(n2398) );
  INVX1 U2985 ( .A(n1380), .Y(n2399) );
  INVX1 U2986 ( .A(n1379), .Y(n2400) );
  INVX1 U2987 ( .A(n1378), .Y(n2401) );
  INVX1 U2988 ( .A(n1779), .Y(n2402) );
  INVX1 U2989 ( .A(n1778), .Y(n2403) );
  INVX1 U2990 ( .A(n1777), .Y(n2404) );
  INVX1 U2991 ( .A(n1740), .Y(n2405) );
  INVX1 U2992 ( .A(n1739), .Y(n2406) );
  INVX1 U2993 ( .A(n1738), .Y(n2407) );
  INVX1 U2994 ( .A(n1713), .Y(n2408) );
  INVX1 U2995 ( .A(n1712), .Y(n2409) );
  INVX1 U2996 ( .A(n1711), .Y(n2410) );
  INVX1 U2997 ( .A(n1688), .Y(n2411) );
  INVX1 U2998 ( .A(n1687), .Y(n2412) );
  INVX1 U2999 ( .A(n1686), .Y(n2413) );
  INVX1 U3000 ( .A(n1661), .Y(n2414) );
  INVX1 U3001 ( .A(n1660), .Y(n2415) );
  INVX1 U3002 ( .A(n1659), .Y(n2416) );
  INVX1 U3003 ( .A(n1636), .Y(n2417) );
  INVX1 U3004 ( .A(n1635), .Y(n2418) );
  INVX1 U3005 ( .A(n1634), .Y(n2419) );
  INVX1 U3006 ( .A(n1609), .Y(n2420) );
  INVX1 U3007 ( .A(n1608), .Y(n2421) );
  INVX1 U3008 ( .A(n1607), .Y(n2422) );
  INVX1 U3009 ( .A(n1584), .Y(n2423) );
  INVX1 U3010 ( .A(n1583), .Y(n2424) );
  INVX1 U3011 ( .A(n1582), .Y(n2425) );
  INVX1 U3012 ( .A(n1557), .Y(n2426) );
  INVX1 U3013 ( .A(n1556), .Y(n2427) );
  INVX1 U3014 ( .A(n1555), .Y(n2428) );
  INVX1 U3015 ( .A(n1532), .Y(n2429) );
  INVX1 U3016 ( .A(n1531), .Y(n2430) );
  INVX1 U3017 ( .A(n1530), .Y(n2431) );
  INVX1 U3018 ( .A(n1505), .Y(n2432) );
  INVX1 U3019 ( .A(n1504), .Y(n2433) );
  INVX1 U3020 ( .A(n1503), .Y(n2434) );
  INVX1 U3021 ( .A(n1480), .Y(n2435) );
  INVX1 U3022 ( .A(n1479), .Y(n2436) );
  INVX1 U3023 ( .A(n1478), .Y(n2437) );
  INVX1 U3024 ( .A(n1453), .Y(n2438) );
  INVX1 U3025 ( .A(n1452), .Y(n2439) );
  INVX1 U3026 ( .A(n1451), .Y(n2440) );
  INVX1 U3027 ( .A(n1428), .Y(n2441) );
  INVX1 U3028 ( .A(n1427), .Y(n2442) );
  INVX1 U3029 ( .A(n1426), .Y(n2443) );
  INVX1 U3030 ( .A(n1400), .Y(n2444) );
  INVX1 U3031 ( .A(n1399), .Y(n2445) );
  INVX1 U3032 ( .A(n1398), .Y(n2446) );
  INVX1 U3033 ( .A(n1375), .Y(n2447) );
  INVX1 U3034 ( .A(n1374), .Y(n2448) );
  INVX1 U3035 ( .A(n1373), .Y(n2449) );
  BUFX2 U3036 ( .A(n1334), .Y(n3115) );
  BUFX2 U3037 ( .A(n1322), .Y(n3116) );
  BUFX2 U3038 ( .A(n1310), .Y(n3117) );
  BUFX2 U3039 ( .A(n1298), .Y(n3118) );
  BUFX2 U3040 ( .A(n1286), .Y(n3119) );
  BUFX2 U3041 ( .A(n1274), .Y(n3120) );
  BUFX2 U3042 ( .A(n1262), .Y(n3121) );
  BUFX2 U3043 ( .A(n1250), .Y(n3122) );
  BUFX2 U3044 ( .A(n1238), .Y(n3123) );
  BUFX2 U3045 ( .A(n1226), .Y(n3124) );
  BUFX2 U3046 ( .A(n1214), .Y(n3125) );
  BUFX2 U3047 ( .A(n1202), .Y(n3126) );
  BUFX2 U3048 ( .A(n1190), .Y(n3127) );
  BUFX2 U3049 ( .A(n1178), .Y(n3128) );
  BUFX2 U3050 ( .A(n1166), .Y(n3129) );
  BUFX2 U3051 ( .A(n1154), .Y(n3130) );
  BUFX2 U3052 ( .A(n1142), .Y(n3131) );
  BUFX2 U3053 ( .A(n1130), .Y(n3132) );
  BUFX2 U3054 ( .A(n1118), .Y(n3133) );
  BUFX2 U3055 ( .A(n1106), .Y(n3134) );
  BUFX2 U3056 ( .A(n1094), .Y(n3135) );
  BUFX2 U3057 ( .A(n1082), .Y(n3136) );
  BUFX2 U3058 ( .A(n1070), .Y(n3137) );
  BUFX2 U3059 ( .A(n1058), .Y(n3138) );
  BUFX2 U3060 ( .A(n1046), .Y(n3139) );
  BUFX2 U3061 ( .A(n1034), .Y(n3140) );
  BUFX2 U3062 ( .A(n1022), .Y(n3141) );
  BUFX2 U3063 ( .A(n1010), .Y(n3142) );
  BUFX2 U3064 ( .A(n998), .Y(n3143) );
  BUFX2 U3065 ( .A(n986), .Y(n3144) );
  BUFX2 U3066 ( .A(n974), .Y(n3145) );
  BUFX2 U3067 ( .A(n962), .Y(n3146) );
  BUFX2 U3068 ( .A(n950), .Y(n3147) );
  BUFX2 U3069 ( .A(n938), .Y(n3148) );
  BUFX2 U3070 ( .A(n926), .Y(n3149) );
  BUFX2 U3071 ( .A(n914), .Y(n3150) );
  BUFX2 U3072 ( .A(n902), .Y(n3151) );
  BUFX2 U3073 ( .A(n890), .Y(n3152) );
  BUFX2 U3074 ( .A(n878), .Y(n3153) );
  BUFX2 U3075 ( .A(n866), .Y(n3154) );
  BUFX2 U3076 ( .A(n854), .Y(n3155) );
  BUFX2 U3077 ( .A(n842), .Y(n3156) );
  BUFX2 U3078 ( .A(n830), .Y(n3157) );
  BUFX2 U3079 ( .A(n818), .Y(n3158) );
  BUFX2 U3080 ( .A(n806), .Y(n3159) );
  BUFX2 U3081 ( .A(n794), .Y(n3160) );
  BUFX2 U3082 ( .A(n782), .Y(n3161) );
  BUFX2 U3083 ( .A(n770), .Y(n3162) );
  BUFX2 U3084 ( .A(n758), .Y(n3163) );
  BUFX2 U3085 ( .A(n746), .Y(n3164) );
  BUFX2 U3086 ( .A(n734), .Y(n3165) );
  BUFX2 U3087 ( .A(n722), .Y(n3166) );
  BUFX2 U3088 ( .A(n710), .Y(n3167) );
  BUFX2 U3089 ( .A(n698), .Y(n3168) );
  BUFX2 U3090 ( .A(n686), .Y(n3169) );
  BUFX2 U3091 ( .A(n674), .Y(n3170) );
  BUFX2 U3092 ( .A(n662), .Y(n3171) );
  BUFX2 U3093 ( .A(n650), .Y(n3172) );
  BUFX2 U3094 ( .A(n638), .Y(n3173) );
  BUFX2 U3095 ( .A(n626), .Y(n3174) );
  BUFX2 U3096 ( .A(n613), .Y(n3175) );
  AND2X1 U3097 ( .A(enable), .B(n3711), .Y(n2450) );
  INVX1 U3098 ( .A(n2450), .Y(n2451) );
  BUFX2 U3099 ( .A(n625), .Y(n2452) );
  INVX1 U3100 ( .A(n2452), .Y(n3183) );
  AND2X1 U3101 ( .A(n1756), .B(n3195), .Y(n2453) );
  INVX1 U3102 ( .A(n2453), .Y(n2454) );
  AND2X1 U3103 ( .A(n164), .B(n1749), .Y(n2455) );
  INVX1 U3104 ( .A(n2455), .Y(n2456) );
  AND2X1 U3105 ( .A(n2455), .B(n3183), .Y(n2457) );
  INVX1 U3106 ( .A(n2457), .Y(n2458) );
  AND2X1 U3107 ( .A(n1744), .B(n2453), .Y(n2459) );
  INVX1 U3108 ( .A(n2459), .Y(n2460) );
  AND2X1 U3109 ( .A(n3191), .B(n1749), .Y(n2461) );
  INVX1 U3110 ( .A(n2461), .Y(n2462) );
  INVX1 U3111 ( .A(n2464), .Y(n2463) );
  AND2X1 U3112 ( .A(n3196), .B(n3189), .Y(n2464) );
  AND2X1 U3113 ( .A(n3191), .B(n1748), .Y(n2465) );
  INVX1 U3114 ( .A(n2465), .Y(n2466) );
  INVX1 U3115 ( .A(n2468), .Y(n2467) );
  AND2X1 U3116 ( .A(n3191), .B(n1747), .Y(n2468) );
  AND2X1 U3117 ( .A(n3191), .B(n1746), .Y(n2469) );
  INVX1 U3118 ( .A(n2469), .Y(n2470) );
  INVX1 U3119 ( .A(n2472), .Y(n2471) );
  AND2X1 U3120 ( .A(n3191), .B(n1745), .Y(n2472) );
  AND2X1 U3121 ( .A(n3191), .B(n1744), .Y(n2473) );
  INVX1 U3122 ( .A(n2473), .Y(n2474) );
  INVX1 U3123 ( .A(n2476), .Y(n2475) );
  AND2X1 U3124 ( .A(n3191), .B(n1743), .Y(n2476) );
  AND2X1 U3125 ( .A(n3196), .B(n1749), .Y(n2477) );
  INVX1 U3126 ( .A(n2477), .Y(n2478) );
  INVX1 U3127 ( .A(n2480), .Y(n2479) );
  AND2X1 U3128 ( .A(n162), .B(n3189), .Y(n2480) );
  AND2X1 U3129 ( .A(n3196), .B(n1748), .Y(n2481) );
  INVX1 U3130 ( .A(n2481), .Y(n2482) );
  INVX1 U3131 ( .A(n2484), .Y(n2483) );
  AND2X1 U3132 ( .A(n3196), .B(n1747), .Y(n2484) );
  AND2X1 U3133 ( .A(n3196), .B(n1746), .Y(n2485) );
  INVX1 U3134 ( .A(n2485), .Y(n2486) );
  INVX1 U3135 ( .A(n2488), .Y(n2487) );
  AND2X1 U3136 ( .A(n3196), .B(n1745), .Y(n2488) );
  AND2X1 U3137 ( .A(n3196), .B(n1744), .Y(n2489) );
  INVX1 U3138 ( .A(n2489), .Y(n2490) );
  INVX1 U3139 ( .A(n2492), .Y(n2491) );
  AND2X1 U3140 ( .A(n3196), .B(n1743), .Y(n2492) );
  AND2X1 U3141 ( .A(n162), .B(n1749), .Y(n2493) );
  INVX1 U3142 ( .A(n2493), .Y(n2494) );
  AND2X1 U3143 ( .A(n164), .B(n3189), .Y(n2495) );
  INVX1 U3144 ( .A(n2495), .Y(n2496) );
  AND2X1 U3145 ( .A(n162), .B(n1748), .Y(n2497) );
  INVX1 U3146 ( .A(n2497), .Y(n2498) );
  AND2X1 U3147 ( .A(n162), .B(n1747), .Y(n2499) );
  INVX1 U3148 ( .A(n2499), .Y(n2500) );
  AND2X1 U3149 ( .A(n162), .B(n1746), .Y(n2501) );
  INVX1 U3150 ( .A(n2501), .Y(n2502) );
  AND2X1 U3151 ( .A(n162), .B(n1745), .Y(n2503) );
  INVX1 U3152 ( .A(n2503), .Y(n2504) );
  AND2X1 U3153 ( .A(n162), .B(n1744), .Y(n2505) );
  INVX1 U3154 ( .A(n2505), .Y(n2506) );
  AND2X1 U3155 ( .A(n162), .B(n1743), .Y(n2507) );
  INVX1 U3156 ( .A(n2507), .Y(n2508) );
  AND2X1 U3157 ( .A(n164), .B(n1748), .Y(n2509) );
  INVX1 U3158 ( .A(n2509), .Y(n2510) );
  AND2X1 U3159 ( .A(n164), .B(n1746), .Y(n2511) );
  INVX1 U3160 ( .A(n2511), .Y(n2512) );
  AND2X1 U3161 ( .A(n164), .B(n1745), .Y(n2513) );
  INVX1 U3162 ( .A(n2513), .Y(n2514) );
  AND2X1 U3163 ( .A(n164), .B(n1744), .Y(n2515) );
  INVX1 U3164 ( .A(n2515), .Y(n2516) );
  AND2X1 U3165 ( .A(n164), .B(n1743), .Y(n2517) );
  INVX1 U3166 ( .A(n2517), .Y(n2518) );
  AND2X1 U3167 ( .A(n3192), .B(n1749), .Y(n2519) );
  INVX1 U3168 ( .A(n2519), .Y(n2520) );
  INVX1 U3169 ( .A(n2522), .Y(n2521) );
  AND2X1 U3170 ( .A(n3194), .B(n3189), .Y(n2522) );
  AND2X1 U3171 ( .A(n3192), .B(n1748), .Y(n2523) );
  INVX1 U3172 ( .A(n2523), .Y(n2524) );
  INVX1 U3173 ( .A(n2526), .Y(n2525) );
  AND2X1 U3174 ( .A(n3192), .B(n1747), .Y(n2526) );
  AND2X1 U3175 ( .A(n3192), .B(n1746), .Y(n2527) );
  INVX1 U3176 ( .A(n2527), .Y(n2528) );
  INVX1 U3177 ( .A(n2530), .Y(n2529) );
  AND2X1 U3178 ( .A(n3192), .B(n1745), .Y(n2530) );
  AND2X1 U3179 ( .A(n3192), .B(n1744), .Y(n2531) );
  INVX1 U3180 ( .A(n2531), .Y(n2532) );
  INVX1 U3181 ( .A(n2534), .Y(n2533) );
  AND2X1 U3182 ( .A(n3192), .B(n1743), .Y(n2534) );
  INVX1 U3183 ( .A(n2536), .Y(n2535) );
  AND2X1 U3184 ( .A(n3194), .B(n1749), .Y(n2536) );
  AND2X1 U3185 ( .A(n3191), .B(n3189), .Y(n2537) );
  INVX1 U3186 ( .A(n2537), .Y(n2538) );
  AND2X1 U3187 ( .A(n3194), .B(n1748), .Y(n2539) );
  INVX1 U3188 ( .A(n2539), .Y(n2540) );
  INVX1 U3189 ( .A(n2542), .Y(n2541) );
  AND2X1 U3190 ( .A(n3194), .B(n1747), .Y(n2542) );
  AND2X1 U3191 ( .A(n3194), .B(n1746), .Y(n2543) );
  INVX1 U3192 ( .A(n2543), .Y(n2544) );
  INVX1 U3193 ( .A(n2546), .Y(n2545) );
  AND2X1 U3194 ( .A(n3194), .B(n1745), .Y(n2546) );
  AND2X1 U3195 ( .A(n3194), .B(n1744), .Y(n2547) );
  INVX1 U3196 ( .A(n2547), .Y(n2548) );
  INVX1 U3197 ( .A(n2550), .Y(n2549) );
  AND2X1 U3198 ( .A(n3194), .B(n1743), .Y(n2550) );
  AND2X1 U3199 ( .A(n1749), .B(n2453), .Y(n2551) );
  INVX1 U3200 ( .A(n2551), .Y(n2552) );
  INVX1 U3201 ( .A(n2554), .Y(n2553) );
  AND2X1 U3202 ( .A(n3193), .B(n3189), .Y(n2554) );
  AND2X1 U3203 ( .A(n1748), .B(n2453), .Y(n2555) );
  INVX1 U3204 ( .A(n2555), .Y(n2556) );
  INVX1 U3205 ( .A(n2558), .Y(n2557) );
  AND2X1 U3206 ( .A(n1747), .B(n2453), .Y(n2558) );
  AND2X1 U3207 ( .A(n1746), .B(n2453), .Y(n2559) );
  INVX1 U3208 ( .A(n2559), .Y(n2560) );
  INVX1 U3209 ( .A(n2562), .Y(n2561) );
  AND2X1 U3210 ( .A(n1745), .B(n2453), .Y(n2562) );
  INVX1 U3211 ( .A(n2564), .Y(n2563) );
  AND2X1 U3212 ( .A(n1743), .B(n2453), .Y(n2564) );
  AND2X1 U3213 ( .A(n3193), .B(n1749), .Y(n2565) );
  INVX1 U3214 ( .A(n2565), .Y(n2566) );
  INVX1 U3215 ( .A(n2568), .Y(n2567) );
  AND2X1 U3216 ( .A(n3192), .B(n3189), .Y(n2568) );
  AND2X1 U3217 ( .A(n3193), .B(n1748), .Y(n2569) );
  INVX1 U3218 ( .A(n2569), .Y(n2570) );
  INVX1 U3219 ( .A(n2572), .Y(n2571) );
  AND2X1 U3220 ( .A(n3193), .B(n1747), .Y(n2572) );
  AND2X1 U3221 ( .A(n3193), .B(n1746), .Y(n2573) );
  INVX1 U3222 ( .A(n2573), .Y(n2574) );
  INVX1 U3223 ( .A(n2576), .Y(n2575) );
  AND2X1 U3224 ( .A(n3193), .B(n1745), .Y(n2576) );
  AND2X1 U3225 ( .A(n3193), .B(n1744), .Y(n2577) );
  INVX1 U3226 ( .A(n2577), .Y(n2578) );
  INVX1 U3227 ( .A(n2580), .Y(n2579) );
  AND2X1 U3228 ( .A(n3193), .B(n1743), .Y(n2580) );
  AND2X1 U3229 ( .A(n164), .B(n1747), .Y(n2581) );
  INVX1 U3230 ( .A(n2581), .Y(n2582) );
  MUX2X1 U3231 ( .B(n2584), .A(n2585), .S(n3084), .Y(n2583) );
  MUX2X1 U3232 ( .B(n2587), .A(n2588), .S(n3089), .Y(n2586) );
  MUX2X1 U3233 ( .B(n2590), .A(n2591), .S(n3090), .Y(n2589) );
  MUX2X1 U3234 ( .B(n2593), .A(n2594), .S(n3090), .Y(n2592) );
  MUX2X1 U3235 ( .B(n2596), .A(n2597), .S(N180), .Y(n2595) );
  MUX2X1 U3236 ( .B(n2599), .A(n2600), .S(n3084), .Y(n2598) );
  MUX2X1 U3237 ( .B(n2602), .A(n2603), .S(n3084), .Y(n2601) );
  MUX2X1 U3238 ( .B(n2605), .A(n2606), .S(n3084), .Y(n2604) );
  MUX2X1 U3239 ( .B(n2608), .A(n2609), .S(n3090), .Y(n2607) );
  MUX2X1 U3240 ( .B(n2611), .A(n2612), .S(N180), .Y(n2610) );
  MUX2X1 U3241 ( .B(n2614), .A(n2615), .S(n3084), .Y(n2613) );
  MUX2X1 U3242 ( .B(n2617), .A(n2618), .S(n3084), .Y(n2616) );
  MUX2X1 U3243 ( .B(n2620), .A(n2621), .S(n3084), .Y(n2619) );
  MUX2X1 U3244 ( .B(n2623), .A(n2624), .S(n3084), .Y(n2622) );
  MUX2X1 U3245 ( .B(n2626), .A(n2627), .S(N180), .Y(n2625) );
  MUX2X1 U3246 ( .B(n2629), .A(n2630), .S(n3084), .Y(n2628) );
  MUX2X1 U3247 ( .B(n2632), .A(n2633), .S(n3084), .Y(n2631) );
  MUX2X1 U3248 ( .B(n2635), .A(n2636), .S(n3084), .Y(n2634) );
  MUX2X1 U3249 ( .B(n2638), .A(n2639), .S(n3084), .Y(n2637) );
  MUX2X1 U3250 ( .B(n2641), .A(n2642), .S(N180), .Y(n2640) );
  MUX2X1 U3251 ( .B(n2643), .A(n2644), .S(N182), .Y(N192) );
  MUX2X1 U3252 ( .B(n2646), .A(n2647), .S(n3084), .Y(n2645) );
  MUX2X1 U3253 ( .B(n2649), .A(n2650), .S(n3084), .Y(n2648) );
  MUX2X1 U3254 ( .B(n2652), .A(n2653), .S(n3084), .Y(n2651) );
  MUX2X1 U3255 ( .B(n2655), .A(n2656), .S(n3084), .Y(n2654) );
  MUX2X1 U3256 ( .B(n2658), .A(n2659), .S(N180), .Y(n2657) );
  MUX2X1 U3257 ( .B(n2661), .A(n2662), .S(n3088), .Y(n2660) );
  MUX2X1 U3258 ( .B(n2664), .A(n2665), .S(n3090), .Y(n2663) );
  MUX2X1 U3259 ( .B(n2667), .A(n2668), .S(n3088), .Y(n2666) );
  MUX2X1 U3260 ( .B(n2670), .A(n2671), .S(n3090), .Y(n2669) );
  MUX2X1 U3261 ( .B(n2673), .A(n2674), .S(N180), .Y(n2672) );
  MUX2X1 U3262 ( .B(n2676), .A(n2677), .S(n3090), .Y(n2675) );
  MUX2X1 U3263 ( .B(n2679), .A(n2680), .S(n3090), .Y(n2678) );
  MUX2X1 U3264 ( .B(n2682), .A(n2683), .S(n3084), .Y(n2681) );
  MUX2X1 U3265 ( .B(n2685), .A(n2686), .S(n3087), .Y(n2684) );
  MUX2X1 U3266 ( .B(n2688), .A(n2689), .S(N180), .Y(n2687) );
  MUX2X1 U3267 ( .B(n2691), .A(n2692), .S(n3087), .Y(n2690) );
  MUX2X1 U3268 ( .B(n2694), .A(n2695), .S(n3084), .Y(n2693) );
  MUX2X1 U3269 ( .B(n2697), .A(n2698), .S(n3089), .Y(n2696) );
  MUX2X1 U3270 ( .B(n2700), .A(n2701), .S(n3084), .Y(n2699) );
  MUX2X1 U3271 ( .B(n2703), .A(n2704), .S(N180), .Y(n2702) );
  MUX2X1 U3272 ( .B(n2705), .A(n2706), .S(N182), .Y(N191) );
  MUX2X1 U3273 ( .B(n2708), .A(n2709), .S(n3085), .Y(n2707) );
  MUX2X1 U3274 ( .B(n2711), .A(n2712), .S(n3085), .Y(n2710) );
  MUX2X1 U3275 ( .B(n2714), .A(n2715), .S(n3085), .Y(n2713) );
  MUX2X1 U3276 ( .B(n2717), .A(n2718), .S(n3085), .Y(n2716) );
  MUX2X1 U3277 ( .B(n2720), .A(n2721), .S(N180), .Y(n2719) );
  MUX2X1 U3278 ( .B(n2723), .A(n2724), .S(n3085), .Y(n2722) );
  MUX2X1 U3279 ( .B(n2726), .A(n2727), .S(n3085), .Y(n2725) );
  MUX2X1 U3280 ( .B(n2729), .A(n2730), .S(n3085), .Y(n2728) );
  MUX2X1 U3281 ( .B(n2732), .A(n2733), .S(n3085), .Y(n2731) );
  MUX2X1 U3282 ( .B(n2735), .A(n2736), .S(N180), .Y(n2734) );
  MUX2X1 U3283 ( .B(n2738), .A(n2739), .S(n3085), .Y(n2737) );
  MUX2X1 U3284 ( .B(n2741), .A(n2742), .S(n3085), .Y(n2740) );
  MUX2X1 U3285 ( .B(n2744), .A(n2745), .S(n3085), .Y(n2743) );
  MUX2X1 U3286 ( .B(n2747), .A(n2748), .S(n3085), .Y(n2746) );
  MUX2X1 U3287 ( .B(n2750), .A(n2751), .S(N180), .Y(n2749) );
  MUX2X1 U3288 ( .B(n2753), .A(n2754), .S(n3086), .Y(n2752) );
  MUX2X1 U3289 ( .B(n2756), .A(n2757), .S(n3086), .Y(n2755) );
  MUX2X1 U3290 ( .B(n2759), .A(n2760), .S(n3086), .Y(n2758) );
  MUX2X1 U3291 ( .B(n2762), .A(n2763), .S(n3086), .Y(n2761) );
  MUX2X1 U3292 ( .B(n2765), .A(n2766), .S(N180), .Y(n2764) );
  MUX2X1 U3293 ( .B(n2767), .A(n2768), .S(N182), .Y(N190) );
  MUX2X1 U3294 ( .B(n2770), .A(n2771), .S(n3086), .Y(n2769) );
  MUX2X1 U3295 ( .B(n2773), .A(n2774), .S(n3086), .Y(n2772) );
  MUX2X1 U3296 ( .B(n2776), .A(n2777), .S(n3086), .Y(n2775) );
  MUX2X1 U3297 ( .B(n2779), .A(n2780), .S(n3086), .Y(n2778) );
  MUX2X1 U3298 ( .B(n2782), .A(n2783), .S(N180), .Y(n2781) );
  MUX2X1 U3299 ( .B(n2785), .A(n2786), .S(n3086), .Y(n2784) );
  MUX2X1 U3300 ( .B(n2788), .A(n2789), .S(n3086), .Y(n2787) );
  MUX2X1 U3301 ( .B(n2791), .A(n2792), .S(n3086), .Y(n2790) );
  MUX2X1 U3302 ( .B(n2794), .A(n2795), .S(n3086), .Y(n2793) );
  MUX2X1 U3303 ( .B(n2797), .A(n2798), .S(N180), .Y(n2796) );
  MUX2X1 U3304 ( .B(n2800), .A(n2801), .S(n3085), .Y(n2799) );
  MUX2X1 U3305 ( .B(n2803), .A(n2804), .S(n3086), .Y(n2802) );
  MUX2X1 U3306 ( .B(n2806), .A(n2807), .S(n3086), .Y(n2805) );
  MUX2X1 U3307 ( .B(n2809), .A(n2810), .S(n3085), .Y(n2808) );
  MUX2X1 U3308 ( .B(n2812), .A(n2813), .S(N180), .Y(n2811) );
  MUX2X1 U3309 ( .B(n2815), .A(n2816), .S(n3085), .Y(n2814) );
  MUX2X1 U3310 ( .B(n2818), .A(n2819), .S(n3085), .Y(n2817) );
  MUX2X1 U3311 ( .B(n2821), .A(n2822), .S(n3086), .Y(n2820) );
  MUX2X1 U3312 ( .B(n2824), .A(n2825), .S(n3085), .Y(n2823) );
  MUX2X1 U3313 ( .B(n2827), .A(n2828), .S(N180), .Y(n2826) );
  MUX2X1 U3314 ( .B(n2829), .A(n2830), .S(N182), .Y(N189) );
  MUX2X1 U3315 ( .B(n2832), .A(n2833), .S(n3085), .Y(n2831) );
  MUX2X1 U3316 ( .B(n2835), .A(n2836), .S(n3085), .Y(n2834) );
  MUX2X1 U3317 ( .B(n2838), .A(n2839), .S(n3086), .Y(n2837) );
  MUX2X1 U3318 ( .B(n2841), .A(n2842), .S(n3086), .Y(n2840) );
  MUX2X1 U3319 ( .B(n2844), .A(n2845), .S(N180), .Y(n2843) );
  MUX2X1 U3320 ( .B(n2847), .A(n2848), .S(n3087), .Y(n2846) );
  MUX2X1 U3321 ( .B(n2850), .A(n2851), .S(n3087), .Y(n2849) );
  MUX2X1 U3322 ( .B(n2853), .A(n2854), .S(n3087), .Y(n2852) );
  MUX2X1 U3323 ( .B(n2856), .A(n2857), .S(n3087), .Y(n2855) );
  MUX2X1 U3324 ( .B(n2859), .A(n2860), .S(N180), .Y(n2858) );
  MUX2X1 U3325 ( .B(n2862), .A(n2863), .S(n3087), .Y(n2861) );
  MUX2X1 U3326 ( .B(n2865), .A(n2866), .S(n3087), .Y(n2864) );
  MUX2X1 U3327 ( .B(n2868), .A(n2869), .S(n3087), .Y(n2867) );
  MUX2X1 U3328 ( .B(n2871), .A(n2872), .S(n3087), .Y(n2870) );
  MUX2X1 U3329 ( .B(n2874), .A(n2875), .S(N180), .Y(n2873) );
  MUX2X1 U3330 ( .B(n2877), .A(n2878), .S(n3087), .Y(n2876) );
  MUX2X1 U3331 ( .B(n2880), .A(n2881), .S(n3087), .Y(n2879) );
  MUX2X1 U3332 ( .B(n2883), .A(n2884), .S(n3087), .Y(n2882) );
  MUX2X1 U3333 ( .B(n2886), .A(n2887), .S(n3087), .Y(n2885) );
  MUX2X1 U3334 ( .B(n2889), .A(n2890), .S(N180), .Y(n2888) );
  MUX2X1 U3335 ( .B(n2891), .A(n2892), .S(N182), .Y(N188) );
  MUX2X1 U3336 ( .B(n2894), .A(n2895), .S(n3088), .Y(n2893) );
  MUX2X1 U3337 ( .B(n2897), .A(n2898), .S(n3088), .Y(n2896) );
  MUX2X1 U3338 ( .B(n2900), .A(n2901), .S(n3088), .Y(n2899) );
  MUX2X1 U3339 ( .B(n2903), .A(n2904), .S(n3088), .Y(n2902) );
  MUX2X1 U3340 ( .B(n2906), .A(n2907), .S(N180), .Y(n2905) );
  MUX2X1 U3341 ( .B(n2909), .A(n2910), .S(n3088), .Y(n2908) );
  MUX2X1 U3342 ( .B(n2912), .A(n2913), .S(n3088), .Y(n2911) );
  MUX2X1 U3343 ( .B(n2915), .A(n2916), .S(n3088), .Y(n2914) );
  MUX2X1 U3344 ( .B(n2918), .A(n2919), .S(n3088), .Y(n2917) );
  MUX2X1 U3345 ( .B(n2921), .A(n2922), .S(N180), .Y(n2920) );
  MUX2X1 U3346 ( .B(n2924), .A(n2925), .S(n3088), .Y(n2923) );
  MUX2X1 U3347 ( .B(n2927), .A(n2928), .S(n3088), .Y(n2926) );
  MUX2X1 U3348 ( .B(n2930), .A(n2931), .S(n3088), .Y(n2929) );
  MUX2X1 U3349 ( .B(n2933), .A(n2934), .S(n3088), .Y(n2932) );
  MUX2X1 U3350 ( .B(n2936), .A(n2937), .S(N180), .Y(n2935) );
  MUX2X1 U3351 ( .B(n2939), .A(n2940), .S(n3089), .Y(n2938) );
  MUX2X1 U3352 ( .B(n2942), .A(n2943), .S(n3089), .Y(n2941) );
  MUX2X1 U3353 ( .B(n2945), .A(n2946), .S(n3089), .Y(n2944) );
  MUX2X1 U3354 ( .B(n2948), .A(n2949), .S(n3089), .Y(n2947) );
  MUX2X1 U3355 ( .B(n2951), .A(n2952), .S(N180), .Y(n2950) );
  MUX2X1 U3356 ( .B(n2953), .A(n2954), .S(N182), .Y(N187) );
  MUX2X1 U3357 ( .B(n2956), .A(n2957), .S(n3089), .Y(n2955) );
  MUX2X1 U3358 ( .B(n2959), .A(n2960), .S(n3089), .Y(n2958) );
  MUX2X1 U3359 ( .B(n2962), .A(n2963), .S(n3089), .Y(n2961) );
  MUX2X1 U3360 ( .B(n2965), .A(n2966), .S(n3089), .Y(n2964) );
  MUX2X1 U3361 ( .B(n2968), .A(n2969), .S(N180), .Y(n2967) );
  MUX2X1 U3362 ( .B(n2971), .A(n2972), .S(n3089), .Y(n2970) );
  MUX2X1 U3363 ( .B(n2974), .A(n2975), .S(n3089), .Y(n2973) );
  MUX2X1 U3364 ( .B(n2977), .A(n2978), .S(n3089), .Y(n2976) );
  MUX2X1 U3365 ( .B(n2980), .A(n2981), .S(n3089), .Y(n2979) );
  MUX2X1 U3366 ( .B(n2983), .A(n2984), .S(N180), .Y(n2982) );
  MUX2X1 U3367 ( .B(n2986), .A(n2987), .S(n3088), .Y(n2985) );
  MUX2X1 U3368 ( .B(n2989), .A(n2990), .S(n3088), .Y(n2988) );
  MUX2X1 U3369 ( .B(n2992), .A(n2993), .S(n3089), .Y(n2991) );
  MUX2X1 U3370 ( .B(n2995), .A(n2996), .S(n3088), .Y(n2994) );
  MUX2X1 U3371 ( .B(n2998), .A(n2999), .S(N180), .Y(n2997) );
  MUX2X1 U3372 ( .B(n3001), .A(n3002), .S(n3089), .Y(n3000) );
  MUX2X1 U3373 ( .B(n3004), .A(n3005), .S(n3088), .Y(n3003) );
  MUX2X1 U3374 ( .B(n3007), .A(n3008), .S(n3087), .Y(n3006) );
  MUX2X1 U3375 ( .B(n3010), .A(n3011), .S(n3087), .Y(n3009) );
  MUX2X1 U3376 ( .B(n3013), .A(n3014), .S(N180), .Y(n3012) );
  MUX2X1 U3377 ( .B(n3015), .A(n3016), .S(N182), .Y(N186) );
  MUX2X1 U3378 ( .B(n3018), .A(n3019), .S(n3089), .Y(n3017) );
  MUX2X1 U3379 ( .B(n3021), .A(n3022), .S(n3089), .Y(n3020) );
  MUX2X1 U3380 ( .B(n3024), .A(n3025), .S(n3087), .Y(n3023) );
  MUX2X1 U3381 ( .B(n3027), .A(n3028), .S(n3087), .Y(n3026) );
  MUX2X1 U3382 ( .B(n3030), .A(n3031), .S(N180), .Y(n3029) );
  MUX2X1 U3383 ( .B(n3033), .A(n3034), .S(n3090), .Y(n3032) );
  MUX2X1 U3384 ( .B(n3036), .A(n3037), .S(n3090), .Y(n3035) );
  MUX2X1 U3385 ( .B(n3039), .A(n3040), .S(n3090), .Y(n3038) );
  MUX2X1 U3386 ( .B(n3042), .A(n3043), .S(n3090), .Y(n3041) );
  MUX2X1 U3387 ( .B(n3045), .A(n3046), .S(N180), .Y(n3044) );
  MUX2X1 U3388 ( .B(n3048), .A(n3049), .S(n3090), .Y(n3047) );
  MUX2X1 U3389 ( .B(n3051), .A(n3052), .S(n3090), .Y(n3050) );
  MUX2X1 U3390 ( .B(n3054), .A(n3055), .S(n3090), .Y(n3053) );
  MUX2X1 U3391 ( .B(n3057), .A(n3058), .S(n3090), .Y(n3056) );
  MUX2X1 U3392 ( .B(n3060), .A(n3061), .S(N180), .Y(n3059) );
  MUX2X1 U3393 ( .B(n3063), .A(n3064), .S(n3090), .Y(n3062) );
  MUX2X1 U3394 ( .B(n3066), .A(n3067), .S(n3090), .Y(n3065) );
  MUX2X1 U3395 ( .B(n3069), .A(n3070), .S(n3090), .Y(n3068) );
  MUX2X1 U3396 ( .B(n3072), .A(n3073), .S(n3090), .Y(n3071) );
  MUX2X1 U3397 ( .B(n3075), .A(n3076), .S(N180), .Y(n3074) );
  MUX2X1 U3398 ( .B(n3077), .A(n3078), .S(N182), .Y(N185) );
  MUX2X1 U3399 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n3096), .Y(n2585) );
  MUX2X1 U3400 ( .B(\mem<60><0> ), .A(\mem<61><0> ), .S(n3095), .Y(n2584) );
  MUX2X1 U3401 ( .B(\mem<58><0> ), .A(\mem<59><0> ), .S(n3096), .Y(n2588) );
  MUX2X1 U3402 ( .B(\mem<56><0> ), .A(\mem<57><0> ), .S(n3095), .Y(n2587) );
  MUX2X1 U3403 ( .B(n2586), .A(n2583), .S(n3083), .Y(n2597) );
  MUX2X1 U3404 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n3095), .Y(n2591) );
  MUX2X1 U3405 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n3095), .Y(n2590) );
  MUX2X1 U3406 ( .B(\mem<50><0> ), .A(\mem<51><0> ), .S(n3095), .Y(n2594) );
  MUX2X1 U3407 ( .B(\mem<48><0> ), .A(\mem<49><0> ), .S(n3095), .Y(n2593) );
  MUX2X1 U3408 ( .B(n2592), .A(n2589), .S(n3083), .Y(n2596) );
  MUX2X1 U3409 ( .B(\mem<46><0> ), .A(\mem<47><0> ), .S(n3095), .Y(n2600) );
  MUX2X1 U3410 ( .B(\mem<44><0> ), .A(\mem<45><0> ), .S(n3095), .Y(n2599) );
  MUX2X1 U3411 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n3095), .Y(n2603) );
  MUX2X1 U3412 ( .B(\mem<40><0> ), .A(\mem<41><0> ), .S(n3095), .Y(n2602) );
  MUX2X1 U3413 ( .B(n2601), .A(n2598), .S(n3083), .Y(n2612) );
  MUX2X1 U3414 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n3095), .Y(n2606) );
  MUX2X1 U3415 ( .B(\mem<36><0> ), .A(\mem<37><0> ), .S(n3095), .Y(n2605) );
  MUX2X1 U3416 ( .B(\mem<34><0> ), .A(\mem<35><0> ), .S(n3095), .Y(n2609) );
  MUX2X1 U3417 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n3095), .Y(n2608) );
  MUX2X1 U3418 ( .B(n2607), .A(n2604), .S(n3083), .Y(n2611) );
  MUX2X1 U3419 ( .B(n2610), .A(n2595), .S(N181), .Y(n2644) );
  MUX2X1 U3420 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n3096), .Y(n2615) );
  MUX2X1 U3421 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n3096), .Y(n2614) );
  MUX2X1 U3422 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n3096), .Y(n2618) );
  MUX2X1 U3423 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n3096), .Y(n2617) );
  MUX2X1 U3424 ( .B(n2616), .A(n2613), .S(n3083), .Y(n2627) );
  MUX2X1 U3425 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n3096), .Y(n2621) );
  MUX2X1 U3426 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n3096), .Y(n2620) );
  MUX2X1 U3427 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n3096), .Y(n2624) );
  MUX2X1 U3428 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n3096), .Y(n2623) );
  MUX2X1 U3429 ( .B(n2622), .A(n2619), .S(n3083), .Y(n2626) );
  MUX2X1 U3430 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n3096), .Y(n2630) );
  MUX2X1 U3431 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n3096), .Y(n2629) );
  MUX2X1 U3432 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n3096), .Y(n2633) );
  MUX2X1 U3433 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n3096), .Y(n2632) );
  MUX2X1 U3434 ( .B(n2631), .A(n2628), .S(n3083), .Y(n2642) );
  MUX2X1 U3435 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n3097), .Y(n2636) );
  MUX2X1 U3436 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n3097), .Y(n2635) );
  MUX2X1 U3437 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n3097), .Y(n2639) );
  MUX2X1 U3438 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n3097), .Y(n2638) );
  MUX2X1 U3439 ( .B(n2637), .A(n2634), .S(n3083), .Y(n2641) );
  MUX2X1 U3440 ( .B(n2640), .A(n2625), .S(N181), .Y(n2643) );
  MUX2X1 U3441 ( .B(\mem<62><1> ), .A(\mem<63><1> ), .S(n3097), .Y(n2647) );
  MUX2X1 U3442 ( .B(\mem<60><1> ), .A(\mem<61><1> ), .S(n3097), .Y(n2646) );
  MUX2X1 U3443 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n3097), .Y(n2650) );
  MUX2X1 U3444 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n3097), .Y(n2649) );
  MUX2X1 U3445 ( .B(n2648), .A(n2645), .S(n3083), .Y(n2659) );
  MUX2X1 U3446 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n3097), .Y(n2653) );
  MUX2X1 U3447 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n3097), .Y(n2652) );
  MUX2X1 U3448 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n3097), .Y(n2656) );
  MUX2X1 U3449 ( .B(\mem<48><1> ), .A(\mem<49><1> ), .S(n3097), .Y(n2655) );
  MUX2X1 U3450 ( .B(n2654), .A(n2651), .S(n3083), .Y(n2658) );
  MUX2X1 U3451 ( .B(\mem<46><1> ), .A(\mem<47><1> ), .S(n3098), .Y(n2662) );
  MUX2X1 U3452 ( .B(\mem<44><1> ), .A(\mem<45><1> ), .S(n3098), .Y(n2661) );
  MUX2X1 U3453 ( .B(\mem<42><1> ), .A(\mem<43><1> ), .S(n3098), .Y(n2665) );
  MUX2X1 U3454 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n3098), .Y(n2664) );
  MUX2X1 U3455 ( .B(n2663), .A(n2660), .S(n3083), .Y(n2674) );
  MUX2X1 U3456 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n3098), .Y(n2668) );
  MUX2X1 U3457 ( .B(\mem<36><1> ), .A(\mem<37><1> ), .S(n3098), .Y(n2667) );
  MUX2X1 U3458 ( .B(\mem<34><1> ), .A(\mem<35><1> ), .S(n3098), .Y(n2671) );
  MUX2X1 U3459 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n3098), .Y(n2670) );
  MUX2X1 U3460 ( .B(n2669), .A(n2666), .S(n3083), .Y(n2673) );
  MUX2X1 U3461 ( .B(n2672), .A(n2657), .S(N181), .Y(n2706) );
  MUX2X1 U3462 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n3098), .Y(n2677) );
  MUX2X1 U3463 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n3098), .Y(n2676) );
  MUX2X1 U3464 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n3098), .Y(n2680) );
  MUX2X1 U3465 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n3098), .Y(n2679) );
  MUX2X1 U3466 ( .B(n2678), .A(n2675), .S(n3082), .Y(n2689) );
  MUX2X1 U3467 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n3099), .Y(n2683) );
  MUX2X1 U3468 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n3099), .Y(n2682) );
  MUX2X1 U3469 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n3099), .Y(n2686) );
  MUX2X1 U3470 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n3099), .Y(n2685) );
  MUX2X1 U3471 ( .B(n2684), .A(n2681), .S(n3082), .Y(n2688) );
  MUX2X1 U3472 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n3099), .Y(n2692) );
  MUX2X1 U3473 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n3099), .Y(n2691) );
  MUX2X1 U3474 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n3099), .Y(n2695) );
  MUX2X1 U3475 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n3099), .Y(n2694) );
  MUX2X1 U3476 ( .B(n2693), .A(n2690), .S(n3082), .Y(n2704) );
  MUX2X1 U3477 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n3099), .Y(n2698) );
  MUX2X1 U3478 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n3099), .Y(n2697) );
  MUX2X1 U3479 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n3099), .Y(n2701) );
  MUX2X1 U3480 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n3099), .Y(n2700) );
  MUX2X1 U3481 ( .B(n2699), .A(n2696), .S(n3082), .Y(n2703) );
  MUX2X1 U3482 ( .B(n2702), .A(n2687), .S(N181), .Y(n2705) );
  MUX2X1 U3483 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n3100), .Y(n2709) );
  MUX2X1 U3484 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n3100), .Y(n2708) );
  MUX2X1 U3485 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n3100), .Y(n2712) );
  MUX2X1 U3486 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n3100), .Y(n2711) );
  MUX2X1 U3487 ( .B(n2710), .A(n2707), .S(n3082), .Y(n2721) );
  MUX2X1 U3488 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n3100), .Y(n2715) );
  MUX2X1 U3489 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n3100), .Y(n2714) );
  MUX2X1 U3490 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n3100), .Y(n2718) );
  MUX2X1 U3491 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n3100), .Y(n2717) );
  MUX2X1 U3492 ( .B(n2716), .A(n2713), .S(n3082), .Y(n2720) );
  MUX2X1 U3493 ( .B(\mem<46><2> ), .A(\mem<47><2> ), .S(n3100), .Y(n2724) );
  MUX2X1 U3494 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n3100), .Y(n2723) );
  MUX2X1 U3495 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n3100), .Y(n2727) );
  MUX2X1 U3496 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n3100), .Y(n2726) );
  MUX2X1 U3497 ( .B(n2725), .A(n2722), .S(n3082), .Y(n2736) );
  MUX2X1 U3498 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n3101), .Y(n2730) );
  MUX2X1 U3499 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n3101), .Y(n2729) );
  MUX2X1 U3500 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n3101), .Y(n2733) );
  MUX2X1 U3501 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n3101), .Y(n2732) );
  MUX2X1 U3502 ( .B(n2731), .A(n2728), .S(n3082), .Y(n2735) );
  MUX2X1 U3503 ( .B(n2734), .A(n2719), .S(N181), .Y(n2768) );
  MUX2X1 U3504 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n3101), .Y(n2739) );
  MUX2X1 U3505 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n3101), .Y(n2738) );
  MUX2X1 U3506 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n3101), .Y(n2742) );
  MUX2X1 U3507 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n3101), .Y(n2741) );
  MUX2X1 U3508 ( .B(n2740), .A(n2737), .S(n3082), .Y(n2751) );
  MUX2X1 U3509 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n3101), .Y(n2745) );
  MUX2X1 U3510 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n3101), .Y(n2744) );
  MUX2X1 U3511 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n3101), .Y(n2748) );
  MUX2X1 U3512 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n3101), .Y(n2747) );
  MUX2X1 U3513 ( .B(n2746), .A(n2743), .S(n3082), .Y(n2750) );
  MUX2X1 U3514 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n3097), .Y(n2754) );
  MUX2X1 U3515 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n3099), .Y(n2753) );
  MUX2X1 U3516 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n3097), .Y(n2757) );
  MUX2X1 U3517 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n3097), .Y(n2756) );
  MUX2X1 U3518 ( .B(n2755), .A(n2752), .S(n3082), .Y(n2766) );
  MUX2X1 U3519 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n3097), .Y(n2760) );
  MUX2X1 U3520 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n3099), .Y(n2759) );
  MUX2X1 U3521 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n3097), .Y(n2763) );
  MUX2X1 U3522 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n3097), .Y(n2762) );
  MUX2X1 U3523 ( .B(n2761), .A(n2758), .S(n3082), .Y(n2765) );
  MUX2X1 U3524 ( .B(n2764), .A(n2749), .S(N181), .Y(n2767) );
  MUX2X1 U3525 ( .B(\mem<62><3> ), .A(\mem<63><3> ), .S(n3098), .Y(n2771) );
  MUX2X1 U3526 ( .B(\mem<60><3> ), .A(\mem<61><3> ), .S(n3099), .Y(n2770) );
  MUX2X1 U3527 ( .B(\mem<58><3> ), .A(\mem<59><3> ), .S(n3100), .Y(n2774) );
  MUX2X1 U3528 ( .B(\mem<56><3> ), .A(\mem<57><3> ), .S(n3101), .Y(n2773) );
  MUX2X1 U3529 ( .B(n2772), .A(n2769), .S(n3083), .Y(n2783) );
  MUX2X1 U3530 ( .B(\mem<54><3> ), .A(\mem<55><3> ), .S(n3102), .Y(n2777) );
  MUX2X1 U3531 ( .B(\mem<52><3> ), .A(\mem<53><3> ), .S(n3102), .Y(n2776) );
  MUX2X1 U3532 ( .B(\mem<50><3> ), .A(\mem<51><3> ), .S(n3102), .Y(n2780) );
  MUX2X1 U3533 ( .B(\mem<48><3> ), .A(\mem<49><3> ), .S(n3102), .Y(n2779) );
  MUX2X1 U3534 ( .B(n2778), .A(n2775), .S(n3082), .Y(n2782) );
  MUX2X1 U3535 ( .B(\mem<46><3> ), .A(\mem<47><3> ), .S(n3102), .Y(n2786) );
  MUX2X1 U3536 ( .B(\mem<44><3> ), .A(\mem<45><3> ), .S(n3102), .Y(n2785) );
  MUX2X1 U3537 ( .B(\mem<42><3> ), .A(\mem<43><3> ), .S(n3102), .Y(n2789) );
  MUX2X1 U3538 ( .B(\mem<40><3> ), .A(\mem<41><3> ), .S(n3102), .Y(n2788) );
  MUX2X1 U3539 ( .B(n2787), .A(n2784), .S(n3083), .Y(n2798) );
  MUX2X1 U3540 ( .B(\mem<38><3> ), .A(\mem<39><3> ), .S(n3102), .Y(n2792) );
  MUX2X1 U3541 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n3102), .Y(n2791) );
  MUX2X1 U3542 ( .B(\mem<34><3> ), .A(\mem<35><3> ), .S(n3102), .Y(n2795) );
  MUX2X1 U3543 ( .B(\mem<32><3> ), .A(\mem<33><3> ), .S(n3102), .Y(n2794) );
  MUX2X1 U3544 ( .B(n2793), .A(n2790), .S(n3082), .Y(n2797) );
  MUX2X1 U3545 ( .B(n2796), .A(n2781), .S(N181), .Y(n2830) );
  MUX2X1 U3546 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n3103), .Y(n2801) );
  MUX2X1 U3547 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n3103), .Y(n2800) );
  MUX2X1 U3548 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n3103), .Y(n2804) );
  MUX2X1 U3549 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n3103), .Y(n2803) );
  MUX2X1 U3550 ( .B(n2802), .A(n2799), .S(n3083), .Y(n2813) );
  MUX2X1 U3551 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n3103), .Y(n2807) );
  MUX2X1 U3552 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n3103), .Y(n2806) );
  MUX2X1 U3553 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n3103), .Y(n2810) );
  MUX2X1 U3554 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n3103), .Y(n2809) );
  MUX2X1 U3555 ( .B(n2808), .A(n2805), .S(n3082), .Y(n2812) );
  MUX2X1 U3556 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n3103), .Y(n2816) );
  MUX2X1 U3557 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n3103), .Y(n2815) );
  MUX2X1 U3558 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n3103), .Y(n2819) );
  MUX2X1 U3559 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n3103), .Y(n2818) );
  MUX2X1 U3560 ( .B(n2817), .A(n2814), .S(n3082), .Y(n2828) );
  MUX2X1 U3561 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n3099), .Y(n2822) );
  MUX2X1 U3562 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n3097), .Y(n2821) );
  MUX2X1 U3563 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n3099), .Y(n2825) );
  MUX2X1 U3564 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n3097), .Y(n2824) );
  MUX2X1 U3565 ( .B(n2823), .A(n2820), .S(n3082), .Y(n2827) );
  MUX2X1 U3566 ( .B(n2826), .A(n2811), .S(N181), .Y(n2829) );
  MUX2X1 U3567 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n3099), .Y(n2833) );
  MUX2X1 U3568 ( .B(\mem<60><4> ), .A(\mem<61><4> ), .S(n3097), .Y(n2832) );
  MUX2X1 U3569 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n3099), .Y(n2836) );
  MUX2X1 U3570 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n3097), .Y(n2835) );
  MUX2X1 U3571 ( .B(n2834), .A(n2831), .S(n3083), .Y(n2845) );
  MUX2X1 U3572 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n3099), .Y(n2839) );
  MUX2X1 U3573 ( .B(\mem<52><4> ), .A(\mem<53><4> ), .S(n3097), .Y(n2838) );
  MUX2X1 U3574 ( .B(\mem<50><4> ), .A(\mem<51><4> ), .S(n3099), .Y(n2842) );
  MUX2X1 U3575 ( .B(\mem<48><4> ), .A(\mem<49><4> ), .S(n3097), .Y(n2841) );
  MUX2X1 U3576 ( .B(n2840), .A(n2837), .S(n3082), .Y(n2844) );
  MUX2X1 U3577 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n3104), .Y(n2848) );
  MUX2X1 U3578 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n3104), .Y(n2847) );
  MUX2X1 U3579 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n3104), .Y(n2851) );
  MUX2X1 U3580 ( .B(\mem<40><4> ), .A(\mem<41><4> ), .S(n3104), .Y(n2850) );
  MUX2X1 U3581 ( .B(n2849), .A(n2846), .S(n3083), .Y(n2860) );
  MUX2X1 U3582 ( .B(\mem<38><4> ), .A(\mem<39><4> ), .S(n3104), .Y(n2854) );
  MUX2X1 U3583 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n3104), .Y(n2853) );
  MUX2X1 U3584 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n3104), .Y(n2857) );
  MUX2X1 U3585 ( .B(\mem<32><4> ), .A(\mem<33><4> ), .S(n3104), .Y(n2856) );
  MUX2X1 U3586 ( .B(n2855), .A(n2852), .S(n3082), .Y(n2859) );
  MUX2X1 U3587 ( .B(n2858), .A(n2843), .S(N181), .Y(n2892) );
  MUX2X1 U3588 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n3104), .Y(n2863) );
  MUX2X1 U3589 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n3104), .Y(n2862) );
  MUX2X1 U3590 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n3104), .Y(n2866) );
  MUX2X1 U3591 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n3104), .Y(n2865) );
  MUX2X1 U3592 ( .B(n2864), .A(n2861), .S(n3081), .Y(n2875) );
  MUX2X1 U3593 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n3105), .Y(n2869) );
  MUX2X1 U3594 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n3105), .Y(n2868) );
  MUX2X1 U3595 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n3105), .Y(n2872) );
  MUX2X1 U3596 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n3105), .Y(n2871) );
  MUX2X1 U3597 ( .B(n2870), .A(n2867), .S(n3081), .Y(n2874) );
  MUX2X1 U3598 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n3105), .Y(n2878) );
  MUX2X1 U3599 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n3105), .Y(n2877) );
  MUX2X1 U3600 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n3105), .Y(n2881) );
  MUX2X1 U3601 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n3105), .Y(n2880) );
  MUX2X1 U3602 ( .B(n2879), .A(n2876), .S(n3081), .Y(n2890) );
  MUX2X1 U3603 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n3105), .Y(n2884) );
  MUX2X1 U3604 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n3105), .Y(n2883) );
  MUX2X1 U3605 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n3105), .Y(n2887) );
  MUX2X1 U3606 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n3105), .Y(n2886) );
  MUX2X1 U3607 ( .B(n2885), .A(n2882), .S(n3081), .Y(n2889) );
  MUX2X1 U3608 ( .B(n2888), .A(n2873), .S(N181), .Y(n2891) );
  MUX2X1 U3609 ( .B(\mem<62><5> ), .A(\mem<63><5> ), .S(n3106), .Y(n2895) );
  MUX2X1 U3610 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n3106), .Y(n2894) );
  MUX2X1 U3611 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n3106), .Y(n2898) );
  MUX2X1 U3612 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n3106), .Y(n2897) );
  MUX2X1 U3613 ( .B(n2896), .A(n2893), .S(n3081), .Y(n2907) );
  MUX2X1 U3614 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n3106), .Y(n2901) );
  MUX2X1 U3615 ( .B(\mem<52><5> ), .A(\mem<53><5> ), .S(n3106), .Y(n2900) );
  MUX2X1 U3616 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n3106), .Y(n2904) );
  MUX2X1 U3617 ( .B(\mem<48><5> ), .A(\mem<49><5> ), .S(n3106), .Y(n2903) );
  MUX2X1 U3618 ( .B(n2902), .A(n2899), .S(n3081), .Y(n2906) );
  MUX2X1 U3619 ( .B(\mem<46><5> ), .A(\mem<47><5> ), .S(n3106), .Y(n2910) );
  MUX2X1 U3620 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n3106), .Y(n2909) );
  MUX2X1 U3621 ( .B(\mem<42><5> ), .A(\mem<43><5> ), .S(n3106), .Y(n2913) );
  MUX2X1 U3622 ( .B(\mem<40><5> ), .A(\mem<41><5> ), .S(n3106), .Y(n2912) );
  MUX2X1 U3623 ( .B(n2911), .A(n2908), .S(n3081), .Y(n2922) );
  MUX2X1 U3624 ( .B(\mem<38><5> ), .A(\mem<39><5> ), .S(n3107), .Y(n2916) );
  MUX2X1 U3625 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n3107), .Y(n2915) );
  MUX2X1 U3626 ( .B(\mem<34><5> ), .A(\mem<35><5> ), .S(n3107), .Y(n2919) );
  MUX2X1 U3627 ( .B(\mem<32><5> ), .A(\mem<33><5> ), .S(n3107), .Y(n2918) );
  MUX2X1 U3628 ( .B(n2917), .A(n2914), .S(n3081), .Y(n2921) );
  MUX2X1 U3629 ( .B(n2920), .A(n2905), .S(N181), .Y(n2954) );
  MUX2X1 U3630 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n3107), .Y(n2925) );
  MUX2X1 U3631 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n3107), .Y(n2924) );
  MUX2X1 U3632 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n3107), .Y(n2928) );
  MUX2X1 U3633 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n3107), .Y(n2927) );
  MUX2X1 U3634 ( .B(n2926), .A(n2923), .S(n3081), .Y(n2937) );
  MUX2X1 U3635 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n3107), .Y(n2931) );
  MUX2X1 U3636 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n3107), .Y(n2930) );
  MUX2X1 U3637 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n3107), .Y(n2934) );
  MUX2X1 U3638 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n3107), .Y(n2933) );
  MUX2X1 U3639 ( .B(n2932), .A(n2929), .S(n3081), .Y(n2936) );
  MUX2X1 U3640 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n3108), .Y(n2940) );
  MUX2X1 U3641 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n3108), .Y(n2939) );
  MUX2X1 U3642 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n3108), .Y(n2943) );
  MUX2X1 U3643 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n3108), .Y(n2942) );
  MUX2X1 U3644 ( .B(n2941), .A(n2938), .S(n3081), .Y(n2952) );
  MUX2X1 U3645 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n3108), .Y(n2946) );
  MUX2X1 U3646 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n3108), .Y(n2945) );
  MUX2X1 U3647 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n3108), .Y(n2949) );
  MUX2X1 U3648 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n3108), .Y(n2948) );
  MUX2X1 U3649 ( .B(n2947), .A(n2944), .S(n3081), .Y(n2951) );
  MUX2X1 U3650 ( .B(n2950), .A(n2935), .S(N181), .Y(n2953) );
  MUX2X1 U3651 ( .B(\mem<62><6> ), .A(\mem<63><6> ), .S(n3108), .Y(n2957) );
  MUX2X1 U3652 ( .B(\mem<60><6> ), .A(\mem<61><6> ), .S(n3108), .Y(n2956) );
  MUX2X1 U3653 ( .B(\mem<58><6> ), .A(\mem<59><6> ), .S(n3108), .Y(n2960) );
  MUX2X1 U3654 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n3108), .Y(n2959) );
  MUX2X1 U3655 ( .B(n2958), .A(n2955), .S(n3080), .Y(n2969) );
  MUX2X1 U3656 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n3109), .Y(n2963) );
  MUX2X1 U3657 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n3109), .Y(n2962) );
  MUX2X1 U3658 ( .B(\mem<50><6> ), .A(\mem<51><6> ), .S(n3109), .Y(n2966) );
  MUX2X1 U3659 ( .B(\mem<48><6> ), .A(\mem<49><6> ), .S(n3109), .Y(n2965) );
  MUX2X1 U3660 ( .B(n2964), .A(n2961), .S(n3080), .Y(n2968) );
  MUX2X1 U3661 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n3109), .Y(n2972) );
  MUX2X1 U3662 ( .B(\mem<44><6> ), .A(\mem<45><6> ), .S(n3109), .Y(n2971) );
  MUX2X1 U3663 ( .B(\mem<42><6> ), .A(\mem<43><6> ), .S(n3109), .Y(n2975) );
  MUX2X1 U3664 ( .B(\mem<40><6> ), .A(\mem<41><6> ), .S(n3109), .Y(n2974) );
  MUX2X1 U3665 ( .B(n2973), .A(n2970), .S(n3080), .Y(n2984) );
  MUX2X1 U3666 ( .B(\mem<38><6> ), .A(\mem<39><6> ), .S(n3109), .Y(n2978) );
  MUX2X1 U3667 ( .B(\mem<36><6> ), .A(\mem<37><6> ), .S(n3109), .Y(n2977) );
  MUX2X1 U3668 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n3109), .Y(n2981) );
  MUX2X1 U3669 ( .B(\mem<32><6> ), .A(\mem<33><6> ), .S(n3109), .Y(n2980) );
  MUX2X1 U3670 ( .B(n2979), .A(n2976), .S(n3080), .Y(n2983) );
  MUX2X1 U3671 ( .B(n2982), .A(n2967), .S(N181), .Y(n3016) );
  MUX2X1 U3672 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n3110), .Y(n2987) );
  MUX2X1 U3673 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n3110), .Y(n2986) );
  MUX2X1 U3674 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n3110), .Y(n2990) );
  MUX2X1 U3675 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n3110), .Y(n2989) );
  MUX2X1 U3676 ( .B(n2988), .A(n2985), .S(n3080), .Y(n2999) );
  MUX2X1 U3677 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n3110), .Y(n2993) );
  MUX2X1 U3678 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n3110), .Y(n2992) );
  MUX2X1 U3679 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n3110), .Y(n2996) );
  MUX2X1 U3680 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n3110), .Y(n2995) );
  MUX2X1 U3681 ( .B(n2994), .A(n2991), .S(n3080), .Y(n2998) );
  MUX2X1 U3682 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n3110), .Y(n3002) );
  MUX2X1 U3683 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n3110), .Y(n3001) );
  MUX2X1 U3684 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n3110), .Y(n3005) );
  MUX2X1 U3685 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n3110), .Y(n3004) );
  MUX2X1 U3686 ( .B(n3003), .A(n3000), .S(n3080), .Y(n3014) );
  MUX2X1 U3687 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n3111), .Y(n3008) );
  MUX2X1 U3688 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n3111), .Y(n3007) );
  MUX2X1 U3689 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n3111), .Y(n3011) );
  MUX2X1 U3690 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n3111), .Y(n3010) );
  MUX2X1 U3691 ( .B(n3009), .A(n3006), .S(n3080), .Y(n3013) );
  MUX2X1 U3692 ( .B(n3012), .A(n2997), .S(N181), .Y(n3015) );
  MUX2X1 U3693 ( .B(\mem<62><7> ), .A(\mem<63><7> ), .S(n3111), .Y(n3019) );
  MUX2X1 U3694 ( .B(\mem<60><7> ), .A(\mem<61><7> ), .S(n3111), .Y(n3018) );
  MUX2X1 U3695 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n3111), .Y(n3022) );
  MUX2X1 U3696 ( .B(\mem<56><7> ), .A(\mem<57><7> ), .S(n3111), .Y(n3021) );
  MUX2X1 U3697 ( .B(n3020), .A(n3017), .S(n3080), .Y(n3031) );
  MUX2X1 U3698 ( .B(\mem<54><7> ), .A(\mem<55><7> ), .S(n3111), .Y(n3025) );
  MUX2X1 U3699 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n3111), .Y(n3024) );
  MUX2X1 U3700 ( .B(\mem<50><7> ), .A(\mem<51><7> ), .S(n3111), .Y(n3028) );
  MUX2X1 U3701 ( .B(\mem<48><7> ), .A(\mem<49><7> ), .S(n3111), .Y(n3027) );
  MUX2X1 U3702 ( .B(n3026), .A(n3023), .S(n3080), .Y(n3030) );
  MUX2X1 U3703 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n3112), .Y(n3034) );
  MUX2X1 U3704 ( .B(\mem<44><7> ), .A(\mem<45><7> ), .S(n3112), .Y(n3033) );
  MUX2X1 U3705 ( .B(\mem<42><7> ), .A(\mem<43><7> ), .S(n3112), .Y(n3037) );
  MUX2X1 U3706 ( .B(\mem<40><7> ), .A(\mem<41><7> ), .S(n3112), .Y(n3036) );
  MUX2X1 U3707 ( .B(n3035), .A(n3032), .S(n3080), .Y(n3046) );
  MUX2X1 U3708 ( .B(\mem<38><7> ), .A(\mem<39><7> ), .S(n3112), .Y(n3040) );
  MUX2X1 U3709 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n3112), .Y(n3039) );
  MUX2X1 U3710 ( .B(\mem<34><7> ), .A(\mem<35><7> ), .S(n3112), .Y(n3043) );
  MUX2X1 U3711 ( .B(\mem<32><7> ), .A(\mem<33><7> ), .S(n3112), .Y(n3042) );
  MUX2X1 U3712 ( .B(n3041), .A(n3038), .S(n3080), .Y(n3045) );
  MUX2X1 U3713 ( .B(n3044), .A(n3029), .S(N181), .Y(n3078) );
  MUX2X1 U3714 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n3112), .Y(n3049) );
  MUX2X1 U3715 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n3112), .Y(n3048) );
  MUX2X1 U3716 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n3112), .Y(n3052) );
  MUX2X1 U3717 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n3112), .Y(n3051) );
  MUX2X1 U3718 ( .B(n3050), .A(n3047), .S(n3081), .Y(n3061) );
  MUX2X1 U3719 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n3096), .Y(n3055) );
  MUX2X1 U3720 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n3095), .Y(n3054) );
  MUX2X1 U3721 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n3095), .Y(n3058) );
  MUX2X1 U3722 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n3095), .Y(n3057) );
  MUX2X1 U3723 ( .B(n3056), .A(n3053), .S(n3080), .Y(n3060) );
  MUX2X1 U3724 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n3096), .Y(n3064) );
  MUX2X1 U3725 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n3096), .Y(n3063) );
  MUX2X1 U3726 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n3095), .Y(n3067) );
  MUX2X1 U3727 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n3096), .Y(n3066) );
  MUX2X1 U3728 ( .B(n3065), .A(n3062), .S(n3081), .Y(n3076) );
  MUX2X1 U3729 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n3095), .Y(n3070) );
  MUX2X1 U3730 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n3096), .Y(n3069) );
  MUX2X1 U3731 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n3096), .Y(n3073) );
  MUX2X1 U3732 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n3096), .Y(n3072) );
  MUX2X1 U3733 ( .B(n3071), .A(n3068), .S(n3080), .Y(n3075) );
  MUX2X1 U3734 ( .B(n3074), .A(n3059), .S(N181), .Y(n3077) );
  INVX8 U3735 ( .A(n3183), .Y(n3176) );
  INVX8 U3736 ( .A(n3180), .Y(n3177) );
  INVX4 U3737 ( .A(n2452), .Y(n3180) );
endmodule


module cla16_2 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n5,
         n6, n7, n8, n1, n2, n4, n9, n10;

  AOI21X1 U5 ( .A(\P<3> ), .B(n4), .C(\G<3> ), .Y(n5) );
  AOI21X1 U6 ( .A(\P<2> ), .B(n9), .C(\G<2> ), .Y(n6) );
  AOI21X1 U7 ( .A(\P<1> ), .B(n10), .C(\G<1> ), .Y(n7) );
  AOI21X1 U8 ( .A(\P<0> ), .B(Cin), .C(\G<0> ), .Y(n8) );
  cla4_11 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_10 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n10), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_9 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n9), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_8 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n4), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  BUFX2 U1 ( .A(n7), .Y(n1) );
  INVX1 U2 ( .A(n6), .Y(n4) );
  INVX1 U3 ( .A(n8), .Y(n10) );
  BUFX2 U4 ( .A(n5), .Y(n2) );
  INVX1 U9 ( .A(n2), .Y(Cout) );
  INVX2 U10 ( .A(n1), .Y(n9) );
endmodule


module dff_355 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_356 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_357 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_358 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_359 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_360 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_361 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_362 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_363 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_364 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_365 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_366 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_367 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_368 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_369 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_370 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_339 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_340 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_341 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_342 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_343 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_344 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_345 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_346 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_347 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_348 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_349 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_350 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_351 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_352 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_353 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_354 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_371 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module rf_bypass ( .read1data({\read1data<15> , \read1data<14> , 
        \read1data<13> , \read1data<12> , \read1data<11> , \read1data<10> , 
        \read1data<9> , \read1data<8> , \read1data<7> , \read1data<6> , 
        \read1data<5> , \read1data<4> , \read1data<3> , \read1data<2> , 
        \read1data<1> , \read1data<0> }), .read2data({\read2data<15> , 
        \read2data<14> , \read2data<13> , \read2data<12> , \read2data<11> , 
        \read2data<10> , \read2data<9> , \read2data<8> , \read2data<7> , 
        \read2data<6> , \read2data<5> , \read2data<4> , \read2data<3> , 
        \read2data<2> , \read2data<1> , \read2data<0> }), err, clk, rst, 
    .read1regsel({\read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), 
    .read2regsel({\read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), 
    .writeregsel({\writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), 
    .writedata({\writedata<15> , \writedata<14> , \writedata<13> , 
        \writedata<12> , \writedata<11> , \writedata<10> , \writedata<9> , 
        \writedata<8> , \writedata<7> , \writedata<6> , \writedata<5> , 
        \writedata<4> , \writedata<3> , \writedata<2> , \writedata<1> , 
        \writedata<0> }), write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   \rf_r1_out<15> , \rf_r1_out<14> , \rf_r1_out<13> , \rf_r1_out<12> ,
         \rf_r1_out<11> , \rf_r1_out<10> , \rf_r1_out<9> , \rf_r1_out<8> ,
         \rf_r1_out<7> , \rf_r1_out<6> , \rf_r1_out<5> , \rf_r1_out<4> ,
         \rf_r1_out<3> , \rf_r1_out<2> , \rf_r1_out<1> , \rf_r1_out<0> ,
         \rf_r2_out<15> , \rf_r2_out<14> , \rf_r2_out<13> , \rf_r2_out<12> ,
         \rf_r2_out<11> , \rf_r2_out<10> , \rf_r2_out<9> , \rf_r2_out<8> ,
         \rf_r2_out<7> , \rf_r2_out<6> , \rf_r2_out<5> , \rf_r2_out<4> ,
         \rf_r2_out<3> , \rf_r2_out<2> , \rf_r2_out<1> , \rf_r2_out<0> , n19,
         n36, n37, n38, n39, n40, n57, n58, n59, n60, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;
  assign err = 1'b0;

  OAI21X1 U18 ( .A(n76), .B(n91), .C(n74), .Y(\read2data<9> ) );
  OAI21X1 U20 ( .A(n76), .B(n90), .C(n72), .Y(\read2data<8> ) );
  OAI21X1 U22 ( .A(n76), .B(n89), .C(n70), .Y(\read2data<7> ) );
  OAI21X1 U24 ( .A(n76), .B(n88), .C(n68), .Y(\read2data<6> ) );
  OAI21X1 U26 ( .A(n76), .B(n87), .C(n66), .Y(\read2data<5> ) );
  OAI21X1 U28 ( .A(n76), .B(n86), .C(n64), .Y(\read2data<4> ) );
  OAI21X1 U30 ( .A(n76), .B(n85), .C(n62), .Y(\read2data<3> ) );
  OAI21X1 U32 ( .A(n76), .B(n84), .C(n56), .Y(\read2data<2> ) );
  OAI21X1 U34 ( .A(n76), .B(n83), .C(n54), .Y(\read2data<1> ) );
  OAI21X1 U36 ( .A(n76), .B(n97), .C(n52), .Y(\read2data<15> ) );
  OAI21X1 U38 ( .A(n76), .B(n96), .C(n50), .Y(\read2data<14> ) );
  OAI21X1 U40 ( .A(n76), .B(n95), .C(n48), .Y(\read2data<13> ) );
  OAI21X1 U42 ( .A(n76), .B(n94), .C(n46), .Y(\read2data<12> ) );
  OAI21X1 U44 ( .A(n76), .B(n93), .C(n44), .Y(\read2data<11> ) );
  OAI21X1 U46 ( .A(n76), .B(n92), .C(n42), .Y(\read2data<10> ) );
  OAI21X1 U48 ( .A(n76), .B(n82), .C(n35), .Y(\read2data<0> ) );
  NAND3X1 U50 ( .A(n36), .B(n37), .C(n38), .Y(n19) );
  NOR2X1 U51 ( .A(n81), .B(n39), .Y(n38) );
  XOR2X1 U52 ( .A(n79), .B(\read2regsel<2> ), .Y(n39) );
  XNOR2X1 U53 ( .A(n77), .B(\read2regsel<1> ), .Y(n37) );
  XNOR2X1 U54 ( .A(\writeregsel<0> ), .B(\read2regsel<0> ), .Y(n36) );
  OAI21X1 U55 ( .A(n91), .B(n75), .C(n33), .Y(\read1data<9> ) );
  OAI21X1 U57 ( .A(n90), .B(n75), .C(n31), .Y(\read1data<8> ) );
  OAI21X1 U59 ( .A(n89), .B(n75), .C(n29), .Y(\read1data<7> ) );
  OAI21X1 U61 ( .A(n88), .B(n75), .C(n27), .Y(\read1data<6> ) );
  OAI21X1 U63 ( .A(n87), .B(n75), .C(n25), .Y(\read1data<5> ) );
  OAI21X1 U65 ( .A(n86), .B(n75), .C(n23), .Y(\read1data<4> ) );
  OAI21X1 U67 ( .A(n85), .B(n75), .C(n21), .Y(\read1data<3> ) );
  OAI21X1 U69 ( .A(n84), .B(n75), .C(n18), .Y(\read1data<2> ) );
  OAI21X1 U71 ( .A(n83), .B(n75), .C(n16), .Y(\read1data<1> ) );
  OAI21X1 U73 ( .A(n97), .B(n75), .C(n14), .Y(\read1data<15> ) );
  OAI21X1 U75 ( .A(n96), .B(n75), .C(n12), .Y(\read1data<14> ) );
  OAI21X1 U77 ( .A(n95), .B(n75), .C(n10), .Y(\read1data<13> ) );
  OAI21X1 U79 ( .A(n94), .B(n75), .C(n8), .Y(\read1data<12> ) );
  OAI21X1 U81 ( .A(n93), .B(n75), .C(n6), .Y(\read1data<11> ) );
  OAI21X1 U83 ( .A(n92), .B(n75), .C(n4), .Y(\read1data<10> ) );
  OAI21X1 U85 ( .A(n82), .B(n75), .C(n2), .Y(\read1data<0> ) );
  NAND3X1 U87 ( .A(n57), .B(n58), .C(n59), .Y(n40) );
  NOR2X1 U88 ( .A(n81), .B(n60), .Y(n59) );
  XOR2X1 U89 ( .A(n79), .B(\read1regsel<2> ), .Y(n60) );
  XNOR2X1 U90 ( .A(n77), .B(\read1regsel<1> ), .Y(n58) );
  XNOR2X1 U91 ( .A(\writeregsel<0> ), .B(\read1regsel<0> ), .Y(n57) );
  rf regfile ( .read1data({\rf_r1_out<15> , \rf_r1_out<14> , \rf_r1_out<13> , 
        \rf_r1_out<12> , \rf_r1_out<11> , \rf_r1_out<10> , \rf_r1_out<9> , 
        \rf_r1_out<8> , \rf_r1_out<7> , \rf_r1_out<6> , \rf_r1_out<5> , 
        \rf_r1_out<4> , \rf_r1_out<3> , \rf_r1_out<2> , \rf_r1_out<1> , 
        \rf_r1_out<0> }), .read2data({\rf_r2_out<15> , \rf_r2_out<14> , 
        \rf_r2_out<13> , \rf_r2_out<12> , \rf_r2_out<11> , \rf_r2_out<10> , 
        \rf_r2_out<9> , \rf_r2_out<8> , \rf_r2_out<7> , \rf_r2_out<6> , 
        \rf_r2_out<5> , \rf_r2_out<4> , \rf_r2_out<3> , \rf_r2_out<2> , 
        \rf_r2_out<1> , \rf_r2_out<0> }), .err(), .clk(clk), .rst(rst), 
        .read1regsel({\read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), 
        .read2regsel({\read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), 
        .writeregsel({n79, n77, \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        .write(write) );
  INVX1 U1 ( .A(\writedata<2> ), .Y(n84) );
  INVX1 U2 ( .A(\writedata<7> ), .Y(n89) );
  INVX1 U3 ( .A(\writedata<10> ), .Y(n92) );
  INVX1 U4 ( .A(\writedata<15> ), .Y(n97) );
  INVX1 U5 ( .A(write), .Y(n81) );
  INVX1 U6 ( .A(n80), .Y(n79) );
  INVX1 U7 ( .A(\writeregsel<2> ), .Y(n80) );
  INVX1 U8 ( .A(n78), .Y(n77) );
  INVX1 U9 ( .A(\writeregsel<1> ), .Y(n78) );
  INVX1 U10 ( .A(\writedata<0> ), .Y(n82) );
  INVX1 U11 ( .A(\writedata<1> ), .Y(n83) );
  INVX1 U12 ( .A(\writedata<3> ), .Y(n85) );
  INVX1 U13 ( .A(\writedata<4> ), .Y(n86) );
  INVX1 U14 ( .A(\writedata<5> ), .Y(n87) );
  INVX1 U15 ( .A(\writedata<6> ), .Y(n88) );
  INVX1 U16 ( .A(\writedata<8> ), .Y(n90) );
  INVX1 U17 ( .A(\writedata<9> ), .Y(n91) );
  INVX1 U19 ( .A(\writedata<11> ), .Y(n93) );
  INVX1 U21 ( .A(\writedata<12> ), .Y(n94) );
  INVX1 U23 ( .A(\writedata<13> ), .Y(n95) );
  INVX1 U25 ( .A(\writedata<14> ), .Y(n96) );
  AND2X1 U27 ( .A(\rf_r1_out<0> ), .B(n75), .Y(n1) );
  INVX1 U29 ( .A(n1), .Y(n2) );
  AND2X1 U31 ( .A(\rf_r1_out<10> ), .B(n75), .Y(n3) );
  INVX1 U33 ( .A(n3), .Y(n4) );
  AND2X1 U35 ( .A(\rf_r1_out<11> ), .B(n75), .Y(n5) );
  INVX1 U37 ( .A(n5), .Y(n6) );
  AND2X1 U39 ( .A(\rf_r1_out<12> ), .B(n75), .Y(n7) );
  INVX1 U41 ( .A(n7), .Y(n8) );
  AND2X1 U43 ( .A(\rf_r1_out<13> ), .B(n75), .Y(n9) );
  INVX1 U45 ( .A(n9), .Y(n10) );
  AND2X1 U47 ( .A(\rf_r1_out<14> ), .B(n75), .Y(n11) );
  INVX1 U49 ( .A(n11), .Y(n12) );
  AND2X1 U56 ( .A(\rf_r1_out<15> ), .B(n75), .Y(n13) );
  INVX1 U58 ( .A(n13), .Y(n14) );
  AND2X1 U60 ( .A(\rf_r1_out<1> ), .B(n75), .Y(n15) );
  INVX1 U62 ( .A(n15), .Y(n16) );
  AND2X1 U64 ( .A(\rf_r1_out<2> ), .B(n75), .Y(n17) );
  INVX1 U66 ( .A(n17), .Y(n18) );
  AND2X1 U68 ( .A(\rf_r1_out<3> ), .B(n75), .Y(n20) );
  INVX1 U70 ( .A(n20), .Y(n21) );
  AND2X1 U72 ( .A(\rf_r1_out<4> ), .B(n75), .Y(n22) );
  INVX1 U74 ( .A(n22), .Y(n23) );
  AND2X1 U76 ( .A(\rf_r1_out<5> ), .B(n75), .Y(n24) );
  INVX1 U78 ( .A(n24), .Y(n25) );
  AND2X1 U80 ( .A(\rf_r1_out<6> ), .B(n75), .Y(n26) );
  INVX1 U82 ( .A(n26), .Y(n27) );
  AND2X1 U84 ( .A(\rf_r1_out<7> ), .B(n75), .Y(n28) );
  INVX1 U86 ( .A(n28), .Y(n29) );
  AND2X1 U92 ( .A(\rf_r1_out<8> ), .B(n75), .Y(n30) );
  INVX1 U93 ( .A(n30), .Y(n31) );
  AND2X1 U94 ( .A(\rf_r1_out<9> ), .B(n75), .Y(n32) );
  INVX1 U95 ( .A(n32), .Y(n33) );
  AND2X1 U96 ( .A(\rf_r2_out<0> ), .B(n76), .Y(n34) );
  INVX1 U97 ( .A(n34), .Y(n35) );
  AND2X1 U98 ( .A(\rf_r2_out<10> ), .B(n76), .Y(n41) );
  INVX1 U99 ( .A(n41), .Y(n42) );
  AND2X1 U100 ( .A(\rf_r2_out<11> ), .B(n76), .Y(n43) );
  INVX1 U101 ( .A(n43), .Y(n44) );
  AND2X1 U102 ( .A(\rf_r2_out<12> ), .B(n76), .Y(n45) );
  INVX1 U103 ( .A(n45), .Y(n46) );
  AND2X1 U104 ( .A(\rf_r2_out<13> ), .B(n76), .Y(n47) );
  INVX1 U105 ( .A(n47), .Y(n48) );
  AND2X1 U106 ( .A(\rf_r2_out<14> ), .B(n76), .Y(n49) );
  INVX1 U107 ( .A(n49), .Y(n50) );
  AND2X1 U108 ( .A(\rf_r2_out<15> ), .B(n76), .Y(n51) );
  INVX1 U109 ( .A(n51), .Y(n52) );
  AND2X1 U110 ( .A(\rf_r2_out<1> ), .B(n76), .Y(n53) );
  INVX1 U111 ( .A(n53), .Y(n54) );
  AND2X1 U112 ( .A(\rf_r2_out<2> ), .B(n76), .Y(n55) );
  INVX1 U113 ( .A(n55), .Y(n56) );
  AND2X1 U114 ( .A(\rf_r2_out<3> ), .B(n76), .Y(n61) );
  INVX1 U115 ( .A(n61), .Y(n62) );
  AND2X1 U116 ( .A(\rf_r2_out<4> ), .B(n76), .Y(n63) );
  INVX1 U117 ( .A(n63), .Y(n64) );
  AND2X1 U118 ( .A(\rf_r2_out<5> ), .B(n76), .Y(n65) );
  INVX1 U119 ( .A(n65), .Y(n66) );
  AND2X1 U120 ( .A(\rf_r2_out<6> ), .B(n76), .Y(n67) );
  INVX1 U121 ( .A(n67), .Y(n68) );
  AND2X1 U122 ( .A(\rf_r2_out<7> ), .B(n76), .Y(n69) );
  INVX1 U123 ( .A(n69), .Y(n70) );
  AND2X1 U124 ( .A(\rf_r2_out<8> ), .B(n76), .Y(n71) );
  INVX1 U125 ( .A(n71), .Y(n72) );
  AND2X1 U126 ( .A(\rf_r2_out<9> ), .B(n76), .Y(n73) );
  INVX1 U127 ( .A(n73), .Y(n74) );
  BUFX2 U128 ( .A(n40), .Y(n75) );
  BUFX2 U129 ( .A(n19), .Y(n76) );
endmodule


module control_unit ( .opcode({\opcode<4> , \opcode<3> , \opcode<2> , 
        \opcode<1> , \opcode<0> }), .func({\func<1> , \func<0> }), .aluop({
        \aluop<2> , \aluop<1> , \aluop<0> }), alusrc, branch, jump, i1, i2, r, 
        jumpreg, set, btr, regwrite, memwrite, memread, memtoreg, invA, invB, 
        cin, excp, zeroext, halt, slbi, link, lbi, stu, rti );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ,
         \func<1> , \func<0> ;
  output \aluop<2> , \aluop<1> , \aluop<0> , alusrc, branch, jump, i1, i2, r,
         jumpreg, set, btr, regwrite, memwrite, memread, memtoreg, invA, invB,
         cin, excp, zeroext, halt, slbi, link, lbi, stu, rti;
  wire   n88, N34, N55, n24, n25, n26, n28, n32, n36, n37, n38, n39, n40, n41,
         n43, n44, n46, n47, n48, n49, n50, n51, n54, n1, n2, n3, n4, n6, n7,
         n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n27, n29, n30, n31, n33, n35, n45, n53, n55, n56, n57, n61, n62,
         n63, n65, n66, n67, n69, n70, n71, n73, n74, n75, n77, n78, n80, n81,
         n82, n83, n84, n85, n86, n87;

  AND2X2 U1 ( .A(n77), .B(n24), .Y(halt) );
  AND2X2 U2 ( .A(\opcode<1> ), .B(jump), .Y(link) );
  AND2X2 U3 ( .A(\opcode<0> ), .B(jump), .Y(jumpreg) );
  AND2X2 U4 ( .A(n24), .B(\opcode<2> ), .Y(jump) );
  AND2X2 U5 ( .A(n24), .B(n38), .Y(excp) );
  AND2X2 U6 ( .A(n47), .B(n48), .Y(n46) );
  OAI21X1 U26 ( .A(\opcode<4> ), .B(n8), .C(n70), .Y(zeroext) );
  NOR3X1 U27 ( .A(n78), .B(n81), .C(n18), .Y(stu) );
  NOR3X1 U28 ( .A(n29), .B(\opcode<2> ), .C(n81), .Y(rti) );
  NAND3X1 U32 ( .A(\opcode<1> ), .B(n86), .C(\opcode<2> ), .Y(n25) );
  OAI21X1 U36 ( .A(n80), .B(n14), .C(n1), .Y(invB) );
  NAND3X1 U37 ( .A(n66), .B(n36), .C(n70), .Y(n88) );
  AOI21X1 U38 ( .A(n84), .B(\opcode<0> ), .C(n4), .Y(n36) );
  OAI21X1 U40 ( .A(n38), .B(n6), .C(n40), .Y(i1) );
  NAND2X1 U41 ( .A(n82), .B(n87), .Y(n40) );
  NOR2X1 U42 ( .A(\opcode<3> ), .B(\opcode<4> ), .Y(n24) );
  OAI21X1 U43 ( .A(n80), .B(n14), .C(n74), .Y(cin) );
  OAI21X1 U44 ( .A(n41), .B(n23), .C(n43), .Y(invA) );
  NAND3X1 U45 ( .A(n82), .B(n87), .C(n15), .Y(n43) );
  NAND3X1 U47 ( .A(n7), .B(n75), .C(\opcode<4> ), .Y(n41) );
  NOR3X1 U48 ( .A(n16), .B(n12), .C(n87), .Y(btr) );
  OAI21X1 U52 ( .A(n77), .B(n87), .C(\opcode<3> ), .Y(n44) );
  NAND3X1 U53 ( .A(n81), .B(n83), .C(n78), .Y(n28) );
  NAND3X1 U54 ( .A(n1), .B(n70), .C(n46), .Y(N55) );
  NAND3X1 U55 ( .A(\opcode<0> ), .B(n85), .C(\opcode<2> ), .Y(n48) );
  NAND3X1 U56 ( .A(n38), .B(\opcode<4> ), .C(\func<0> ), .Y(n47) );
  NOR3X1 U58 ( .A(\opcode<0> ), .B(\opcode<2> ), .C(n81), .Y(n38) );
  OAI21X1 U60 ( .A(n73), .B(n75), .C(\opcode<4> ), .Y(n49) );
  NAND3X1 U61 ( .A(n50), .B(n51), .C(n62), .Y(N34) );
  NAND3X1 U66 ( .A(n85), .B(\opcode<1> ), .C(\opcode<2> ), .Y(n51) );
  OAI21X1 U67 ( .A(\func<1> ), .B(n87), .C(n7), .Y(n50) );
  NAND2X1 U69 ( .A(\opcode<3> ), .B(n83), .Y(n26) );
  NAND3X1 U72 ( .A(n32), .B(n83), .C(\opcode<4> ), .Y(n54) );
  OAI21X1 U73 ( .A(\opcode<0> ), .B(n81), .C(n16), .Y(n32) );
  NAND2X1 U76 ( .A(\opcode<4> ), .B(n86), .Y(n39) );
  NAND2X1 U77 ( .A(\opcode<2> ), .B(n87), .Y(n37) );
  OR2X1 U7 ( .A(n16), .B(n18), .Y(n63) );
  INVX1 U8 ( .A(invA), .Y(n74) );
  INVX1 U9 ( .A(n66), .Y(lbi) );
  INVX1 U10 ( .A(n70), .Y(slbi) );
  INVX1 U11 ( .A(\func<0> ), .Y(n73) );
  INVX1 U12 ( .A(\func<1> ), .Y(n75) );
  AND2X1 U13 ( .A(n31), .B(set), .Y(n61) );
  INVX1 U14 ( .A(n32), .Y(n80) );
  OR2X1 U15 ( .A(n32), .B(n18), .Y(n57) );
  INVX1 U16 ( .A(\opcode<0> ), .Y(n78) );
  OR2X1 U17 ( .A(n8), .B(n10), .Y(n1) );
  BUFX2 U18 ( .A(n28), .Y(n2) );
  OR2X2 U19 ( .A(n37), .B(n86), .Y(n3) );
  INVX1 U20 ( .A(n3), .Y(n4) );
  INVX1 U21 ( .A(n3), .Y(branch) );
  BUFX2 U22 ( .A(n39), .Y(n6) );
  AND2X2 U23 ( .A(\opcode<1> ), .B(n82), .Y(n7) );
  INVX1 U24 ( .A(n7), .Y(n8) );
  INVX1 U25 ( .A(n49), .Y(n9) );
  NOR2X1 U29 ( .A(n78), .B(n9), .Y(n11) );
  INVX1 U30 ( .A(n11), .Y(n10) );
  BUFX2 U31 ( .A(n26), .Y(n12) );
  AND2X2 U33 ( .A(\opcode<2> ), .B(n33), .Y(set) );
  INVX1 U34 ( .A(set), .Y(n14) );
  AND2X2 U35 ( .A(\opcode<0> ), .B(n81), .Y(n15) );
  INVX1 U39 ( .A(n15), .Y(n16) );
  AND2X2 U46 ( .A(n85), .B(n83), .Y(n17) );
  INVX1 U49 ( .A(n17), .Y(n18) );
  AND2X2 U50 ( .A(\opcode<3> ), .B(n54), .Y(n19) );
  AND2X2 U51 ( .A(\opcode<2> ), .B(n86), .Y(n20) );
  AND2X2 U57 ( .A(\opcode<4> ), .B(n2), .Y(n21) );
  AND2X2 U59 ( .A(\func<0> ), .B(\opcode<0> ), .Y(n22) );
  INVX1 U62 ( .A(n22), .Y(n23) );
  AND2X2 U63 ( .A(n24), .B(\opcode<0> ), .Y(n27) );
  INVX1 U64 ( .A(n27), .Y(n29) );
  OR2X2 U65 ( .A(\opcode<1> ), .B(\opcode<0> ), .Y(n30) );
  INVX1 U68 ( .A(n30), .Y(n31) );
  AND2X1 U70 ( .A(\opcode<4> ), .B(\opcode<3> ), .Y(n33) );
  INVX1 U71 ( .A(n28), .Y(n77) );
  INVX1 U74 ( .A(\opcode<4> ), .Y(n87) );
  INVX1 U75 ( .A(\opcode<3> ), .Y(n86) );
  INVX1 U78 ( .A(\opcode<2> ), .Y(n83) );
  OR2X1 U79 ( .A(n55), .B(n35), .Y(alusrc) );
  OR2X1 U80 ( .A(n20), .B(n85), .Y(n35) );
  OR2X1 U81 ( .A(n56), .B(n45), .Y(regwrite) );
  OR2X1 U82 ( .A(n21), .B(n82), .Y(n45) );
  OR2X1 U83 ( .A(n84), .B(n53), .Y(\aluop<2> ) );
  OR2X1 U84 ( .A(n19), .B(n17), .Y(n53) );
  INVX1 U85 ( .A(n44), .Y(n55) );
  INVX1 U86 ( .A(n25), .Y(n56) );
  INVX1 U87 ( .A(n57), .Y(memwrite) );
  BUFX2 U88 ( .A(N34), .Y(\aluop<1> ) );
  BUFX2 U89 ( .A(N55), .Y(\aluop<0> ) );
  INVX1 U90 ( .A(n37), .Y(n84) );
  INVX1 U91 ( .A(n61), .Y(n62) );
  INVX1 U92 ( .A(n63), .Y(memtoreg) );
  AND2X1 U93 ( .A(n77), .B(n33), .Y(n65) );
  INVX1 U94 ( .A(n65), .Y(n66) );
  INVX1 U95 ( .A(n26), .Y(n82) );
  INVX1 U96 ( .A(n88), .Y(n67) );
  INVX1 U97 ( .A(n67), .Y(i2) );
  AND2X1 U98 ( .A(n85), .B(n38), .Y(n69) );
  INVX1 U99 ( .A(n69), .Y(n70) );
  INVX1 U100 ( .A(n39), .Y(n85) );
  OAI21X1 U101 ( .A(\opcode<2> ), .B(n30), .C(n33), .Y(n71) );
  INVX2 U102 ( .A(n71), .Y(r) );
  BUFX2 U103 ( .A(memtoreg), .Y(memread) );
  INVX2 U104 ( .A(\opcode<1> ), .Y(n81) );
endmodule


module dff_338 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_304 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_305 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_306 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_307 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_308 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_309 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_310 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_311 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_312 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_313 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_314 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_315 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_316 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_317 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_318 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_319 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_337 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_336 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_335 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_301 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_302 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_303 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_285 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_286 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_287 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_288 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_289 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_290 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_291 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_292 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_293 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_294 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_295 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_296 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_297 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_298 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_299 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_300 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_334 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_282 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_283 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_284 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_279 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_280 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_281 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_276 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_277 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_278 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_264 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_265 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_266 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_267 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_268 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_269 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_270 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_271 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_272 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_273 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_274 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_275 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_333 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_332 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_331 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_330 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_329 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_328 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_327 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_326 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_325 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_324 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_323 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_322 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_321 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_320 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module alu ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , 
        \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> 
        }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , 
        \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> 
        }), Cin, .Op({\Op<2> , \Op<1> , \Op<0> }), invA, invB, sign, .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Ofl, Z, Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<2> , \Op<1> , \Op<0> , invA, invB, sign;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Ofl, Z, Cout;
  wire   \A_real<15> , \A_real<14> , \A_real<13> , \A_real<12> , \A_real<11> ,
         \A_real<10> , \A_real<9> , \A_real<8> , \A_real<7> , \A_real<6> ,
         \A_real<5> , \A_real<4> , \A_real<3> , \A_real<2> , \A_real<1> ,
         \A_real<0> , \B_real<15> , \B_real<13> , \B_real<11> , \B_real<10> ,
         \B_real<9> , \B_real<8> , \B_real<7> , \B_real<6> , \B_real<5> ,
         \B_real<4> , \B_real<3> , \B_real<2> , \B_real<1> , \B_real<0> ,
         \op0_out<15> , \op0_out<14> , \op0_out<13> , \op0_out<12> ,
         \op0_out<11> , \op0_out<10> , \op0_out<9> , \op0_out<8> ,
         \op0_out<7> , \op0_out<6> , \op0_out<5> , \op0_out<4> , \op0_out<3> ,
         \op0_out<2> , \op0_out<1> , \op0_out<0> , \op1_out<15> ,
         \op1_out<14> , \op1_out<13> , \op1_out<12> , \op1_out<11> ,
         \op1_out<10> , \op1_out<9> , \op1_out<8> , \op1_out<7> , \op1_out<6> ,
         \op1_out<5> , \op1_out<4> , \op1_out<3> , \op1_out<2> , \op1_out<1> ,
         \op1_out<0> , \op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> ,
         \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> ,
         \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> ,
         \op0_A<1> , \op0_A<0> , \op0_B<15> , \op0_B<14> , \op0_B<13> ,
         \op0_B<12> , \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> ,
         \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> ,
         \op0_B<2> , \op0_B<1> , \op0_B<0> , \op1_A<3> , \op1_A<2> ,
         \op1_A<1> , \op1_A<0> , \op1_B<15> , \op1_B<14> , \op1_B<13> ,
         \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> ,
         \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> ,
         \op1_B<2> , \op1_B<1> , \op1_B<0> , n59, n60, n62, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n61, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n144;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  OR2X2 U4 ( .A(\Op<1> ), .B(n104), .Y(n62) );
  OAI21X1 U74 ( .A(n111), .B(n144), .C(n54), .Y(\Out<0> ) );
  NAND3X1 U76 ( .A(Cout), .B(n111), .C(n90), .Y(n59) );
  demux1to2_16_1 demux0 ( .In({\A_real<15> , \A_real<14> , \A_real<13> , 
        \A_real<12> , \A_real<11> , \A_real<10> , \A_real<9> , \A_real<8> , 
        \A_real<7> , \A_real<6> , \A_real<5> , \A_real<4> , \A_real<3> , 
        \A_real<2> , \A_real<1> , \A_real<0> }), .S(n111), .Out0({\op0_A<15> , 
        \op0_A<14> , \op0_A<13> , \op0_A<12> , \op0_A<11> , \op0_A<10> , 
        \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , \op0_A<5> , \op0_A<4> , 
        \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .Out1({\op0_B<15> , 
        \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , \op0_B<10> , 
        \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , 
        \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }) );
  demux1to2_16_0 demux1 ( .In({\B_real<15> , n24, \B_real<13> , n22, 
        \B_real<11> , \B_real<10> , \B_real<9> , \B_real<8> , \B_real<7> , 
        \B_real<6> , \B_real<5> , \B_real<4> , \B_real<3> , \B_real<2> , 
        \B_real<1> , \B_real<0> }), .S(n111), .Out0({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, \op1_A<3> , \op1_A<2> , \op1_A<1> , 
        \op1_A<0> }), .Out1({\op1_B<15> , \op1_B<14> , \op1_B<13> , 
        \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , 
        \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> , 
        \op1_B<1> , \op1_B<0> }) );
  cla_or_xor_and coxa0 ( .A({\op0_B<15> , \op0_B<14> , \op0_B<13> , 
        \op0_B<12> , \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> , 
        \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , 
        \op0_B<1> , \op0_B<0> }), .B({\op1_B<15> , \op1_B<14> , \op1_B<13> , 
        \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , 
        \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> , 
        \op1_B<1> , \op1_B<0> }), .Cin(Cin), .Op({\Op<1> , \Op<0> }), .Out({
        \op0_out<15> , \op0_out<14> , \op0_out<13> , \op0_out<12> , 
        \op0_out<11> , \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , 
        \op0_out<6> , \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , 
        \op0_out<1> , \op0_out<0> }), .Cout(Cout) );
  shifter shift ( .In({\op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> , 
        \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> , 
        \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> , \op0_A<1> , 
        \op0_A<0> }), .Cnt({\op1_A<3> , \op1_A<2> , \op1_A<1> , \op1_A<0> }), 
        .Op({\Op<1> , n104}), .Out({\op1_out<15> , \op1_out<14> , 
        \op1_out<13> , \op1_out<12> , \op1_out<11> , \op1_out<10> , 
        \op1_out<9> , \op1_out<8> , \op1_out<7> , \op1_out<6> , \op1_out<5> , 
        \op1_out<4> , \op1_out<3> , \op1_out<2> , \op1_out<1> , \op1_out<0> })
         );
  BUFX2 U1 ( .A(\op0_out<8> ), .Y(n1) );
  XNOR2X1 U2 ( .A(\B<2> ), .B(n105), .Y(\B_real<2> ) );
  INVX1 U3 ( .A(n105), .Y(n16) );
  INVX1 U5 ( .A(n109), .Y(n12) );
  INVX1 U6 ( .A(n109), .Y(n19) );
  INVX1 U7 ( .A(n139), .Y(\A_real<15> ) );
  INVX1 U8 ( .A(n107), .Y(n18) );
  OR2X1 U9 ( .A(\op1_out<10> ), .B(\op1_out<11> ), .Y(n49) );
  INVX1 U10 ( .A(n12), .Y(n10) );
  AND2X1 U11 ( .A(n40), .B(n35), .Y(n88) );
  INVX1 U12 ( .A(\op0_out<2> ), .Y(n115) );
  INVX1 U13 ( .A(\op1_out<6> ), .Y(n124) );
  INVX1 U14 ( .A(\op0_out<6> ), .Y(n123) );
  INVX1 U15 ( .A(\op1_out<7> ), .Y(n125) );
  INVX1 U16 ( .A(\op1_out<8> ), .Y(n127) );
  INVX1 U17 ( .A(\op1_out<9> ), .Y(n129) );
  INVX1 U18 ( .A(\op1_out<10> ), .Y(n131) );
  INVX1 U19 ( .A(\op1_out<11> ), .Y(n133) );
  INVX1 U20 ( .A(\op1_out<12> ), .Y(n135) );
  INVX1 U21 ( .A(\op1_out<13> ), .Y(n136) );
  INVX1 U22 ( .A(\op1_out<14> ), .Y(n138) );
  INVX1 U23 ( .A(\op0_out<10> ), .Y(n2) );
  INVX1 U24 ( .A(n2), .Y(n3) );
  MUX2X1 U25 ( .B(n132), .A(n133), .S(n112), .Y(\Out<11> ) );
  INVX1 U26 ( .A(n81), .Y(n4) );
  INVX1 U27 ( .A(n4), .Y(n5) );
  INVX1 U28 ( .A(\op0_out<7> ), .Y(n6) );
  OR2X2 U29 ( .A(n61), .B(n85), .Y(n7) );
  OR2X2 U30 ( .A(\op0_out<13> ), .B(n82), .Y(n8) );
  NOR2X1 U31 ( .A(n8), .B(n9), .Y(n79) );
  OR2X2 U32 ( .A(n14), .B(n3), .Y(n9) );
  XOR2X1 U33 ( .A(\A<2> ), .B(n10), .Y(\A_real<2> ) );
  XOR2X1 U34 ( .A(\B<4> ), .B(n106), .Y(\B_real<4> ) );
  INVX1 U35 ( .A(\op0_out<13> ), .Y(n11) );
  MUX2X1 U36 ( .B(n11), .A(n136), .S(n112), .Y(\Out<13> ) );
  BUFX2 U37 ( .A(\op0_out<4> ), .Y(n13) );
  XOR2X1 U38 ( .A(\B<7> ), .B(n107), .Y(\B_real<7> ) );
  OR2X2 U39 ( .A(\op0_out<11> ), .B(n112), .Y(n14) );
  XNOR2X1 U40 ( .A(n15), .B(n110), .Y(\A_real<1> ) );
  INVX1 U41 ( .A(\A<1> ), .Y(n15) );
  INVX2 U42 ( .A(n108), .Y(n110) );
  XOR2X1 U43 ( .A(\B<1> ), .B(n16), .Y(\B_real<1> ) );
  XOR2X1 U44 ( .A(\B<6> ), .B(n17), .Y(\B_real<6> ) );
  INVX1 U45 ( .A(n105), .Y(n17) );
  XNOR2X1 U46 ( .A(\A<8> ), .B(n94), .Y(\A_real<8> ) );
  INVX1 U47 ( .A(n109), .Y(n94) );
  XNOR2X1 U48 ( .A(\A<9> ), .B(n99), .Y(\A_real<9> ) );
  XOR2X1 U49 ( .A(\B<5> ), .B(n17), .Y(\B_real<5> ) );
  XNOR2X1 U50 ( .A(\B<9> ), .B(n18), .Y(\B_real<9> ) );
  OR2X2 U51 ( .A(\op0_out<1> ), .B(\op0_out<0> ), .Y(n85) );
  XNOR2X1 U52 ( .A(\A<10> ), .B(n19), .Y(\A_real<10> ) );
  XNOR2X1 U53 ( .A(\B<0> ), .B(n105), .Y(\B_real<0> ) );
  XOR2X1 U54 ( .A(\B<10> ), .B(n106), .Y(\B_real<10> ) );
  XNOR2X1 U55 ( .A(n20), .B(n106), .Y(\B_real<8> ) );
  INVX1 U56 ( .A(\B<8> ), .Y(n20) );
  INVX8 U57 ( .A(n105), .Y(n107) );
  INVX1 U58 ( .A(n13), .Y(n119) );
  AND2X2 U59 ( .A(n66), .B(n56), .Y(n21) );
  INVX1 U60 ( .A(n21), .Y(n22) );
  AND2X2 U61 ( .A(n102), .B(n103), .Y(n23) );
  INVX1 U62 ( .A(n23), .Y(n24) );
  AND2X2 U63 ( .A(n70), .B(n64), .Y(n25) );
  INVX1 U64 ( .A(n25), .Y(\Out<1> ) );
  OR2X2 U65 ( .A(n87), .B(n28), .Y(n27) );
  OR2X2 U66 ( .A(n36), .B(n86), .Y(n28) );
  OR2X2 U67 ( .A(n7), .B(\op0_out<3> ), .Y(n29) );
  OR2X2 U68 ( .A(n29), .B(\op0_out<8> ), .Y(n30) );
  OR2X2 U69 ( .A(n33), .B(n37), .Y(n31) );
  OR2X2 U70 ( .A(\op0_out<9> ), .B(\op0_out<6> ), .Y(n32) );
  OR2X2 U71 ( .A(n72), .B(n32), .Y(n33) );
  OR2X1 U72 ( .A(\op1_out<6> ), .B(\op1_out<7> ), .Y(n34) );
  INVX1 U73 ( .A(n34), .Y(n35) );
  OR2X2 U75 ( .A(\op1_out<3> ), .B(\op1_out<2> ), .Y(n36) );
  OR2X2 U77 ( .A(n91), .B(n5), .Y(n37) );
  AND2X2 U78 ( .A(\op1_out<15> ), .B(n112), .Y(n38) );
  OR2X1 U79 ( .A(\op1_out<4> ), .B(\op1_out<5> ), .Y(n39) );
  INVX1 U80 ( .A(n39), .Y(n40) );
  OR2X2 U81 ( .A(\op1_out<12> ), .B(\op1_out<13> ), .Y(n41) );
  INVX1 U82 ( .A(n41), .Y(n42) );
  OR2X2 U83 ( .A(\op1_out<8> ), .B(\op1_out<9> ), .Y(n43) );
  INVX1 U84 ( .A(n43), .Y(n44) );
  OR2X2 U85 ( .A(\op0_out<12> ), .B(n30), .Y(n45) );
  INVX1 U86 ( .A(n45), .Y(n46) );
  OR2X2 U87 ( .A(\op1_out<14> ), .B(\op1_out<15> ), .Y(n47) );
  INVX1 U88 ( .A(n47), .Y(n48) );
  INVX1 U89 ( .A(n49), .Y(n50) );
  AND2X2 U90 ( .A(n68), .B(n58), .Y(n51) );
  INVX1 U91 ( .A(n51), .Y(n52) );
  AND2X2 U92 ( .A(\op0_out<0> ), .B(n111), .Y(n53) );
  INVX1 U93 ( .A(n53), .Y(n54) );
  AND2X2 U94 ( .A(n97), .B(n106), .Y(n55) );
  INVX1 U95 ( .A(n55), .Y(n56) );
  OR2X2 U96 ( .A(n74), .B(n76), .Y(n57) );
  INVX1 U97 ( .A(n57), .Y(n58) );
  OR2X2 U98 ( .A(\op0_out<4> ), .B(\op0_out<2> ), .Y(n61) );
  AND2X2 U99 ( .A(\op1_out<1> ), .B(n112), .Y(n63) );
  INVX1 U100 ( .A(n63), .Y(n64) );
  AND2X2 U101 ( .A(n84), .B(n101), .Y(n65) );
  INVX1 U102 ( .A(n65), .Y(n66) );
  OR2X2 U103 ( .A(n27), .B(n89), .Y(n67) );
  INVX1 U104 ( .A(n67), .Y(n68) );
  AND2X2 U105 ( .A(\op0_out<1> ), .B(n111), .Y(n69) );
  INVX1 U106 ( .A(n69), .Y(n70) );
  AND2X2 U107 ( .A(n46), .B(n121), .Y(n71) );
  INVX1 U108 ( .A(n71), .Y(n72) );
  AND2X2 U109 ( .A(n42), .B(n48), .Y(n73) );
  INVX1 U110 ( .A(n73), .Y(n74) );
  AND2X2 U111 ( .A(n44), .B(n50), .Y(n75) );
  INVX1 U112 ( .A(n75), .Y(n76) );
  OR2X2 U113 ( .A(n81), .B(n38), .Y(n77) );
  INVX1 U114 ( .A(n77), .Y(n78) );
  INVX1 U115 ( .A(n79), .Y(n80) );
  BUFX2 U116 ( .A(\op0_out<15> ), .Y(n81) );
  BUFX2 U117 ( .A(\op0_out<7> ), .Y(n82) );
  INVX1 U118 ( .A(n38), .Y(n83) );
  INVX1 U119 ( .A(n97), .Y(n84) );
  INVX1 U120 ( .A(n113), .Y(n86) );
  INVX1 U121 ( .A(n114), .Y(n87) );
  INVX1 U122 ( .A(n88), .Y(n89) );
  INVX1 U123 ( .A(\op0_out<5> ), .Y(n121) );
  INVX1 U124 ( .A(n59), .Y(Ofl) );
  BUFX2 U125 ( .A(n60), .Y(n90) );
  OAI21X1 U126 ( .A(n80), .B(n31), .C(n52), .Y(Z) );
  XOR2X1 U127 ( .A(\B<3> ), .B(n92), .Y(\B_real<3> ) );
  INVX1 U128 ( .A(n105), .Y(n92) );
  BUFX2 U129 ( .A(\op0_out<14> ), .Y(n91) );
  INVX1 U130 ( .A(\op0_out<3> ), .Y(n117) );
  INVX1 U131 ( .A(n110), .Y(n99) );
  INVX1 U132 ( .A(n110), .Y(n98) );
  INVX1 U133 ( .A(n110), .Y(n93) );
  XNOR2X1 U134 ( .A(\A<3> ), .B(n108), .Y(\A_real<3> ) );
  INVX4 U135 ( .A(n105), .Y(n106) );
  XNOR2X1 U136 ( .A(\A<11> ), .B(n93), .Y(\A_real<11> ) );
  INVX1 U137 ( .A(\op1_out<3> ), .Y(n118) );
  XNOR2X1 U138 ( .A(\A<6> ), .B(n94), .Y(\A_real<6> ) );
  INVX1 U139 ( .A(n109), .Y(n96) );
  INVX1 U140 ( .A(n109), .Y(n95) );
  INVX1 U141 ( .A(\op1_out<0> ), .Y(n144) );
  INVX1 U142 ( .A(\op1_out<4> ), .Y(n120) );
  XNOR2X1 U143 ( .A(\A<14> ), .B(n95), .Y(\A_real<14> ) );
  INVX1 U144 ( .A(\op1_out<1> ), .Y(n114) );
  INVX1 U145 ( .A(\op1_out<2> ), .Y(n116) );
  INVX1 U146 ( .A(\op0_out<9> ), .Y(n128) );
  XOR2X1 U147 ( .A(\A<0> ), .B(n109), .Y(\A_real<0> ) );
  XNOR2X1 U148 ( .A(\A<4> ), .B(n96), .Y(\A_real<4> ) );
  INVX1 U149 ( .A(\B<12> ), .Y(n97) );
  INVX1 U150 ( .A(\op0_out<11> ), .Y(n132) );
  INVX1 U151 ( .A(\op1_out<5> ), .Y(n122) );
  INVX1 U152 ( .A(\op0_out<10> ), .Y(n130) );
  XNOR2X1 U153 ( .A(\A<7> ), .B(n98), .Y(\A_real<7> ) );
  NAND2X1 U154 ( .A(n101), .B(\B<14> ), .Y(n102) );
  NAND2X1 U155 ( .A(n100), .B(n106), .Y(n103) );
  INVX1 U156 ( .A(\B<14> ), .Y(n100) );
  INVX1 U157 ( .A(n106), .Y(n101) );
  INVX1 U158 ( .A(\op0_out<12> ), .Y(n134) );
  BUFX2 U159 ( .A(\Op<0> ), .Y(n104) );
  INVX1 U160 ( .A(n91), .Y(n137) );
  INVX1 U161 ( .A(n1), .Y(n126) );
  INVX8 U162 ( .A(invB), .Y(n105) );
  INVX8 U163 ( .A(invA), .Y(n108) );
  INVX8 U164 ( .A(n108), .Y(n109) );
  INVX8 U165 ( .A(n112), .Y(n111) );
  INVX8 U166 ( .A(\Op<2> ), .Y(n112) );
  XNOR2X1 U167 ( .A(\B<15> ), .B(n107), .Y(n140) );
  INVX2 U168 ( .A(n140), .Y(\B_real<15> ) );
  XOR2X1 U169 ( .A(\B<13> ), .B(n107), .Y(\B_real<13> ) );
  XOR2X1 U170 ( .A(\B<11> ), .B(n107), .Y(\B_real<11> ) );
  XNOR2X1 U171 ( .A(\A<15> ), .B(n110), .Y(n139) );
  XOR2X1 U172 ( .A(\A<13> ), .B(n110), .Y(\A_real<13> ) );
  XOR2X1 U173 ( .A(\A<12> ), .B(n109), .Y(\A_real<12> ) );
  XOR2X1 U174 ( .A(\A<5> ), .B(n110), .Y(\A_real<5> ) );
  NOR2X1 U175 ( .A(n111), .B(\op1_out<0> ), .Y(n113) );
  MUX2X1 U176 ( .B(n116), .A(n115), .S(n111), .Y(\Out<2> ) );
  MUX2X1 U177 ( .B(n118), .A(n117), .S(n111), .Y(\Out<3> ) );
  MUX2X1 U178 ( .B(n120), .A(n119), .S(n111), .Y(\Out<4> ) );
  MUX2X1 U179 ( .B(n122), .A(n121), .S(n111), .Y(\Out<5> ) );
  MUX2X1 U180 ( .B(n124), .A(n123), .S(n111), .Y(\Out<6> ) );
  MUX2X1 U181 ( .B(n125), .A(n6), .S(n111), .Y(\Out<7> ) );
  MUX2X1 U182 ( .B(n127), .A(n126), .S(n111), .Y(\Out<8> ) );
  MUX2X1 U183 ( .B(n129), .A(n128), .S(n111), .Y(\Out<9> ) );
  MUX2X1 U184 ( .B(n131), .A(n130), .S(n111), .Y(\Out<10> ) );
  MUX2X1 U185 ( .B(n135), .A(n134), .S(n111), .Y(\Out<12> ) );
  MUX2X1 U186 ( .B(n138), .A(n137), .S(n111), .Y(\Out<14> ) );
  AOI21X1 U187 ( .A(n112), .B(n83), .C(n78), .Y(\Out<15> ) );
  XNOR2X1 U188 ( .A(n140), .B(n139), .Y(n141) );
  AOI21X1 U189 ( .A(sign), .B(n141), .C(n62), .Y(n60) );
endmodule


module mux4to1_16_5 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n3, n4, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n1, n2, n5, n6, n7, n8, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72,
         n74, n76, n78, n80, n82, n84, n86, n88, n90, n92, n94, n96, n98, n100,
         n101, n102, n103, n104;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n104), .C(\InB<9> ), .D(n8), .Y(n4) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n38), .C(\InD<9> ), .D(n37), .Y(n3) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n104), .C(\InB<8> ), .D(n8), .Y(n10) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n38), .C(\InD<8> ), .D(n37), .Y(n9) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n104), .C(\InB<7> ), .D(n8), .Y(n12) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n38), .C(\InD<7> ), .D(n37), .Y(n11) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n104), .C(\InB<6> ), .D(n8), .Y(n14) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n38), .C(\InD<6> ), .D(n37), .Y(n13) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n104), .C(\InB<5> ), .D(n8), .Y(n16) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n38), .C(\InD<5> ), .D(n37), .Y(n15) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n104), .C(\InB<4> ), .D(n8), .Y(n18) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n38), .C(\InD<4> ), .D(n37), .Y(n17) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n104), .C(\InB<3> ), .D(n8), .Y(n20) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n38), .C(\InD<3> ), .D(n37), .Y(n19) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n104), .C(\InB<2> ), .D(n8), .Y(n22) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n38), .C(\InD<2> ), .D(n37), .Y(n21) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n104), .C(\InB<1> ), .D(n8), .Y(n24) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n38), .C(\InD<1> ), .D(n37), .Y(n23) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n104), .C(\InB<15> ), .D(n8), .Y(n26) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n38), .C(\InD<15> ), .D(n37), .Y(n25) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n104), .C(\InB<14> ), .D(n8), .Y(n28) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n38), .C(\InD<14> ), .D(n37), .Y(n27) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n104), .C(\InB<13> ), .D(n8), .Y(n30) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n38), .C(\InD<13> ), .D(n37), .Y(n29) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n104), .C(\InB<12> ), .D(n8), .Y(n32) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n38), .C(\InD<12> ), .D(n37), .Y(n31) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n104), .C(\InB<11> ), .D(n8), .Y(n34) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n38), .C(\InD<11> ), .D(n37), .Y(n33) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n104), .C(\InB<10> ), .D(n8), .Y(n36) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n38), .C(\InD<10> ), .D(n37), .Y(n35) );
  INVX1 U1 ( .A(\S<0> ), .Y(n102) );
  OR2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n101) );
  INVX1 U3 ( .A(\S<1> ), .Y(n100) );
  AND2X1 U4 ( .A(n45), .B(n60), .Y(n70) );
  AND2X1 U7 ( .A(n46), .B(n61), .Y(n84) );
  AND2X1 U10 ( .A(n47), .B(n62), .Y(n86) );
  AND2X1 U13 ( .A(n48), .B(n63), .Y(n88) );
  AND2X1 U16 ( .A(n49), .B(n64), .Y(n90) );
  AND2X1 U19 ( .A(n50), .B(n65), .Y(n92) );
  AND2X1 U22 ( .A(n51), .B(n66), .Y(n94) );
  AND2X1 U25 ( .A(n52), .B(n67), .Y(n96) );
  AND2X1 U28 ( .A(n53), .B(n68), .Y(n98) );
  AND2X1 U31 ( .A(n39), .B(n54), .Y(n72) );
  AND2X1 U34 ( .A(n40), .B(n55), .Y(n74) );
  AND2X1 U37 ( .A(n41), .B(n56), .Y(n76) );
  AND2X1 U40 ( .A(n42), .B(n57), .Y(n78) );
  AND2X1 U43 ( .A(n43), .B(n58), .Y(n80) );
  AND2X1 U46 ( .A(n44), .B(n59), .Y(n82) );
  OR2X1 U49 ( .A(n8), .B(n69), .Y(n1) );
  INVX1 U50 ( .A(n1), .Y(n2) );
  BUFX2 U51 ( .A(n103), .Y(n5) );
  OR2X2 U52 ( .A(n69), .B(\InB<0> ), .Y(n6) );
  INVX1 U53 ( .A(n6), .Y(n7) );
  AND2X1 U54 ( .A(\S<0> ), .B(n100), .Y(n8) );
  AND2X1 U55 ( .A(\S<0> ), .B(\S<1> ), .Y(n37) );
  AND2X1 U56 ( .A(n102), .B(\S<1> ), .Y(n38) );
  BUFX2 U57 ( .A(n35), .Y(n39) );
  BUFX2 U58 ( .A(n33), .Y(n40) );
  BUFX2 U59 ( .A(n31), .Y(n41) );
  BUFX2 U60 ( .A(n29), .Y(n42) );
  BUFX2 U61 ( .A(n27), .Y(n43) );
  BUFX2 U62 ( .A(n25), .Y(n44) );
  BUFX2 U63 ( .A(n23), .Y(n45) );
  BUFX2 U64 ( .A(n21), .Y(n46) );
  BUFX2 U65 ( .A(n19), .Y(n47) );
  BUFX2 U66 ( .A(n17), .Y(n48) );
  BUFX2 U67 ( .A(n15), .Y(n49) );
  BUFX2 U68 ( .A(n13), .Y(n50) );
  BUFX2 U69 ( .A(n11), .Y(n51) );
  BUFX2 U70 ( .A(n9), .Y(n52) );
  BUFX2 U71 ( .A(n3), .Y(n53) );
  BUFX2 U72 ( .A(n36), .Y(n54) );
  BUFX2 U73 ( .A(n34), .Y(n55) );
  BUFX2 U74 ( .A(n32), .Y(n56) );
  BUFX2 U75 ( .A(n30), .Y(n57) );
  BUFX2 U76 ( .A(n28), .Y(n58) );
  BUFX2 U77 ( .A(n26), .Y(n59) );
  BUFX2 U78 ( .A(n24), .Y(n60) );
  BUFX2 U79 ( .A(n22), .Y(n61) );
  BUFX2 U80 ( .A(n20), .Y(n62) );
  BUFX2 U81 ( .A(n18), .Y(n63) );
  BUFX2 U82 ( .A(n16), .Y(n64) );
  BUFX2 U83 ( .A(n14), .Y(n65) );
  BUFX2 U84 ( .A(n12), .Y(n66) );
  BUFX2 U85 ( .A(n10), .Y(n67) );
  BUFX2 U86 ( .A(n4), .Y(n68) );
  AND2X1 U87 ( .A(\InD<0> ), .B(n37), .Y(n69) );
  INVX1 U88 ( .A(n70), .Y(\Out<1> ) );
  INVX1 U89 ( .A(n72), .Y(\Out<10> ) );
  INVX1 U90 ( .A(n74), .Y(\Out<11> ) );
  INVX1 U91 ( .A(n76), .Y(\Out<12> ) );
  INVX1 U92 ( .A(n78), .Y(\Out<13> ) );
  INVX1 U93 ( .A(n80), .Y(\Out<14> ) );
  INVX1 U94 ( .A(n82), .Y(\Out<15> ) );
  INVX1 U95 ( .A(n84), .Y(\Out<2> ) );
  INVX1 U96 ( .A(n86), .Y(\Out<3> ) );
  INVX1 U97 ( .A(n88), .Y(\Out<4> ) );
  INVX1 U98 ( .A(n90), .Y(\Out<5> ) );
  INVX1 U99 ( .A(n92), .Y(\Out<6> ) );
  INVX1 U100 ( .A(n94), .Y(\Out<7> ) );
  INVX1 U101 ( .A(n96), .Y(\Out<8> ) );
  INVX1 U102 ( .A(n98), .Y(\Out<9> ) );
  AOI22X1 U103 ( .A(n104), .B(\InA<0> ), .C(n38), .D(\InC<0> ), .Y(n103) );
  INVX1 U104 ( .A(n101), .Y(n104) );
  OAI21X1 U105 ( .A(n2), .B(n7), .C(n5), .Y(\Out<0> ) );
endmodule


module cla16_1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n1,
         n2, n3, n9, n10, n11, n12, n13, n14, n15;

  AOI21X1 U5 ( .A(\P<3> ), .B(n9), .C(\G<3> ), .Y(n15) );
  AOI21X1 U6 ( .A(\P<2> ), .B(n10), .C(\G<2> ), .Y(n14) );
  AOI21X1 U7 ( .A(\P<1> ), .B(n11), .C(\G<1> ), .Y(n13) );
  AOI21X1 U8 ( .A(\P<0> ), .B(Cin), .C(\G<0> ), .Y(n12) );
  cla4_7 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_6 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n2), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_5 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n10), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_4 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n9), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  BUFX2 U1 ( .A(n13), .Y(n1) );
  BUFX2 U2 ( .A(n11), .Y(n2) );
  INVX1 U3 ( .A(n12), .Y(n11) );
  INVX1 U4 ( .A(n14), .Y(n9) );
  BUFX2 U9 ( .A(n15), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(Cout) );
  INVX2 U11 ( .A(n1), .Y(n10) );
endmodule


module mux4to1 ( InA, InB, InC, InD, .S({\S<1> , \S<0> }), Out );
  input InA, InB, InC, InD, \S<1> , \S<0> ;
  output Out;
  wire   n4, n5, n6, n1, n2;

  OAI21X1 U3 ( .A(\S<1> ), .B(n4), .C(n5), .Y(Out) );
  NAND2X1 U4 ( .A(n1), .B(\S<1> ), .Y(n5) );
  AOI22X1 U5 ( .A(InC), .B(n2), .C(InD), .D(\S<0> ), .Y(n6) );
  AOI22X1 U6 ( .A(InA), .B(n2), .C(\S<0> ), .D(InB), .Y(n4) );
  INVX1 U1 ( .A(\S<0> ), .Y(n2) );
  INVX1 U2 ( .A(n6), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module stallmem ( .DataOut({\DataOut<15> , \DataOut<14> , \DataOut<13> , 
        \DataOut<12> , \DataOut<11> , \DataOut<10> , \DataOut<9> , 
        \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , 
        \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), Done, Stall, 
        CacheHit, err, .Addr({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> , \Addr<10> , \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , 
        \Addr<5> , \Addr<4> , \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> }), 
    .DataIn({\DataIn<15> , \DataIn<14> , \DataIn<13> , \DataIn<12> , 
        \DataIn<11> , \DataIn<10> , \DataIn<9> , \DataIn<8> , \DataIn<7> , 
        \DataIn<6> , \DataIn<5> , \DataIn<4> , \DataIn<3> , \DataIn<2> , 
        \DataIn<1> , \DataIn<0> }), Rd, Wr, createdump, clk, rst );
  input \Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , \Addr<11> , \Addr<10> ,
         \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , \Addr<5> , \Addr<4> ,
         \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> , \DataIn<15> ,
         \DataIn<14> , \DataIn<13> , \DataIn<12> , \DataIn<11> , \DataIn<10> ,
         \DataIn<9> , \DataIn<8> , \DataIn<7> , \DataIn<6> , \DataIn<5> ,
         \DataIn<4> , \DataIn<3> , \DataIn<2> , \DataIn<1> , \DataIn<0> , Rd,
         Wr, createdump, clk, rst;
  output \DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> ,
         \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> ,
         \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> ,
         \DataOut<2> , \DataOut<1> , \DataOut<0> , Done, Stall, CacheHit, err;
  wire   N253, N254, N255, N256, N257, N258, n2581, \rand_pat<31> ,
         \rand_pat<30> , \rand_pat<29> , \rand_pat<28> , \rand_pat<27> ,
         \rand_pat<26> , \rand_pat<25> , \rand_pat<24> , \rand_pat<23> ,
         \rand_pat<22> , \rand_pat<21> , \rand_pat<20> , \rand_pat<19> ,
         \rand_pat<18> , \rand_pat<17> , \rand_pat<16> , \rand_pat<15> ,
         \rand_pat<14> , \rand_pat<13> , \rand_pat<12> , \rand_pat<11> ,
         \rand_pat<10> , \rand_pat<9> , \rand_pat<8> , \rand_pat<7> ,
         \rand_pat<6> , \rand_pat<5> , \rand_pat<4> , \rand_pat<3> ,
         \rand_pat<2> , \rand_pat<1> , \rand_pat<0> , \mem<0><7> , \mem<0><6> ,
         \mem<0><5> , \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> ,
         \mem<0><0> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> ,
         \mem<2><6> , \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> ,
         \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> ,
         \mem<4><7> , \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> ,
         \mem<4><2> , \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> ,
         \mem<5><5> , \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> ,
         \mem<5><0> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> ,
         \mem<7><6> , \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> ,
         \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> ,
         \mem<9><7> , \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> ,
         \mem<9><2> , \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> ,
         \mem<10><5> , \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> ,
         \mem<10><0> , \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> ,
         \mem<11><3> , \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> ,
         \mem<12><6> , \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> ,
         \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> ,
         \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> ,
         \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> ,
         \mem<17><6> , \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> ,
         \mem<18><4> , \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> ,
         \mem<19><7> , \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> ,
         \mem<19><2> , \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> ,
         \mem<20><5> , \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> ,
         \mem<20><0> , \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> ,
         \mem<21><3> , \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> ,
         \mem<22><6> , \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> ,
         \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> ,
         \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> ,
         \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> ,
         \mem<27><6> , \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> ,
         \mem<28><4> , \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> ,
         \mem<29><7> , \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> ,
         \mem<29><2> , \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> ,
         \mem<30><5> , \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> ,
         \mem<30><0> , \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> ,
         \mem<31><3> , \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> ,
         \mem<32><6> , \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> ,
         \mem<32><1> , \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> ,
         \mem<33><4> , \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> ,
         \mem<34><7> , \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> ,
         \mem<34><2> , \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> ,
         \mem<35><5> , \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> ,
         \mem<35><0> , \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> ,
         \mem<36><3> , \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> ,
         \mem<37><6> , \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> ,
         \mem<37><1> , \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> ,
         \mem<38><4> , \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> ,
         \mem<39><7> , \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> ,
         \mem<39><2> , \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> ,
         \mem<40><5> , \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> ,
         \mem<40><0> , \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> ,
         \mem<41><3> , \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> ,
         \mem<42><6> , \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> ,
         \mem<42><1> , \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> ,
         \mem<43><4> , \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> ,
         \mem<44><7> , \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> ,
         \mem<44><2> , \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> ,
         \mem<45><5> , \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> ,
         \mem<45><0> , \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> ,
         \mem<46><3> , \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> ,
         \mem<47><6> , \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> ,
         \mem<47><1> , \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> ,
         \mem<48><4> , \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> ,
         \mem<49><7> , \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> ,
         \mem<49><2> , \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> ,
         \mem<50><5> , \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> ,
         \mem<50><0> , \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> ,
         \mem<51><3> , \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> ,
         \mem<52><6> , \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> ,
         \mem<52><1> , \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> ,
         \mem<53><4> , \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> ,
         \mem<54><7> , \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> ,
         \mem<54><2> , \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> ,
         \mem<55><5> , \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> ,
         \mem<55><0> , \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> ,
         \mem<56><3> , \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> ,
         \mem<57><6> , \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> ,
         \mem<57><1> , \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> ,
         \mem<58><4> , \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> ,
         \mem<59><7> , \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> ,
         \mem<59><2> , \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> ,
         \mem<60><5> , \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> ,
         \mem<60><0> , \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> ,
         \mem<61><3> , \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> ,
         \mem<62><6> , \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> ,
         \mem<62><1> , \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> ,
         \mem<63><4> , \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> ,
         N259, N260, N261, N262, N263, N264, N265, N266, n4, n6, n8, n10, n12,
         n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34, n35, n36, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n598, n600, n602, n604,
         n606, n608, n610, n612, n614, n616, n618, n620, n622, n624, n626,
         n628, n630, n632, n634, n636, n638, n640, n642, n644, n646, n648,
         n650, n652, n654, n656, n658, n660, n662, n663, n666, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n725, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n754, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n781, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n808, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n835, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n862, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n889, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n916, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n943, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n970, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n997, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1024,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1051, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1078, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1118, n1121, n1122,
         n1123, n1124, n1125, n1132, n1133, n1134, n1135, n1136, n1139, n1140,
         n1141, n1142, n1143, n1145, n1146, n1147, n1148, n1149, n1150, n1152,
         n1154, n1155, n1156, n1157, n1158, n1159, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1, n2, n3, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25,
         n27, n29, n31, n33, n37, n55, n73, n91, n109, n127, n145, n163, n181,
         n199, n217, n235, n253, n271, n289, n307, n325, n343, n361, n379,
         n397, n415, n433, n451, n469, n487, n505, n523, n541, n559, n577,
         n595, n596, n597, n599, n601, n603, n605, n607, n609, n611, n613,
         n615, n617, n619, n621, n623, n625, n627, n629, n631, n633, n635,
         n637, n639, n641, n643, n645, n647, n649, n651, n653, n655, n657,
         n659, n661, n664, n665, n667, n668, n695, n696, n724, n726, n727,
         n738, n739, n752, n753, n755, n756, n767, n768, n780, n782, n783,
         n794, n795, n807, n809, n810, n821, n822, n834, n836, n837, n848,
         n849, n861, n863, n864, n875, n876, n888, n890, n891, n902, n903,
         n915, n917, n918, n929, n930, n942, n944, n945, n956, n957, n969,
         n971, n972, n983, n984, n996, n998, n999, n1010, n1011, n1023, n1025,
         n1026, n1037, n1038, n1050, n1052, n1053, n1064, n1065, n1077, n1079,
         n1080, n1099, n1100, n1116, n1117, n1119, n1120, n1126, n1127, n1128,
         n1129, n1130, n1131, n1137, n1138, n1144, n1151, n1153, n1160, n1194,
         n1195, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580;
  assign N253 = \Addr<0> ;
  assign N254 = \Addr<1> ;
  assign N255 = \Addr<2> ;
  assign N256 = \Addr<3> ;
  assign N257 = \Addr<4> ;
  assign N258 = \Addr<5> ;
  assign CacheHit = 1'b0;

  DFFPOSX1 \rand_pat_reg<0>  ( .D(n1193), .CLK(clk), .Q(\rand_pat<0> ) );
  DFFPOSX1 \rand_pat_reg<31>  ( .D(n1192), .CLK(clk), .Q(\rand_pat<31> ) );
  DFFPOSX1 \rand_pat_reg<30>  ( .D(n1191), .CLK(clk), .Q(\rand_pat<30> ) );
  DFFPOSX1 \rand_pat_reg<29>  ( .D(n1190), .CLK(clk), .Q(\rand_pat<29> ) );
  DFFPOSX1 \rand_pat_reg<28>  ( .D(n1189), .CLK(clk), .Q(\rand_pat<28> ) );
  DFFPOSX1 \rand_pat_reg<27>  ( .D(n1188), .CLK(clk), .Q(\rand_pat<27> ) );
  DFFPOSX1 \rand_pat_reg<26>  ( .D(n1187), .CLK(clk), .Q(\rand_pat<26> ) );
  DFFPOSX1 \rand_pat_reg<25>  ( .D(n1186), .CLK(clk), .Q(\rand_pat<25> ) );
  DFFPOSX1 \rand_pat_reg<24>  ( .D(n1185), .CLK(clk), .Q(\rand_pat<24> ) );
  DFFPOSX1 \rand_pat_reg<23>  ( .D(n1184), .CLK(clk), .Q(\rand_pat<23> ) );
  DFFPOSX1 \rand_pat_reg<22>  ( .D(n1183), .CLK(clk), .Q(\rand_pat<22> ) );
  DFFPOSX1 \rand_pat_reg<21>  ( .D(n1182), .CLK(clk), .Q(\rand_pat<21> ) );
  DFFPOSX1 \rand_pat_reg<20>  ( .D(n1181), .CLK(clk), .Q(\rand_pat<20> ) );
  DFFPOSX1 \rand_pat_reg<19>  ( .D(n1180), .CLK(clk), .Q(\rand_pat<19> ) );
  DFFPOSX1 \rand_pat_reg<18>  ( .D(n1179), .CLK(clk), .Q(\rand_pat<18> ) );
  DFFPOSX1 \rand_pat_reg<17>  ( .D(n1178), .CLK(clk), .Q(\rand_pat<17> ) );
  DFFPOSX1 \rand_pat_reg<16>  ( .D(n1177), .CLK(clk), .Q(\rand_pat<16> ) );
  DFFPOSX1 \rand_pat_reg<15>  ( .D(n1176), .CLK(clk), .Q(\rand_pat<15> ) );
  DFFPOSX1 \rand_pat_reg<14>  ( .D(n1175), .CLK(clk), .Q(\rand_pat<14> ) );
  DFFPOSX1 \rand_pat_reg<13>  ( .D(n1174), .CLK(clk), .Q(\rand_pat<13> ) );
  DFFPOSX1 \rand_pat_reg<12>  ( .D(n1173), .CLK(clk), .Q(\rand_pat<12> ) );
  DFFPOSX1 \rand_pat_reg<11>  ( .D(n1172), .CLK(clk), .Q(\rand_pat<11> ) );
  DFFPOSX1 \rand_pat_reg<10>  ( .D(n1171), .CLK(clk), .Q(\rand_pat<10> ) );
  DFFPOSX1 \rand_pat_reg<9>  ( .D(n1170), .CLK(clk), .Q(\rand_pat<9> ) );
  DFFPOSX1 \rand_pat_reg<8>  ( .D(n1169), .CLK(clk), .Q(\rand_pat<8> ) );
  DFFPOSX1 \rand_pat_reg<7>  ( .D(n1168), .CLK(clk), .Q(\rand_pat<7> ) );
  DFFPOSX1 \rand_pat_reg<6>  ( .D(n1167), .CLK(clk), .Q(\rand_pat<6> ) );
  DFFPOSX1 \rand_pat_reg<5>  ( .D(n1166), .CLK(clk), .Q(\rand_pat<5> ) );
  DFFPOSX1 \rand_pat_reg<4>  ( .D(n1165), .CLK(clk), .Q(\rand_pat<4> ) );
  DFFPOSX1 \rand_pat_reg<3>  ( .D(n1164), .CLK(clk), .Q(\rand_pat<3> ) );
  DFFPOSX1 \rand_pat_reg<2>  ( .D(n1163), .CLK(clk), .Q(\rand_pat<2> ) );
  DFFPOSX1 \rand_pat_reg<1>  ( .D(n1162), .CLK(clk), .Q(\rand_pat<1> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1707), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1706), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1705), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1704), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1703), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1702), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1701), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1700), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1699), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1698), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1697), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1696), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1695), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1694), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1693), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1692), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1691), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1690), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1689), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1688), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1687), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1686), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1685), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1684), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1683), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1682), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1681), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1680), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1679), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1678), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1677), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1676), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1675), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1674), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1673), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1672), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1671), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1670), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1669), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1668), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1667), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1666), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1665), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1664), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1663), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1662), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1661), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1660), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1659), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1658), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1657), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1656), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1655), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1654), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1653), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1652), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1651), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1650), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1649), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1648), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1647), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1646), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1645), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1644), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1643), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1642), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1641), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1640), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1639), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1638), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1637), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1636), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1635), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1634), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1633), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1632), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1631), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1630), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1629), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1628), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1627), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1626), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1625), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1624), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1623), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1622), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1621), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1620), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1619), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1618), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1617), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1616), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1615), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1614), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1613), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1612), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1611), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1610), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1609), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1608), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1607), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1606), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1605), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1604), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1603), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1602), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1601), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1600), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1599), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1598), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1597), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1596), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1595), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1594), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1593), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1592), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1591), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1590), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1589), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1588), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1587), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1586), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1585), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1584), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1583), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1582), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1581), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1580), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1579), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1578), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1577), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1576), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1575), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1574), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1573), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1572), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1571), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1570), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1569), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1568), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1567), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1566), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1565), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1564), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1563), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1562), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1561), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1560), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1559), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1558), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1557), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1556), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1555), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1554), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1553), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1552), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1551), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1550), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1549), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1548), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1547), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1546), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1545), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1544), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1543), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1542), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1541), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1540), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1539), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1538), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1537), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1536), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1535), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1534), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1533), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1532), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1531), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1530), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1529), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1528), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1527), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1526), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1525), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1524), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1523), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1522), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1521), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1520), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1519), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1518), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1517), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1516), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1515), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1514), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1513), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1512), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1511), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1510), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1509), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1508), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1507), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1506), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1505), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1504), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1503), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1502), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1501), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1500), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1499), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1498), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1497), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1496), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1495), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1494), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1493), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1492), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1491), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1490), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1489), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1488), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1487), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1486), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1485), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1484), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1483), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1482), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1481), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1480), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1479), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1478), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1477), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1476), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1475), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1474), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1473), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1472), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1471), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1470), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1469), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1468), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1467), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1466), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1465), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1464), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1463), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1462), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1461), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1460), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1459), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1458), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1457), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1456), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1455), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1454), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1453), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1452), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1451), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1450), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1449), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1448), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1447), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1446), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1445), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1444), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n1443), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n1442), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n1441), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n1440), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n1439), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n1438), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n1437), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n1436), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n1435), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n1434), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n1433), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n1432), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n1431), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n1430), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n1429), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n1428), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n1427), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n1426), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n1425), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n1424), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n1423), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n1422), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n1421), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n1420), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n1419), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n1418), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n1417), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n1416), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n1415), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n1414), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n1413), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n1412), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n1411), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n1410), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n1409), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n1408), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n1407), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n1406), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n1405), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n1404), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n1403), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n1402), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n1401), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n1400), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n1399), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n1398), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n1397), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n1396), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n1395), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n1394), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n1393), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n1392), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n1391), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n1390), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n1389), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n1388), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n1387), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n1386), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n1385), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n1384), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n1383), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n1382), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n1381), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n1380), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n1379), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n1378), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n1377), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n1376), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n1375), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n1374), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n1373), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n1372), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n1371), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n1370), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n1369), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n1368), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n1367), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n1366), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n1365), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n1364), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n1363), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n1362), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n1361), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n1360), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n1359), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n1358), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n1357), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n1356), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n1355), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n1354), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n1353), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n1352), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n1351), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n1350), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n1349), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n1348), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n1347), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n1346), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n1345), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n1344), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n1343), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n1342), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n1341), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n1340), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n1339), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n1338), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n1337), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n1336), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n1335), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n1334), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n1333), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n1332), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n1331), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n1330), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n1329), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n1328), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n1327), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n1326), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n1325), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n1324), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n1323), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n1322), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n1321), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n1320), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n1319), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n1318), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n1317), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n1316), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n1315), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n1314), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n1313), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n1312), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n1311), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n1310), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n1309), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n1308), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n1307), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n1306), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n1305), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n1304), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n1303), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n1302), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n1301), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n1300), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n1299), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n1298), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n1297), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n1296), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n1295), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n1294), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n1293), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n1292), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n1291), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n1290), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n1289), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n1288), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n1287), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n1286), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n1285), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n1284), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n1283), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n1282), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n1281), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n1280), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n1279), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n1278), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n1277), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n1276), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n1275), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n1274), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n1273), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n1272), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n1271), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n1270), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n1269), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n1268), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n1267), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n1266), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n1265), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n1264), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n1263), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n1262), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n1261), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n1260), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n1259), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n1258), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n1257), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n1256), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n1255), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n1254), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n1253), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n1252), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n1251), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n1250), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n1249), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n1248), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n1247), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n1246), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n1245), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n1244), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n1243), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n1242), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n1241), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n1240), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n1239), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n1238), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n1237), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n1236), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n1235), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n1234), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n1233), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n1232), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n1231), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n1230), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n1229), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n1228), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n1227), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n1226), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n1225), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n1224), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n1223), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n1222), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n1221), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n1220), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n1219), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n1218), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n1217), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n1216), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n1215), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n1214), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n1213), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n1212), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n1211), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n1210), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n1209), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n1208), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n1207), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n1206), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n1205), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n1204), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n1203), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n1202), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n1201), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n1200), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n1199), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n1198), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n1197), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n1196), .CLK(clk), .Q(\mem<63><0> ) );
  OAI21X1 U3 ( .A(n2525), .B(n2449), .C(n4), .Y(n1196) );
  NAND2X1 U4 ( .A(\mem<63><0> ), .B(n2525), .Y(n4) );
  OAI21X1 U5 ( .A(n2525), .B(n2450), .C(n6), .Y(n1197) );
  NAND2X1 U6 ( .A(\mem<63><1> ), .B(n2525), .Y(n6) );
  OAI21X1 U7 ( .A(n2525), .B(n2451), .C(n8), .Y(n1198) );
  NAND2X1 U8 ( .A(\mem<63><2> ), .B(n2525), .Y(n8) );
  OAI21X1 U9 ( .A(n2525), .B(n2452), .C(n10), .Y(n1199) );
  NAND2X1 U10 ( .A(\mem<63><3> ), .B(n2524), .Y(n10) );
  OAI21X1 U11 ( .A(n2525), .B(n2453), .C(n12), .Y(n1200) );
  NAND2X1 U12 ( .A(\mem<63><4> ), .B(n2524), .Y(n12) );
  OAI21X1 U13 ( .A(n2525), .B(n2454), .C(n14), .Y(n1201) );
  NAND2X1 U14 ( .A(\mem<63><5> ), .B(n2524), .Y(n14) );
  OAI21X1 U15 ( .A(n2525), .B(n2455), .C(n16), .Y(n1202) );
  NAND2X1 U16 ( .A(\mem<63><6> ), .B(n2524), .Y(n16) );
  OAI21X1 U17 ( .A(n2525), .B(n2456), .C(n18), .Y(n1203) );
  NAND2X1 U18 ( .A(\mem<63><7> ), .B(n2524), .Y(n18) );
  OAI21X1 U19 ( .A(n2525), .B(n2457), .C(n20), .Y(n1204) );
  NAND2X1 U20 ( .A(\mem<62><0> ), .B(n2524), .Y(n20) );
  OAI21X1 U21 ( .A(n2525), .B(n2458), .C(n22), .Y(n1205) );
  NAND2X1 U22 ( .A(\mem<62><1> ), .B(n2524), .Y(n22) );
  OAI21X1 U23 ( .A(n2525), .B(n2459), .C(n24), .Y(n1206) );
  NAND2X1 U24 ( .A(\mem<62><2> ), .B(n2524), .Y(n24) );
  OAI21X1 U25 ( .A(n2525), .B(n2460), .C(n26), .Y(n1207) );
  NAND2X1 U26 ( .A(\mem<62><3> ), .B(n2524), .Y(n26) );
  OAI21X1 U27 ( .A(n2524), .B(n2461), .C(n28), .Y(n1208) );
  NAND2X1 U28 ( .A(\mem<62><4> ), .B(n2524), .Y(n28) );
  OAI21X1 U29 ( .A(n2524), .B(n2462), .C(n30), .Y(n1209) );
  NAND2X1 U30 ( .A(\mem<62><5> ), .B(n2524), .Y(n30) );
  OAI21X1 U31 ( .A(n2524), .B(n2463), .C(n32), .Y(n1210) );
  NAND2X1 U32 ( .A(\mem<62><6> ), .B(n2525), .Y(n32) );
  OAI21X1 U33 ( .A(n2524), .B(n2464), .C(n34), .Y(n1211) );
  NAND2X1 U34 ( .A(\mem<62><7> ), .B(n2525), .Y(n34) );
  OAI21X1 U36 ( .A(n2449), .B(n2520), .C(n38), .Y(n1212) );
  NAND2X1 U37 ( .A(\mem<61><0> ), .B(n2520), .Y(n38) );
  OAI21X1 U38 ( .A(n2450), .B(n2520), .C(n39), .Y(n1213) );
  NAND2X1 U39 ( .A(\mem<61><1> ), .B(n2520), .Y(n39) );
  OAI21X1 U40 ( .A(n2451), .B(n2520), .C(n40), .Y(n1214) );
  NAND2X1 U41 ( .A(\mem<61><2> ), .B(n2519), .Y(n40) );
  OAI21X1 U42 ( .A(n2452), .B(n2520), .C(n41), .Y(n1215) );
  NAND2X1 U43 ( .A(\mem<61><3> ), .B(n2519), .Y(n41) );
  OAI21X1 U44 ( .A(n2453), .B(n2520), .C(n42), .Y(n1216) );
  NAND2X1 U45 ( .A(\mem<61><4> ), .B(n2519), .Y(n42) );
  OAI21X1 U46 ( .A(n2454), .B(n2520), .C(n43), .Y(n1217) );
  NAND2X1 U47 ( .A(\mem<61><5> ), .B(n2519), .Y(n43) );
  OAI21X1 U48 ( .A(n2455), .B(n2520), .C(n44), .Y(n1218) );
  NAND2X1 U49 ( .A(\mem<61><6> ), .B(n2519), .Y(n44) );
  OAI21X1 U50 ( .A(n2456), .B(n2520), .C(n45), .Y(n1219) );
  NAND2X1 U51 ( .A(\mem<61><7> ), .B(n2519), .Y(n45) );
  OAI21X1 U52 ( .A(n2457), .B(n2520), .C(n46), .Y(n1220) );
  NAND2X1 U53 ( .A(\mem<60><0> ), .B(n2519), .Y(n46) );
  OAI21X1 U54 ( .A(n2458), .B(n2520), .C(n47), .Y(n1221) );
  NAND2X1 U55 ( .A(\mem<60><1> ), .B(n2519), .Y(n47) );
  OAI21X1 U56 ( .A(n2459), .B(n2520), .C(n48), .Y(n1222) );
  NAND2X1 U57 ( .A(\mem<60><2> ), .B(n2519), .Y(n48) );
  OAI21X1 U58 ( .A(n2460), .B(n2520), .C(n49), .Y(n1223) );
  NAND2X1 U59 ( .A(\mem<60><3> ), .B(n2519), .Y(n49) );
  OAI21X1 U60 ( .A(n2461), .B(n2519), .C(n50), .Y(n1224) );
  NAND2X1 U61 ( .A(\mem<60><4> ), .B(n2519), .Y(n50) );
  OAI21X1 U62 ( .A(n2462), .B(n2519), .C(n51), .Y(n1225) );
  NAND2X1 U63 ( .A(\mem<60><5> ), .B(n2519), .Y(n51) );
  OAI21X1 U64 ( .A(n2463), .B(n2519), .C(n52), .Y(n1226) );
  NAND2X1 U65 ( .A(\mem<60><6> ), .B(n2520), .Y(n52) );
  OAI21X1 U66 ( .A(n2464), .B(n2519), .C(n53), .Y(n1227) );
  NAND2X1 U67 ( .A(\mem<60><7> ), .B(n2520), .Y(n53) );
  OAI21X1 U69 ( .A(n2449), .B(n2518), .C(n56), .Y(n1228) );
  NAND2X1 U70 ( .A(\mem<59><0> ), .B(n2518), .Y(n56) );
  OAI21X1 U71 ( .A(n2450), .B(n2518), .C(n57), .Y(n1229) );
  NAND2X1 U72 ( .A(\mem<59><1> ), .B(n2518), .Y(n57) );
  OAI21X1 U73 ( .A(n2451), .B(n2518), .C(n58), .Y(n1230) );
  NAND2X1 U74 ( .A(\mem<59><2> ), .B(n2517), .Y(n58) );
  OAI21X1 U75 ( .A(n2452), .B(n2518), .C(n59), .Y(n1231) );
  NAND2X1 U76 ( .A(\mem<59><3> ), .B(n2517), .Y(n59) );
  OAI21X1 U77 ( .A(n2453), .B(n2518), .C(n60), .Y(n1232) );
  NAND2X1 U78 ( .A(\mem<59><4> ), .B(n2517), .Y(n60) );
  OAI21X1 U79 ( .A(n2454), .B(n2518), .C(n61), .Y(n1233) );
  NAND2X1 U80 ( .A(\mem<59><5> ), .B(n2517), .Y(n61) );
  OAI21X1 U81 ( .A(n2455), .B(n2518), .C(n62), .Y(n1234) );
  NAND2X1 U82 ( .A(\mem<59><6> ), .B(n2517), .Y(n62) );
  OAI21X1 U83 ( .A(n2456), .B(n2518), .C(n63), .Y(n1235) );
  NAND2X1 U84 ( .A(\mem<59><7> ), .B(n2517), .Y(n63) );
  OAI21X1 U85 ( .A(n2457), .B(n2518), .C(n64), .Y(n1236) );
  NAND2X1 U86 ( .A(\mem<58><0> ), .B(n2517), .Y(n64) );
  OAI21X1 U87 ( .A(n2458), .B(n2518), .C(n65), .Y(n1237) );
  NAND2X1 U88 ( .A(\mem<58><1> ), .B(n2517), .Y(n65) );
  OAI21X1 U89 ( .A(n2459), .B(n2518), .C(n66), .Y(n1238) );
  NAND2X1 U90 ( .A(\mem<58><2> ), .B(n2517), .Y(n66) );
  OAI21X1 U91 ( .A(n2460), .B(n2518), .C(n67), .Y(n1239) );
  NAND2X1 U92 ( .A(\mem<58><3> ), .B(n2517), .Y(n67) );
  OAI21X1 U93 ( .A(n2461), .B(n2517), .C(n68), .Y(n1240) );
  NAND2X1 U94 ( .A(\mem<58><4> ), .B(n2517), .Y(n68) );
  OAI21X1 U95 ( .A(n2462), .B(n2517), .C(n69), .Y(n1241) );
  NAND2X1 U96 ( .A(\mem<58><5> ), .B(n2517), .Y(n69) );
  OAI21X1 U97 ( .A(n2463), .B(n2517), .C(n70), .Y(n1242) );
  NAND2X1 U98 ( .A(\mem<58><6> ), .B(n2518), .Y(n70) );
  OAI21X1 U99 ( .A(n2464), .B(n2517), .C(n71), .Y(n1243) );
  NAND2X1 U100 ( .A(\mem<58><7> ), .B(n2518), .Y(n71) );
  OAI21X1 U102 ( .A(n2449), .B(n2516), .C(n74), .Y(n1244) );
  NAND2X1 U103 ( .A(\mem<57><0> ), .B(n2516), .Y(n74) );
  OAI21X1 U104 ( .A(n2450), .B(n2516), .C(n75), .Y(n1245) );
  NAND2X1 U105 ( .A(\mem<57><1> ), .B(n2516), .Y(n75) );
  OAI21X1 U106 ( .A(n2451), .B(n2516), .C(n76), .Y(n1246) );
  NAND2X1 U107 ( .A(\mem<57><2> ), .B(n2515), .Y(n76) );
  OAI21X1 U108 ( .A(n2452), .B(n2516), .C(n77), .Y(n1247) );
  NAND2X1 U109 ( .A(\mem<57><3> ), .B(n2515), .Y(n77) );
  OAI21X1 U110 ( .A(n2453), .B(n2516), .C(n78), .Y(n1248) );
  NAND2X1 U111 ( .A(\mem<57><4> ), .B(n2515), .Y(n78) );
  OAI21X1 U112 ( .A(n2454), .B(n2516), .C(n79), .Y(n1249) );
  NAND2X1 U113 ( .A(\mem<57><5> ), .B(n2515), .Y(n79) );
  OAI21X1 U114 ( .A(n2455), .B(n2516), .C(n80), .Y(n1250) );
  NAND2X1 U115 ( .A(\mem<57><6> ), .B(n2515), .Y(n80) );
  OAI21X1 U116 ( .A(n2456), .B(n2516), .C(n81), .Y(n1251) );
  NAND2X1 U117 ( .A(\mem<57><7> ), .B(n2515), .Y(n81) );
  OAI21X1 U118 ( .A(n2457), .B(n2516), .C(n82), .Y(n1252) );
  NAND2X1 U119 ( .A(\mem<56><0> ), .B(n2515), .Y(n82) );
  OAI21X1 U120 ( .A(n2458), .B(n2516), .C(n83), .Y(n1253) );
  NAND2X1 U121 ( .A(\mem<56><1> ), .B(n2515), .Y(n83) );
  OAI21X1 U122 ( .A(n2459), .B(n2516), .C(n84), .Y(n1254) );
  NAND2X1 U123 ( .A(\mem<56><2> ), .B(n2515), .Y(n84) );
  OAI21X1 U124 ( .A(n2460), .B(n2516), .C(n85), .Y(n1255) );
  NAND2X1 U125 ( .A(\mem<56><3> ), .B(n2515), .Y(n85) );
  OAI21X1 U126 ( .A(n2461), .B(n2515), .C(n86), .Y(n1256) );
  NAND2X1 U127 ( .A(\mem<56><4> ), .B(n2515), .Y(n86) );
  OAI21X1 U128 ( .A(n2462), .B(n2515), .C(n87), .Y(n1257) );
  NAND2X1 U129 ( .A(\mem<56><5> ), .B(n2515), .Y(n87) );
  OAI21X1 U130 ( .A(n2463), .B(n2515), .C(n88), .Y(n1258) );
  NAND2X1 U131 ( .A(\mem<56><6> ), .B(n2516), .Y(n88) );
  OAI21X1 U132 ( .A(n2464), .B(n2515), .C(n89), .Y(n1259) );
  NAND2X1 U133 ( .A(\mem<56><7> ), .B(n2516), .Y(n89) );
  OAI21X1 U135 ( .A(n2449), .B(n2514), .C(n92), .Y(n1260) );
  NAND2X1 U136 ( .A(\mem<55><0> ), .B(n2514), .Y(n92) );
  OAI21X1 U137 ( .A(n2450), .B(n2514), .C(n93), .Y(n1261) );
  NAND2X1 U138 ( .A(\mem<55><1> ), .B(n2514), .Y(n93) );
  OAI21X1 U139 ( .A(n2451), .B(n2514), .C(n94), .Y(n1262) );
  NAND2X1 U140 ( .A(\mem<55><2> ), .B(n2513), .Y(n94) );
  OAI21X1 U141 ( .A(n2452), .B(n2514), .C(n95), .Y(n1263) );
  NAND2X1 U142 ( .A(\mem<55><3> ), .B(n2513), .Y(n95) );
  OAI21X1 U143 ( .A(n2453), .B(n2514), .C(n96), .Y(n1264) );
  NAND2X1 U144 ( .A(\mem<55><4> ), .B(n2513), .Y(n96) );
  OAI21X1 U145 ( .A(n2454), .B(n2514), .C(n97), .Y(n1265) );
  NAND2X1 U146 ( .A(\mem<55><5> ), .B(n2513), .Y(n97) );
  OAI21X1 U147 ( .A(n2455), .B(n2514), .C(n98), .Y(n1266) );
  NAND2X1 U148 ( .A(\mem<55><6> ), .B(n2513), .Y(n98) );
  OAI21X1 U149 ( .A(n2456), .B(n2514), .C(n99), .Y(n1267) );
  NAND2X1 U150 ( .A(\mem<55><7> ), .B(n2513), .Y(n99) );
  OAI21X1 U151 ( .A(n2457), .B(n2514), .C(n100), .Y(n1268) );
  NAND2X1 U152 ( .A(\mem<54><0> ), .B(n2513), .Y(n100) );
  OAI21X1 U153 ( .A(n2458), .B(n2514), .C(n101), .Y(n1269) );
  NAND2X1 U154 ( .A(\mem<54><1> ), .B(n2513), .Y(n101) );
  OAI21X1 U155 ( .A(n2459), .B(n2514), .C(n102), .Y(n1270) );
  NAND2X1 U156 ( .A(\mem<54><2> ), .B(n2513), .Y(n102) );
  OAI21X1 U157 ( .A(n2460), .B(n2514), .C(n103), .Y(n1271) );
  NAND2X1 U158 ( .A(\mem<54><3> ), .B(n2513), .Y(n103) );
  OAI21X1 U159 ( .A(n2461), .B(n2513), .C(n104), .Y(n1272) );
  NAND2X1 U160 ( .A(\mem<54><4> ), .B(n2513), .Y(n104) );
  OAI21X1 U161 ( .A(n2462), .B(n2513), .C(n105), .Y(n1273) );
  NAND2X1 U162 ( .A(\mem<54><5> ), .B(n2513), .Y(n105) );
  OAI21X1 U163 ( .A(n2463), .B(n2513), .C(n106), .Y(n1274) );
  NAND2X1 U164 ( .A(\mem<54><6> ), .B(n2514), .Y(n106) );
  OAI21X1 U165 ( .A(n2464), .B(n2513), .C(n107), .Y(n1275) );
  NAND2X1 U166 ( .A(\mem<54><7> ), .B(n2514), .Y(n107) );
  OAI21X1 U168 ( .A(n2449), .B(n2512), .C(n110), .Y(n1276) );
  NAND2X1 U169 ( .A(\mem<53><0> ), .B(n2512), .Y(n110) );
  OAI21X1 U170 ( .A(n2450), .B(n2512), .C(n111), .Y(n1277) );
  NAND2X1 U171 ( .A(\mem<53><1> ), .B(n2512), .Y(n111) );
  OAI21X1 U172 ( .A(n2451), .B(n2512), .C(n112), .Y(n1278) );
  NAND2X1 U173 ( .A(\mem<53><2> ), .B(n2511), .Y(n112) );
  OAI21X1 U174 ( .A(n2452), .B(n2512), .C(n113), .Y(n1279) );
  NAND2X1 U175 ( .A(\mem<53><3> ), .B(n2511), .Y(n113) );
  OAI21X1 U176 ( .A(n2453), .B(n2512), .C(n114), .Y(n1280) );
  NAND2X1 U177 ( .A(\mem<53><4> ), .B(n2511), .Y(n114) );
  OAI21X1 U178 ( .A(n2454), .B(n2512), .C(n115), .Y(n1281) );
  NAND2X1 U179 ( .A(\mem<53><5> ), .B(n2511), .Y(n115) );
  OAI21X1 U180 ( .A(n2455), .B(n2512), .C(n116), .Y(n1282) );
  NAND2X1 U181 ( .A(\mem<53><6> ), .B(n2511), .Y(n116) );
  OAI21X1 U182 ( .A(n2456), .B(n2512), .C(n117), .Y(n1283) );
  NAND2X1 U183 ( .A(\mem<53><7> ), .B(n2511), .Y(n117) );
  OAI21X1 U184 ( .A(n2457), .B(n2512), .C(n118), .Y(n1284) );
  NAND2X1 U185 ( .A(\mem<52><0> ), .B(n2511), .Y(n118) );
  OAI21X1 U186 ( .A(n2458), .B(n2512), .C(n119), .Y(n1285) );
  NAND2X1 U187 ( .A(\mem<52><1> ), .B(n2511), .Y(n119) );
  OAI21X1 U188 ( .A(n2459), .B(n2512), .C(n120), .Y(n1286) );
  NAND2X1 U189 ( .A(\mem<52><2> ), .B(n2511), .Y(n120) );
  OAI21X1 U190 ( .A(n2460), .B(n2512), .C(n121), .Y(n1287) );
  NAND2X1 U191 ( .A(\mem<52><3> ), .B(n2511), .Y(n121) );
  OAI21X1 U192 ( .A(n2461), .B(n2511), .C(n122), .Y(n1288) );
  NAND2X1 U193 ( .A(\mem<52><4> ), .B(n2511), .Y(n122) );
  OAI21X1 U194 ( .A(n2462), .B(n2511), .C(n123), .Y(n1289) );
  NAND2X1 U195 ( .A(\mem<52><5> ), .B(n2511), .Y(n123) );
  OAI21X1 U196 ( .A(n2463), .B(n2511), .C(n124), .Y(n1290) );
  NAND2X1 U197 ( .A(\mem<52><6> ), .B(n2512), .Y(n124) );
  OAI21X1 U198 ( .A(n2464), .B(n2511), .C(n125), .Y(n1291) );
  NAND2X1 U199 ( .A(\mem<52><7> ), .B(n2512), .Y(n125) );
  OAI21X1 U201 ( .A(n2449), .B(n2510), .C(n128), .Y(n1292) );
  NAND2X1 U202 ( .A(\mem<51><0> ), .B(n2510), .Y(n128) );
  OAI21X1 U203 ( .A(n2450), .B(n2510), .C(n129), .Y(n1293) );
  NAND2X1 U204 ( .A(\mem<51><1> ), .B(n2510), .Y(n129) );
  OAI21X1 U205 ( .A(n2451), .B(n2510), .C(n130), .Y(n1294) );
  NAND2X1 U206 ( .A(\mem<51><2> ), .B(n2509), .Y(n130) );
  OAI21X1 U207 ( .A(n2452), .B(n2510), .C(n131), .Y(n1295) );
  NAND2X1 U208 ( .A(\mem<51><3> ), .B(n2509), .Y(n131) );
  OAI21X1 U209 ( .A(n2453), .B(n2510), .C(n132), .Y(n1296) );
  NAND2X1 U210 ( .A(\mem<51><4> ), .B(n2509), .Y(n132) );
  OAI21X1 U211 ( .A(n2454), .B(n2510), .C(n133), .Y(n1297) );
  NAND2X1 U212 ( .A(\mem<51><5> ), .B(n2509), .Y(n133) );
  OAI21X1 U213 ( .A(n2455), .B(n2510), .C(n134), .Y(n1298) );
  NAND2X1 U214 ( .A(\mem<51><6> ), .B(n2509), .Y(n134) );
  OAI21X1 U215 ( .A(n2456), .B(n2510), .C(n135), .Y(n1299) );
  NAND2X1 U216 ( .A(\mem<51><7> ), .B(n2509), .Y(n135) );
  OAI21X1 U217 ( .A(n2457), .B(n2510), .C(n136), .Y(n1300) );
  NAND2X1 U218 ( .A(\mem<50><0> ), .B(n2509), .Y(n136) );
  OAI21X1 U219 ( .A(n2458), .B(n2510), .C(n137), .Y(n1301) );
  NAND2X1 U220 ( .A(\mem<50><1> ), .B(n2509), .Y(n137) );
  OAI21X1 U221 ( .A(n2459), .B(n2510), .C(n138), .Y(n1302) );
  NAND2X1 U222 ( .A(\mem<50><2> ), .B(n2509), .Y(n138) );
  OAI21X1 U223 ( .A(n2460), .B(n2510), .C(n139), .Y(n1303) );
  NAND2X1 U224 ( .A(\mem<50><3> ), .B(n2509), .Y(n139) );
  OAI21X1 U225 ( .A(n2461), .B(n2509), .C(n140), .Y(n1304) );
  NAND2X1 U226 ( .A(\mem<50><4> ), .B(n2509), .Y(n140) );
  OAI21X1 U227 ( .A(n2462), .B(n2509), .C(n141), .Y(n1305) );
  NAND2X1 U228 ( .A(\mem<50><5> ), .B(n2509), .Y(n141) );
  OAI21X1 U229 ( .A(n2463), .B(n2509), .C(n142), .Y(n1306) );
  NAND2X1 U230 ( .A(\mem<50><6> ), .B(n2510), .Y(n142) );
  OAI21X1 U231 ( .A(n2464), .B(n2509), .C(n143), .Y(n1307) );
  NAND2X1 U232 ( .A(\mem<50><7> ), .B(n2510), .Y(n143) );
  OAI21X1 U234 ( .A(n2449), .B(n2508), .C(n146), .Y(n1308) );
  NAND2X1 U235 ( .A(\mem<49><0> ), .B(n2508), .Y(n146) );
  OAI21X1 U236 ( .A(n2450), .B(n2508), .C(n147), .Y(n1309) );
  NAND2X1 U237 ( .A(\mem<49><1> ), .B(n2508), .Y(n147) );
  OAI21X1 U238 ( .A(n2451), .B(n2508), .C(n148), .Y(n1310) );
  NAND2X1 U239 ( .A(\mem<49><2> ), .B(n2507), .Y(n148) );
  OAI21X1 U240 ( .A(n2452), .B(n2508), .C(n149), .Y(n1311) );
  NAND2X1 U241 ( .A(\mem<49><3> ), .B(n2507), .Y(n149) );
  OAI21X1 U242 ( .A(n2453), .B(n2508), .C(n150), .Y(n1312) );
  NAND2X1 U243 ( .A(\mem<49><4> ), .B(n2507), .Y(n150) );
  OAI21X1 U244 ( .A(n2454), .B(n2508), .C(n151), .Y(n1313) );
  NAND2X1 U245 ( .A(\mem<49><5> ), .B(n2507), .Y(n151) );
  OAI21X1 U246 ( .A(n2455), .B(n2508), .C(n152), .Y(n1314) );
  NAND2X1 U247 ( .A(\mem<49><6> ), .B(n2507), .Y(n152) );
  OAI21X1 U248 ( .A(n2456), .B(n2508), .C(n153), .Y(n1315) );
  NAND2X1 U249 ( .A(\mem<49><7> ), .B(n2507), .Y(n153) );
  OAI21X1 U250 ( .A(n2457), .B(n2508), .C(n154), .Y(n1316) );
  NAND2X1 U251 ( .A(\mem<48><0> ), .B(n2507), .Y(n154) );
  OAI21X1 U252 ( .A(n2458), .B(n2508), .C(n155), .Y(n1317) );
  NAND2X1 U253 ( .A(\mem<48><1> ), .B(n2507), .Y(n155) );
  OAI21X1 U254 ( .A(n2459), .B(n2508), .C(n156), .Y(n1318) );
  NAND2X1 U255 ( .A(\mem<48><2> ), .B(n2507), .Y(n156) );
  OAI21X1 U256 ( .A(n2460), .B(n2508), .C(n157), .Y(n1319) );
  NAND2X1 U257 ( .A(\mem<48><3> ), .B(n2507), .Y(n157) );
  OAI21X1 U258 ( .A(n2461), .B(n2507), .C(n158), .Y(n1320) );
  NAND2X1 U259 ( .A(\mem<48><4> ), .B(n2507), .Y(n158) );
  OAI21X1 U260 ( .A(n2462), .B(n2507), .C(n159), .Y(n1321) );
  NAND2X1 U261 ( .A(\mem<48><5> ), .B(n2507), .Y(n159) );
  OAI21X1 U262 ( .A(n2463), .B(n2507), .C(n160), .Y(n1322) );
  NAND2X1 U263 ( .A(\mem<48><6> ), .B(n2508), .Y(n160) );
  OAI21X1 U264 ( .A(n2464), .B(n2507), .C(n161), .Y(n1323) );
  NAND2X1 U265 ( .A(\mem<48><7> ), .B(n2508), .Y(n161) );
  OAI21X1 U267 ( .A(n2449), .B(n2506), .C(n164), .Y(n1324) );
  NAND2X1 U268 ( .A(\mem<47><0> ), .B(n2506), .Y(n164) );
  OAI21X1 U269 ( .A(n2450), .B(n2506), .C(n165), .Y(n1325) );
  NAND2X1 U270 ( .A(\mem<47><1> ), .B(n2506), .Y(n165) );
  OAI21X1 U271 ( .A(n2451), .B(n2506), .C(n166), .Y(n1326) );
  NAND2X1 U272 ( .A(\mem<47><2> ), .B(n2505), .Y(n166) );
  OAI21X1 U273 ( .A(n2452), .B(n2506), .C(n167), .Y(n1327) );
  NAND2X1 U274 ( .A(\mem<47><3> ), .B(n2505), .Y(n167) );
  OAI21X1 U275 ( .A(n2453), .B(n2506), .C(n168), .Y(n1328) );
  NAND2X1 U276 ( .A(\mem<47><4> ), .B(n2505), .Y(n168) );
  OAI21X1 U277 ( .A(n2454), .B(n2506), .C(n169), .Y(n1329) );
  NAND2X1 U278 ( .A(\mem<47><5> ), .B(n2505), .Y(n169) );
  OAI21X1 U279 ( .A(n2455), .B(n2506), .C(n170), .Y(n1330) );
  NAND2X1 U280 ( .A(\mem<47><6> ), .B(n2505), .Y(n170) );
  OAI21X1 U281 ( .A(n2456), .B(n2506), .C(n171), .Y(n1331) );
  NAND2X1 U282 ( .A(\mem<47><7> ), .B(n2505), .Y(n171) );
  OAI21X1 U283 ( .A(n2457), .B(n2506), .C(n172), .Y(n1332) );
  NAND2X1 U284 ( .A(\mem<46><0> ), .B(n2505), .Y(n172) );
  OAI21X1 U285 ( .A(n2458), .B(n2506), .C(n173), .Y(n1333) );
  NAND2X1 U286 ( .A(\mem<46><1> ), .B(n2505), .Y(n173) );
  OAI21X1 U287 ( .A(n2459), .B(n2506), .C(n174), .Y(n1334) );
  NAND2X1 U288 ( .A(\mem<46><2> ), .B(n2505), .Y(n174) );
  OAI21X1 U289 ( .A(n2460), .B(n2506), .C(n175), .Y(n1335) );
  NAND2X1 U290 ( .A(\mem<46><3> ), .B(n2505), .Y(n175) );
  OAI21X1 U291 ( .A(n2461), .B(n2505), .C(n176), .Y(n1336) );
  NAND2X1 U292 ( .A(\mem<46><4> ), .B(n2505), .Y(n176) );
  OAI21X1 U293 ( .A(n2462), .B(n2505), .C(n177), .Y(n1337) );
  NAND2X1 U294 ( .A(\mem<46><5> ), .B(n2505), .Y(n177) );
  OAI21X1 U295 ( .A(n2463), .B(n2505), .C(n178), .Y(n1338) );
  NAND2X1 U296 ( .A(\mem<46><6> ), .B(n2506), .Y(n178) );
  OAI21X1 U297 ( .A(n2464), .B(n2505), .C(n179), .Y(n1339) );
  NAND2X1 U298 ( .A(\mem<46><7> ), .B(n2506), .Y(n179) );
  OAI21X1 U300 ( .A(n2449), .B(n2504), .C(n182), .Y(n1340) );
  NAND2X1 U301 ( .A(\mem<45><0> ), .B(n2504), .Y(n182) );
  OAI21X1 U302 ( .A(n2450), .B(n2504), .C(n183), .Y(n1341) );
  NAND2X1 U303 ( .A(\mem<45><1> ), .B(n2504), .Y(n183) );
  OAI21X1 U304 ( .A(n2451), .B(n2504), .C(n184), .Y(n1342) );
  NAND2X1 U305 ( .A(\mem<45><2> ), .B(n2503), .Y(n184) );
  OAI21X1 U306 ( .A(n2452), .B(n2504), .C(n185), .Y(n1343) );
  NAND2X1 U307 ( .A(\mem<45><3> ), .B(n2503), .Y(n185) );
  OAI21X1 U308 ( .A(n2453), .B(n2504), .C(n186), .Y(n1344) );
  NAND2X1 U309 ( .A(\mem<45><4> ), .B(n2503), .Y(n186) );
  OAI21X1 U310 ( .A(n2454), .B(n2504), .C(n187), .Y(n1345) );
  NAND2X1 U311 ( .A(\mem<45><5> ), .B(n2503), .Y(n187) );
  OAI21X1 U312 ( .A(n2455), .B(n2504), .C(n188), .Y(n1346) );
  NAND2X1 U313 ( .A(\mem<45><6> ), .B(n2503), .Y(n188) );
  OAI21X1 U314 ( .A(n2456), .B(n2504), .C(n189), .Y(n1347) );
  NAND2X1 U315 ( .A(\mem<45><7> ), .B(n2503), .Y(n189) );
  OAI21X1 U316 ( .A(n2457), .B(n2504), .C(n190), .Y(n1348) );
  NAND2X1 U317 ( .A(\mem<44><0> ), .B(n2503), .Y(n190) );
  OAI21X1 U318 ( .A(n2458), .B(n2504), .C(n191), .Y(n1349) );
  NAND2X1 U319 ( .A(\mem<44><1> ), .B(n2503), .Y(n191) );
  OAI21X1 U320 ( .A(n2459), .B(n2504), .C(n192), .Y(n1350) );
  NAND2X1 U321 ( .A(\mem<44><2> ), .B(n2503), .Y(n192) );
  OAI21X1 U322 ( .A(n2460), .B(n2504), .C(n193), .Y(n1351) );
  NAND2X1 U323 ( .A(\mem<44><3> ), .B(n2503), .Y(n193) );
  OAI21X1 U324 ( .A(n2461), .B(n2503), .C(n194), .Y(n1352) );
  NAND2X1 U325 ( .A(\mem<44><4> ), .B(n2503), .Y(n194) );
  OAI21X1 U326 ( .A(n2462), .B(n2503), .C(n195), .Y(n1353) );
  NAND2X1 U327 ( .A(\mem<44><5> ), .B(n2503), .Y(n195) );
  OAI21X1 U328 ( .A(n2463), .B(n2503), .C(n196), .Y(n1354) );
  NAND2X1 U329 ( .A(\mem<44><6> ), .B(n2504), .Y(n196) );
  OAI21X1 U330 ( .A(n2464), .B(n2503), .C(n197), .Y(n1355) );
  NAND2X1 U331 ( .A(\mem<44><7> ), .B(n2504), .Y(n197) );
  OAI21X1 U333 ( .A(n2449), .B(n2502), .C(n200), .Y(n1356) );
  NAND2X1 U334 ( .A(\mem<43><0> ), .B(n2502), .Y(n200) );
  OAI21X1 U335 ( .A(n2450), .B(n2502), .C(n201), .Y(n1357) );
  NAND2X1 U336 ( .A(\mem<43><1> ), .B(n2502), .Y(n201) );
  OAI21X1 U337 ( .A(n2451), .B(n2502), .C(n202), .Y(n1358) );
  NAND2X1 U338 ( .A(\mem<43><2> ), .B(n2501), .Y(n202) );
  OAI21X1 U339 ( .A(n2452), .B(n2502), .C(n203), .Y(n1359) );
  NAND2X1 U340 ( .A(\mem<43><3> ), .B(n2501), .Y(n203) );
  OAI21X1 U341 ( .A(n2453), .B(n2502), .C(n204), .Y(n1360) );
  NAND2X1 U342 ( .A(\mem<43><4> ), .B(n2501), .Y(n204) );
  OAI21X1 U343 ( .A(n2454), .B(n2502), .C(n205), .Y(n1361) );
  NAND2X1 U344 ( .A(\mem<43><5> ), .B(n2501), .Y(n205) );
  OAI21X1 U345 ( .A(n2455), .B(n2502), .C(n206), .Y(n1362) );
  NAND2X1 U346 ( .A(\mem<43><6> ), .B(n2501), .Y(n206) );
  OAI21X1 U347 ( .A(n2456), .B(n2502), .C(n207), .Y(n1363) );
  NAND2X1 U348 ( .A(\mem<43><7> ), .B(n2501), .Y(n207) );
  OAI21X1 U349 ( .A(n2457), .B(n2502), .C(n208), .Y(n1364) );
  NAND2X1 U350 ( .A(\mem<42><0> ), .B(n2501), .Y(n208) );
  OAI21X1 U351 ( .A(n2458), .B(n2502), .C(n209), .Y(n1365) );
  NAND2X1 U352 ( .A(\mem<42><1> ), .B(n2501), .Y(n209) );
  OAI21X1 U353 ( .A(n2459), .B(n2502), .C(n210), .Y(n1366) );
  NAND2X1 U354 ( .A(\mem<42><2> ), .B(n2501), .Y(n210) );
  OAI21X1 U355 ( .A(n2460), .B(n2502), .C(n211), .Y(n1367) );
  NAND2X1 U356 ( .A(\mem<42><3> ), .B(n2501), .Y(n211) );
  OAI21X1 U357 ( .A(n2461), .B(n2501), .C(n212), .Y(n1368) );
  NAND2X1 U358 ( .A(\mem<42><4> ), .B(n2501), .Y(n212) );
  OAI21X1 U359 ( .A(n2462), .B(n2501), .C(n213), .Y(n1369) );
  NAND2X1 U360 ( .A(\mem<42><5> ), .B(n2501), .Y(n213) );
  OAI21X1 U361 ( .A(n2463), .B(n2501), .C(n214), .Y(n1370) );
  NAND2X1 U362 ( .A(\mem<42><6> ), .B(n2502), .Y(n214) );
  OAI21X1 U363 ( .A(n2464), .B(n2501), .C(n215), .Y(n1371) );
  NAND2X1 U364 ( .A(\mem<42><7> ), .B(n2502), .Y(n215) );
  OAI21X1 U366 ( .A(n2449), .B(n2500), .C(n218), .Y(n1372) );
  NAND2X1 U367 ( .A(\mem<41><0> ), .B(n2500), .Y(n218) );
  OAI21X1 U368 ( .A(n2450), .B(n2500), .C(n219), .Y(n1373) );
  NAND2X1 U369 ( .A(\mem<41><1> ), .B(n2500), .Y(n219) );
  OAI21X1 U370 ( .A(n2451), .B(n2500), .C(n220), .Y(n1374) );
  NAND2X1 U371 ( .A(\mem<41><2> ), .B(n2499), .Y(n220) );
  OAI21X1 U372 ( .A(n2452), .B(n2500), .C(n221), .Y(n1375) );
  NAND2X1 U373 ( .A(\mem<41><3> ), .B(n2499), .Y(n221) );
  OAI21X1 U374 ( .A(n2453), .B(n2500), .C(n222), .Y(n1376) );
  NAND2X1 U375 ( .A(\mem<41><4> ), .B(n2499), .Y(n222) );
  OAI21X1 U376 ( .A(n2454), .B(n2500), .C(n223), .Y(n1377) );
  NAND2X1 U377 ( .A(\mem<41><5> ), .B(n2499), .Y(n223) );
  OAI21X1 U378 ( .A(n2455), .B(n2500), .C(n224), .Y(n1378) );
  NAND2X1 U379 ( .A(\mem<41><6> ), .B(n2499), .Y(n224) );
  OAI21X1 U380 ( .A(n2456), .B(n2500), .C(n225), .Y(n1379) );
  NAND2X1 U381 ( .A(\mem<41><7> ), .B(n2499), .Y(n225) );
  OAI21X1 U382 ( .A(n2457), .B(n2500), .C(n226), .Y(n1380) );
  NAND2X1 U383 ( .A(\mem<40><0> ), .B(n2499), .Y(n226) );
  OAI21X1 U384 ( .A(n2458), .B(n2500), .C(n227), .Y(n1381) );
  NAND2X1 U385 ( .A(\mem<40><1> ), .B(n2499), .Y(n227) );
  OAI21X1 U386 ( .A(n2459), .B(n2500), .C(n228), .Y(n1382) );
  NAND2X1 U387 ( .A(\mem<40><2> ), .B(n2499), .Y(n228) );
  OAI21X1 U388 ( .A(n2460), .B(n2500), .C(n229), .Y(n1383) );
  NAND2X1 U389 ( .A(\mem<40><3> ), .B(n2499), .Y(n229) );
  OAI21X1 U390 ( .A(n2461), .B(n2499), .C(n230), .Y(n1384) );
  NAND2X1 U391 ( .A(\mem<40><4> ), .B(n2499), .Y(n230) );
  OAI21X1 U392 ( .A(n2462), .B(n2499), .C(n231), .Y(n1385) );
  NAND2X1 U393 ( .A(\mem<40><5> ), .B(n2499), .Y(n231) );
  OAI21X1 U394 ( .A(n2463), .B(n2499), .C(n232), .Y(n1386) );
  NAND2X1 U395 ( .A(\mem<40><6> ), .B(n2500), .Y(n232) );
  OAI21X1 U396 ( .A(n2464), .B(n2499), .C(n233), .Y(n1387) );
  NAND2X1 U397 ( .A(\mem<40><7> ), .B(n2500), .Y(n233) );
  OAI21X1 U399 ( .A(n2449), .B(n2498), .C(n236), .Y(n1388) );
  NAND2X1 U400 ( .A(\mem<39><0> ), .B(n2498), .Y(n236) );
  OAI21X1 U401 ( .A(n2450), .B(n2498), .C(n237), .Y(n1389) );
  NAND2X1 U402 ( .A(\mem<39><1> ), .B(n2498), .Y(n237) );
  OAI21X1 U403 ( .A(n2451), .B(n2498), .C(n238), .Y(n1390) );
  NAND2X1 U404 ( .A(\mem<39><2> ), .B(n2497), .Y(n238) );
  OAI21X1 U405 ( .A(n2452), .B(n2498), .C(n239), .Y(n1391) );
  NAND2X1 U406 ( .A(\mem<39><3> ), .B(n2497), .Y(n239) );
  OAI21X1 U407 ( .A(n2453), .B(n2498), .C(n240), .Y(n1392) );
  NAND2X1 U408 ( .A(\mem<39><4> ), .B(n2497), .Y(n240) );
  OAI21X1 U409 ( .A(n2454), .B(n2498), .C(n241), .Y(n1393) );
  NAND2X1 U410 ( .A(\mem<39><5> ), .B(n2497), .Y(n241) );
  OAI21X1 U411 ( .A(n2455), .B(n2498), .C(n242), .Y(n1394) );
  NAND2X1 U412 ( .A(\mem<39><6> ), .B(n2497), .Y(n242) );
  OAI21X1 U413 ( .A(n2456), .B(n2498), .C(n243), .Y(n1395) );
  NAND2X1 U414 ( .A(\mem<39><7> ), .B(n2497), .Y(n243) );
  OAI21X1 U415 ( .A(n2457), .B(n2498), .C(n244), .Y(n1396) );
  NAND2X1 U416 ( .A(\mem<38><0> ), .B(n2497), .Y(n244) );
  OAI21X1 U417 ( .A(n2458), .B(n2498), .C(n245), .Y(n1397) );
  NAND2X1 U418 ( .A(\mem<38><1> ), .B(n2497), .Y(n245) );
  OAI21X1 U419 ( .A(n2459), .B(n2498), .C(n246), .Y(n1398) );
  NAND2X1 U420 ( .A(\mem<38><2> ), .B(n2497), .Y(n246) );
  OAI21X1 U421 ( .A(n2460), .B(n2498), .C(n247), .Y(n1399) );
  NAND2X1 U422 ( .A(\mem<38><3> ), .B(n2497), .Y(n247) );
  OAI21X1 U423 ( .A(n2461), .B(n2497), .C(n248), .Y(n1400) );
  NAND2X1 U424 ( .A(\mem<38><4> ), .B(n2497), .Y(n248) );
  OAI21X1 U425 ( .A(n2462), .B(n2497), .C(n249), .Y(n1401) );
  NAND2X1 U426 ( .A(\mem<38><5> ), .B(n2497), .Y(n249) );
  OAI21X1 U427 ( .A(n2463), .B(n2497), .C(n250), .Y(n1402) );
  NAND2X1 U428 ( .A(\mem<38><6> ), .B(n2498), .Y(n250) );
  OAI21X1 U429 ( .A(n2464), .B(n2497), .C(n251), .Y(n1403) );
  NAND2X1 U430 ( .A(\mem<38><7> ), .B(n2498), .Y(n251) );
  OAI21X1 U432 ( .A(n2449), .B(n2496), .C(n254), .Y(n1404) );
  NAND2X1 U433 ( .A(\mem<37><0> ), .B(n2496), .Y(n254) );
  OAI21X1 U434 ( .A(n2450), .B(n2496), .C(n255), .Y(n1405) );
  NAND2X1 U435 ( .A(\mem<37><1> ), .B(n2496), .Y(n255) );
  OAI21X1 U436 ( .A(n2451), .B(n2496), .C(n256), .Y(n1406) );
  NAND2X1 U437 ( .A(\mem<37><2> ), .B(n2495), .Y(n256) );
  OAI21X1 U438 ( .A(n2452), .B(n2496), .C(n257), .Y(n1407) );
  NAND2X1 U439 ( .A(\mem<37><3> ), .B(n2495), .Y(n257) );
  OAI21X1 U440 ( .A(n2453), .B(n2496), .C(n258), .Y(n1408) );
  NAND2X1 U441 ( .A(\mem<37><4> ), .B(n2495), .Y(n258) );
  OAI21X1 U442 ( .A(n2454), .B(n2496), .C(n259), .Y(n1409) );
  NAND2X1 U443 ( .A(\mem<37><5> ), .B(n2495), .Y(n259) );
  OAI21X1 U444 ( .A(n2455), .B(n2496), .C(n260), .Y(n1410) );
  NAND2X1 U445 ( .A(\mem<37><6> ), .B(n2495), .Y(n260) );
  OAI21X1 U446 ( .A(n2456), .B(n2496), .C(n261), .Y(n1411) );
  NAND2X1 U447 ( .A(\mem<37><7> ), .B(n2495), .Y(n261) );
  OAI21X1 U448 ( .A(n2457), .B(n2496), .C(n262), .Y(n1412) );
  NAND2X1 U449 ( .A(\mem<36><0> ), .B(n2495), .Y(n262) );
  OAI21X1 U450 ( .A(n2458), .B(n2496), .C(n263), .Y(n1413) );
  NAND2X1 U451 ( .A(\mem<36><1> ), .B(n2495), .Y(n263) );
  OAI21X1 U452 ( .A(n2459), .B(n2496), .C(n264), .Y(n1414) );
  NAND2X1 U453 ( .A(\mem<36><2> ), .B(n2495), .Y(n264) );
  OAI21X1 U454 ( .A(n2460), .B(n2496), .C(n265), .Y(n1415) );
  NAND2X1 U455 ( .A(\mem<36><3> ), .B(n2495), .Y(n265) );
  OAI21X1 U456 ( .A(n2461), .B(n2495), .C(n266), .Y(n1416) );
  NAND2X1 U457 ( .A(\mem<36><4> ), .B(n2495), .Y(n266) );
  OAI21X1 U458 ( .A(n2462), .B(n2495), .C(n267), .Y(n1417) );
  NAND2X1 U459 ( .A(\mem<36><5> ), .B(n2495), .Y(n267) );
  OAI21X1 U460 ( .A(n2463), .B(n2495), .C(n268), .Y(n1418) );
  NAND2X1 U461 ( .A(\mem<36><6> ), .B(n2496), .Y(n268) );
  OAI21X1 U462 ( .A(n2464), .B(n2495), .C(n269), .Y(n1419) );
  NAND2X1 U463 ( .A(\mem<36><7> ), .B(n2496), .Y(n269) );
  OAI21X1 U465 ( .A(n2449), .B(n2494), .C(n272), .Y(n1420) );
  NAND2X1 U466 ( .A(\mem<35><0> ), .B(n2494), .Y(n272) );
  OAI21X1 U467 ( .A(n2450), .B(n2494), .C(n273), .Y(n1421) );
  NAND2X1 U468 ( .A(\mem<35><1> ), .B(n2494), .Y(n273) );
  OAI21X1 U469 ( .A(n2451), .B(n2494), .C(n274), .Y(n1422) );
  NAND2X1 U470 ( .A(\mem<35><2> ), .B(n2493), .Y(n274) );
  OAI21X1 U471 ( .A(n2452), .B(n2494), .C(n275), .Y(n1423) );
  NAND2X1 U472 ( .A(\mem<35><3> ), .B(n2493), .Y(n275) );
  OAI21X1 U473 ( .A(n2453), .B(n2494), .C(n276), .Y(n1424) );
  NAND2X1 U474 ( .A(\mem<35><4> ), .B(n2493), .Y(n276) );
  OAI21X1 U475 ( .A(n2454), .B(n2494), .C(n277), .Y(n1425) );
  NAND2X1 U476 ( .A(\mem<35><5> ), .B(n2493), .Y(n277) );
  OAI21X1 U477 ( .A(n2455), .B(n2494), .C(n278), .Y(n1426) );
  NAND2X1 U478 ( .A(\mem<35><6> ), .B(n2493), .Y(n278) );
  OAI21X1 U479 ( .A(n2456), .B(n2494), .C(n279), .Y(n1427) );
  NAND2X1 U480 ( .A(\mem<35><7> ), .B(n2493), .Y(n279) );
  OAI21X1 U481 ( .A(n2457), .B(n2494), .C(n280), .Y(n1428) );
  NAND2X1 U482 ( .A(\mem<34><0> ), .B(n2493), .Y(n280) );
  OAI21X1 U483 ( .A(n2458), .B(n2494), .C(n281), .Y(n1429) );
  NAND2X1 U484 ( .A(\mem<34><1> ), .B(n2493), .Y(n281) );
  OAI21X1 U485 ( .A(n2459), .B(n2494), .C(n282), .Y(n1430) );
  NAND2X1 U486 ( .A(\mem<34><2> ), .B(n2493), .Y(n282) );
  OAI21X1 U487 ( .A(n2460), .B(n2494), .C(n283), .Y(n1431) );
  NAND2X1 U488 ( .A(\mem<34><3> ), .B(n2493), .Y(n283) );
  OAI21X1 U489 ( .A(n2461), .B(n2493), .C(n284), .Y(n1432) );
  NAND2X1 U490 ( .A(\mem<34><4> ), .B(n2493), .Y(n284) );
  OAI21X1 U491 ( .A(n2462), .B(n2493), .C(n285), .Y(n1433) );
  NAND2X1 U492 ( .A(\mem<34><5> ), .B(n2493), .Y(n285) );
  OAI21X1 U493 ( .A(n2463), .B(n2493), .C(n286), .Y(n1434) );
  NAND2X1 U494 ( .A(\mem<34><6> ), .B(n2494), .Y(n286) );
  OAI21X1 U495 ( .A(n2464), .B(n2493), .C(n287), .Y(n1435) );
  NAND2X1 U496 ( .A(\mem<34><7> ), .B(n2494), .Y(n287) );
  OAI21X1 U498 ( .A(n2449), .B(n2492), .C(n290), .Y(n1436) );
  NAND2X1 U499 ( .A(\mem<33><0> ), .B(n2492), .Y(n290) );
  OAI21X1 U500 ( .A(n2450), .B(n2492), .C(n291), .Y(n1437) );
  NAND2X1 U501 ( .A(\mem<33><1> ), .B(n2492), .Y(n291) );
  OAI21X1 U502 ( .A(n2451), .B(n2492), .C(n292), .Y(n1438) );
  NAND2X1 U503 ( .A(\mem<33><2> ), .B(n2491), .Y(n292) );
  OAI21X1 U504 ( .A(n2452), .B(n2492), .C(n293), .Y(n1439) );
  NAND2X1 U505 ( .A(\mem<33><3> ), .B(n2491), .Y(n293) );
  OAI21X1 U506 ( .A(n2453), .B(n2492), .C(n294), .Y(n1440) );
  NAND2X1 U507 ( .A(\mem<33><4> ), .B(n2491), .Y(n294) );
  OAI21X1 U508 ( .A(n2454), .B(n2492), .C(n295), .Y(n1441) );
  NAND2X1 U509 ( .A(\mem<33><5> ), .B(n2491), .Y(n295) );
  OAI21X1 U510 ( .A(n2455), .B(n2492), .C(n296), .Y(n1442) );
  NAND2X1 U511 ( .A(\mem<33><6> ), .B(n2491), .Y(n296) );
  OAI21X1 U512 ( .A(n2456), .B(n2492), .C(n297), .Y(n1443) );
  NAND2X1 U513 ( .A(\mem<33><7> ), .B(n2491), .Y(n297) );
  OAI21X1 U514 ( .A(n2457), .B(n2492), .C(n298), .Y(n1444) );
  NAND2X1 U515 ( .A(\mem<32><0> ), .B(n2491), .Y(n298) );
  OAI21X1 U516 ( .A(n2458), .B(n2492), .C(n299), .Y(n1445) );
  NAND2X1 U517 ( .A(\mem<32><1> ), .B(n2491), .Y(n299) );
  OAI21X1 U518 ( .A(n2459), .B(n2492), .C(n300), .Y(n1446) );
  NAND2X1 U519 ( .A(\mem<32><2> ), .B(n2491), .Y(n300) );
  OAI21X1 U520 ( .A(n2460), .B(n2492), .C(n301), .Y(n1447) );
  NAND2X1 U521 ( .A(\mem<32><3> ), .B(n2491), .Y(n301) );
  OAI21X1 U522 ( .A(n2461), .B(n2491), .C(n302), .Y(n1448) );
  NAND2X1 U523 ( .A(\mem<32><4> ), .B(n2491), .Y(n302) );
  OAI21X1 U524 ( .A(n2462), .B(n2491), .C(n303), .Y(n1449) );
  NAND2X1 U525 ( .A(\mem<32><5> ), .B(n2491), .Y(n303) );
  OAI21X1 U526 ( .A(n2463), .B(n2491), .C(n304), .Y(n1450) );
  NAND2X1 U527 ( .A(\mem<32><6> ), .B(n2492), .Y(n304) );
  OAI21X1 U528 ( .A(n2464), .B(n2491), .C(n305), .Y(n1451) );
  NAND2X1 U529 ( .A(\mem<32><7> ), .B(n2492), .Y(n305) );
  OAI21X1 U531 ( .A(n2449), .B(n2490), .C(n308), .Y(n1452) );
  NAND2X1 U532 ( .A(\mem<31><0> ), .B(n2490), .Y(n308) );
  OAI21X1 U533 ( .A(n2450), .B(n2490), .C(n309), .Y(n1453) );
  NAND2X1 U534 ( .A(\mem<31><1> ), .B(n2490), .Y(n309) );
  OAI21X1 U535 ( .A(n2451), .B(n2490), .C(n310), .Y(n1454) );
  NAND2X1 U536 ( .A(\mem<31><2> ), .B(n2489), .Y(n310) );
  OAI21X1 U537 ( .A(n2452), .B(n2490), .C(n311), .Y(n1455) );
  NAND2X1 U538 ( .A(\mem<31><3> ), .B(n2489), .Y(n311) );
  OAI21X1 U539 ( .A(n2453), .B(n2490), .C(n312), .Y(n1456) );
  NAND2X1 U540 ( .A(\mem<31><4> ), .B(n2489), .Y(n312) );
  OAI21X1 U541 ( .A(n2454), .B(n2490), .C(n313), .Y(n1457) );
  NAND2X1 U542 ( .A(\mem<31><5> ), .B(n2489), .Y(n313) );
  OAI21X1 U543 ( .A(n2455), .B(n2490), .C(n314), .Y(n1458) );
  NAND2X1 U544 ( .A(\mem<31><6> ), .B(n2489), .Y(n314) );
  OAI21X1 U545 ( .A(n2456), .B(n2490), .C(n315), .Y(n1459) );
  NAND2X1 U546 ( .A(\mem<31><7> ), .B(n2489), .Y(n315) );
  OAI21X1 U547 ( .A(n2457), .B(n2490), .C(n316), .Y(n1460) );
  NAND2X1 U548 ( .A(\mem<30><0> ), .B(n2489), .Y(n316) );
  OAI21X1 U549 ( .A(n2458), .B(n2490), .C(n317), .Y(n1461) );
  NAND2X1 U550 ( .A(\mem<30><1> ), .B(n2489), .Y(n317) );
  OAI21X1 U551 ( .A(n2459), .B(n2490), .C(n318), .Y(n1462) );
  NAND2X1 U552 ( .A(\mem<30><2> ), .B(n2489), .Y(n318) );
  OAI21X1 U553 ( .A(n2460), .B(n2490), .C(n319), .Y(n1463) );
  NAND2X1 U554 ( .A(\mem<30><3> ), .B(n2489), .Y(n319) );
  OAI21X1 U555 ( .A(n2461), .B(n2489), .C(n320), .Y(n1464) );
  NAND2X1 U556 ( .A(\mem<30><4> ), .B(n2489), .Y(n320) );
  OAI21X1 U557 ( .A(n2462), .B(n2489), .C(n321), .Y(n1465) );
  NAND2X1 U558 ( .A(\mem<30><5> ), .B(n2489), .Y(n321) );
  OAI21X1 U559 ( .A(n2463), .B(n2489), .C(n322), .Y(n1466) );
  NAND2X1 U560 ( .A(\mem<30><6> ), .B(n2490), .Y(n322) );
  OAI21X1 U561 ( .A(n2464), .B(n2489), .C(n323), .Y(n1467) );
  NAND2X1 U562 ( .A(\mem<30><7> ), .B(n2490), .Y(n323) );
  OAI21X1 U564 ( .A(n2449), .B(n2488), .C(n326), .Y(n1468) );
  NAND2X1 U565 ( .A(\mem<29><0> ), .B(n2488), .Y(n326) );
  OAI21X1 U566 ( .A(n2450), .B(n2488), .C(n327), .Y(n1469) );
  NAND2X1 U567 ( .A(\mem<29><1> ), .B(n2488), .Y(n327) );
  OAI21X1 U568 ( .A(n2451), .B(n2488), .C(n328), .Y(n1470) );
  NAND2X1 U569 ( .A(\mem<29><2> ), .B(n2487), .Y(n328) );
  OAI21X1 U570 ( .A(n2452), .B(n2488), .C(n329), .Y(n1471) );
  NAND2X1 U571 ( .A(\mem<29><3> ), .B(n2487), .Y(n329) );
  OAI21X1 U572 ( .A(n2453), .B(n2488), .C(n330), .Y(n1472) );
  NAND2X1 U573 ( .A(\mem<29><4> ), .B(n2487), .Y(n330) );
  OAI21X1 U574 ( .A(n2454), .B(n2488), .C(n331), .Y(n1473) );
  NAND2X1 U575 ( .A(\mem<29><5> ), .B(n2487), .Y(n331) );
  OAI21X1 U576 ( .A(n2455), .B(n2488), .C(n332), .Y(n1474) );
  NAND2X1 U577 ( .A(\mem<29><6> ), .B(n2487), .Y(n332) );
  OAI21X1 U578 ( .A(n2456), .B(n2488), .C(n333), .Y(n1475) );
  NAND2X1 U579 ( .A(\mem<29><7> ), .B(n2487), .Y(n333) );
  OAI21X1 U580 ( .A(n2457), .B(n2488), .C(n334), .Y(n1476) );
  NAND2X1 U581 ( .A(\mem<28><0> ), .B(n2487), .Y(n334) );
  OAI21X1 U582 ( .A(n2458), .B(n2488), .C(n335), .Y(n1477) );
  NAND2X1 U583 ( .A(\mem<28><1> ), .B(n2487), .Y(n335) );
  OAI21X1 U584 ( .A(n2459), .B(n2488), .C(n336), .Y(n1478) );
  NAND2X1 U585 ( .A(\mem<28><2> ), .B(n2487), .Y(n336) );
  OAI21X1 U586 ( .A(n2460), .B(n2488), .C(n337), .Y(n1479) );
  NAND2X1 U587 ( .A(\mem<28><3> ), .B(n2487), .Y(n337) );
  OAI21X1 U588 ( .A(n2461), .B(n2487), .C(n338), .Y(n1480) );
  NAND2X1 U589 ( .A(\mem<28><4> ), .B(n2487), .Y(n338) );
  OAI21X1 U590 ( .A(n2462), .B(n2487), .C(n339), .Y(n1481) );
  NAND2X1 U591 ( .A(\mem<28><5> ), .B(n2487), .Y(n339) );
  OAI21X1 U592 ( .A(n2463), .B(n2487), .C(n340), .Y(n1482) );
  NAND2X1 U593 ( .A(\mem<28><6> ), .B(n2488), .Y(n340) );
  OAI21X1 U594 ( .A(n2464), .B(n2487), .C(n341), .Y(n1483) );
  NAND2X1 U595 ( .A(\mem<28><7> ), .B(n2488), .Y(n341) );
  OAI21X1 U597 ( .A(n2449), .B(n2486), .C(n344), .Y(n1484) );
  NAND2X1 U598 ( .A(\mem<27><0> ), .B(n2486), .Y(n344) );
  OAI21X1 U599 ( .A(n2450), .B(n2486), .C(n345), .Y(n1485) );
  NAND2X1 U600 ( .A(\mem<27><1> ), .B(n2486), .Y(n345) );
  OAI21X1 U601 ( .A(n2451), .B(n2486), .C(n346), .Y(n1486) );
  NAND2X1 U602 ( .A(\mem<27><2> ), .B(n2485), .Y(n346) );
  OAI21X1 U603 ( .A(n2452), .B(n2486), .C(n347), .Y(n1487) );
  NAND2X1 U604 ( .A(\mem<27><3> ), .B(n2485), .Y(n347) );
  OAI21X1 U605 ( .A(n2453), .B(n2486), .C(n348), .Y(n1488) );
  NAND2X1 U606 ( .A(\mem<27><4> ), .B(n2485), .Y(n348) );
  OAI21X1 U607 ( .A(n2454), .B(n2486), .C(n349), .Y(n1489) );
  NAND2X1 U608 ( .A(\mem<27><5> ), .B(n2485), .Y(n349) );
  OAI21X1 U609 ( .A(n2455), .B(n2486), .C(n350), .Y(n1490) );
  NAND2X1 U610 ( .A(\mem<27><6> ), .B(n2485), .Y(n350) );
  OAI21X1 U611 ( .A(n2456), .B(n2486), .C(n351), .Y(n1491) );
  NAND2X1 U612 ( .A(\mem<27><7> ), .B(n2485), .Y(n351) );
  OAI21X1 U613 ( .A(n2457), .B(n2486), .C(n352), .Y(n1492) );
  NAND2X1 U614 ( .A(\mem<26><0> ), .B(n2485), .Y(n352) );
  OAI21X1 U615 ( .A(n2458), .B(n2486), .C(n353), .Y(n1493) );
  NAND2X1 U616 ( .A(\mem<26><1> ), .B(n2485), .Y(n353) );
  OAI21X1 U617 ( .A(n2459), .B(n2486), .C(n354), .Y(n1494) );
  NAND2X1 U618 ( .A(\mem<26><2> ), .B(n2485), .Y(n354) );
  OAI21X1 U619 ( .A(n2460), .B(n2486), .C(n355), .Y(n1495) );
  NAND2X1 U620 ( .A(\mem<26><3> ), .B(n2485), .Y(n355) );
  OAI21X1 U621 ( .A(n2461), .B(n2485), .C(n356), .Y(n1496) );
  NAND2X1 U622 ( .A(\mem<26><4> ), .B(n2485), .Y(n356) );
  OAI21X1 U623 ( .A(n2462), .B(n2485), .C(n357), .Y(n1497) );
  NAND2X1 U624 ( .A(\mem<26><5> ), .B(n2485), .Y(n357) );
  OAI21X1 U625 ( .A(n2463), .B(n2485), .C(n358), .Y(n1498) );
  NAND2X1 U626 ( .A(\mem<26><6> ), .B(n2486), .Y(n358) );
  OAI21X1 U627 ( .A(n2464), .B(n2485), .C(n359), .Y(n1499) );
  NAND2X1 U628 ( .A(\mem<26><7> ), .B(n2486), .Y(n359) );
  OAI21X1 U630 ( .A(n2449), .B(n2484), .C(n362), .Y(n1500) );
  NAND2X1 U631 ( .A(\mem<25><0> ), .B(n2484), .Y(n362) );
  OAI21X1 U632 ( .A(n2450), .B(n2484), .C(n363), .Y(n1501) );
  NAND2X1 U633 ( .A(\mem<25><1> ), .B(n2484), .Y(n363) );
  OAI21X1 U634 ( .A(n2451), .B(n2484), .C(n364), .Y(n1502) );
  NAND2X1 U635 ( .A(\mem<25><2> ), .B(n2483), .Y(n364) );
  OAI21X1 U636 ( .A(n2452), .B(n2484), .C(n365), .Y(n1503) );
  NAND2X1 U637 ( .A(\mem<25><3> ), .B(n2483), .Y(n365) );
  OAI21X1 U638 ( .A(n2453), .B(n2484), .C(n366), .Y(n1504) );
  NAND2X1 U639 ( .A(\mem<25><4> ), .B(n2483), .Y(n366) );
  OAI21X1 U640 ( .A(n2454), .B(n2484), .C(n367), .Y(n1505) );
  NAND2X1 U641 ( .A(\mem<25><5> ), .B(n2483), .Y(n367) );
  OAI21X1 U642 ( .A(n2455), .B(n2484), .C(n368), .Y(n1506) );
  NAND2X1 U643 ( .A(\mem<25><6> ), .B(n2483), .Y(n368) );
  OAI21X1 U644 ( .A(n2456), .B(n2484), .C(n369), .Y(n1507) );
  NAND2X1 U645 ( .A(\mem<25><7> ), .B(n2483), .Y(n369) );
  OAI21X1 U646 ( .A(n2457), .B(n2484), .C(n370), .Y(n1508) );
  NAND2X1 U647 ( .A(\mem<24><0> ), .B(n2483), .Y(n370) );
  OAI21X1 U648 ( .A(n2458), .B(n2484), .C(n371), .Y(n1509) );
  NAND2X1 U649 ( .A(\mem<24><1> ), .B(n2483), .Y(n371) );
  OAI21X1 U650 ( .A(n2459), .B(n2484), .C(n372), .Y(n1510) );
  NAND2X1 U651 ( .A(\mem<24><2> ), .B(n2483), .Y(n372) );
  OAI21X1 U652 ( .A(n2460), .B(n2484), .C(n373), .Y(n1511) );
  NAND2X1 U653 ( .A(\mem<24><3> ), .B(n2483), .Y(n373) );
  OAI21X1 U654 ( .A(n2461), .B(n2483), .C(n374), .Y(n1512) );
  NAND2X1 U655 ( .A(\mem<24><4> ), .B(n2483), .Y(n374) );
  OAI21X1 U656 ( .A(n2462), .B(n2483), .C(n375), .Y(n1513) );
  NAND2X1 U657 ( .A(\mem<24><5> ), .B(n2483), .Y(n375) );
  OAI21X1 U658 ( .A(n2463), .B(n2483), .C(n376), .Y(n1514) );
  NAND2X1 U659 ( .A(\mem<24><6> ), .B(n2484), .Y(n376) );
  OAI21X1 U660 ( .A(n2464), .B(n2483), .C(n377), .Y(n1515) );
  NAND2X1 U661 ( .A(\mem<24><7> ), .B(n2484), .Y(n377) );
  OAI21X1 U663 ( .A(n2449), .B(n2482), .C(n380), .Y(n1516) );
  NAND2X1 U664 ( .A(\mem<23><0> ), .B(n2482), .Y(n380) );
  OAI21X1 U665 ( .A(n2450), .B(n2482), .C(n381), .Y(n1517) );
  NAND2X1 U666 ( .A(\mem<23><1> ), .B(n2482), .Y(n381) );
  OAI21X1 U667 ( .A(n2451), .B(n2482), .C(n382), .Y(n1518) );
  NAND2X1 U668 ( .A(\mem<23><2> ), .B(n2481), .Y(n382) );
  OAI21X1 U669 ( .A(n2452), .B(n2482), .C(n383), .Y(n1519) );
  NAND2X1 U670 ( .A(\mem<23><3> ), .B(n2481), .Y(n383) );
  OAI21X1 U671 ( .A(n2453), .B(n2482), .C(n384), .Y(n1520) );
  NAND2X1 U672 ( .A(\mem<23><4> ), .B(n2481), .Y(n384) );
  OAI21X1 U673 ( .A(n2454), .B(n2482), .C(n385), .Y(n1521) );
  NAND2X1 U674 ( .A(\mem<23><5> ), .B(n2481), .Y(n385) );
  OAI21X1 U675 ( .A(n2455), .B(n2482), .C(n386), .Y(n1522) );
  NAND2X1 U676 ( .A(\mem<23><6> ), .B(n2481), .Y(n386) );
  OAI21X1 U677 ( .A(n2456), .B(n2482), .C(n387), .Y(n1523) );
  NAND2X1 U678 ( .A(\mem<23><7> ), .B(n2481), .Y(n387) );
  OAI21X1 U679 ( .A(n2457), .B(n2482), .C(n388), .Y(n1524) );
  NAND2X1 U680 ( .A(\mem<22><0> ), .B(n2481), .Y(n388) );
  OAI21X1 U681 ( .A(n2458), .B(n2482), .C(n389), .Y(n1525) );
  NAND2X1 U682 ( .A(\mem<22><1> ), .B(n2481), .Y(n389) );
  OAI21X1 U683 ( .A(n2459), .B(n2482), .C(n390), .Y(n1526) );
  NAND2X1 U684 ( .A(\mem<22><2> ), .B(n2481), .Y(n390) );
  OAI21X1 U685 ( .A(n2460), .B(n2482), .C(n391), .Y(n1527) );
  NAND2X1 U686 ( .A(\mem<22><3> ), .B(n2481), .Y(n391) );
  OAI21X1 U687 ( .A(n2461), .B(n2481), .C(n392), .Y(n1528) );
  NAND2X1 U688 ( .A(\mem<22><4> ), .B(n2481), .Y(n392) );
  OAI21X1 U689 ( .A(n2462), .B(n2481), .C(n393), .Y(n1529) );
  NAND2X1 U690 ( .A(\mem<22><5> ), .B(n2481), .Y(n393) );
  OAI21X1 U691 ( .A(n2463), .B(n2481), .C(n394), .Y(n1530) );
  NAND2X1 U692 ( .A(\mem<22><6> ), .B(n2482), .Y(n394) );
  OAI21X1 U693 ( .A(n2464), .B(n2481), .C(n395), .Y(n1531) );
  NAND2X1 U694 ( .A(\mem<22><7> ), .B(n2482), .Y(n395) );
  OAI21X1 U696 ( .A(n2449), .B(n2480), .C(n398), .Y(n1532) );
  NAND2X1 U697 ( .A(\mem<21><0> ), .B(n2480), .Y(n398) );
  OAI21X1 U698 ( .A(n2450), .B(n2480), .C(n399), .Y(n1533) );
  NAND2X1 U699 ( .A(\mem<21><1> ), .B(n2480), .Y(n399) );
  OAI21X1 U700 ( .A(n2451), .B(n2480), .C(n400), .Y(n1534) );
  NAND2X1 U701 ( .A(\mem<21><2> ), .B(n2479), .Y(n400) );
  OAI21X1 U702 ( .A(n2452), .B(n2480), .C(n401), .Y(n1535) );
  NAND2X1 U703 ( .A(\mem<21><3> ), .B(n2479), .Y(n401) );
  OAI21X1 U704 ( .A(n2453), .B(n2480), .C(n402), .Y(n1536) );
  NAND2X1 U705 ( .A(\mem<21><4> ), .B(n2479), .Y(n402) );
  OAI21X1 U706 ( .A(n2454), .B(n2480), .C(n403), .Y(n1537) );
  NAND2X1 U707 ( .A(\mem<21><5> ), .B(n2479), .Y(n403) );
  OAI21X1 U708 ( .A(n2455), .B(n2480), .C(n404), .Y(n1538) );
  NAND2X1 U709 ( .A(\mem<21><6> ), .B(n2479), .Y(n404) );
  OAI21X1 U710 ( .A(n2456), .B(n2480), .C(n405), .Y(n1539) );
  NAND2X1 U711 ( .A(\mem<21><7> ), .B(n2479), .Y(n405) );
  OAI21X1 U712 ( .A(n2457), .B(n2480), .C(n406), .Y(n1540) );
  NAND2X1 U713 ( .A(\mem<20><0> ), .B(n2479), .Y(n406) );
  OAI21X1 U714 ( .A(n2458), .B(n2480), .C(n407), .Y(n1541) );
  NAND2X1 U715 ( .A(\mem<20><1> ), .B(n2479), .Y(n407) );
  OAI21X1 U716 ( .A(n2459), .B(n2480), .C(n408), .Y(n1542) );
  NAND2X1 U717 ( .A(\mem<20><2> ), .B(n2479), .Y(n408) );
  OAI21X1 U718 ( .A(n2460), .B(n2480), .C(n409), .Y(n1543) );
  NAND2X1 U719 ( .A(\mem<20><3> ), .B(n2479), .Y(n409) );
  OAI21X1 U720 ( .A(n2461), .B(n2479), .C(n410), .Y(n1544) );
  NAND2X1 U721 ( .A(\mem<20><4> ), .B(n2479), .Y(n410) );
  OAI21X1 U722 ( .A(n2462), .B(n2479), .C(n411), .Y(n1545) );
  NAND2X1 U723 ( .A(\mem<20><5> ), .B(n2479), .Y(n411) );
  OAI21X1 U724 ( .A(n2463), .B(n2479), .C(n412), .Y(n1546) );
  NAND2X1 U725 ( .A(\mem<20><6> ), .B(n2480), .Y(n412) );
  OAI21X1 U726 ( .A(n2464), .B(n2479), .C(n413), .Y(n1547) );
  NAND2X1 U727 ( .A(\mem<20><7> ), .B(n2480), .Y(n413) );
  OAI21X1 U729 ( .A(n2449), .B(n2478), .C(n416), .Y(n1548) );
  NAND2X1 U730 ( .A(\mem<19><0> ), .B(n2478), .Y(n416) );
  OAI21X1 U731 ( .A(n2450), .B(n2478), .C(n417), .Y(n1549) );
  NAND2X1 U732 ( .A(\mem<19><1> ), .B(n2478), .Y(n417) );
  OAI21X1 U733 ( .A(n2451), .B(n2478), .C(n418), .Y(n1550) );
  NAND2X1 U734 ( .A(\mem<19><2> ), .B(n2477), .Y(n418) );
  OAI21X1 U735 ( .A(n2452), .B(n2478), .C(n419), .Y(n1551) );
  NAND2X1 U736 ( .A(\mem<19><3> ), .B(n2477), .Y(n419) );
  OAI21X1 U737 ( .A(n2453), .B(n2478), .C(n420), .Y(n1552) );
  NAND2X1 U738 ( .A(\mem<19><4> ), .B(n2477), .Y(n420) );
  OAI21X1 U739 ( .A(n2454), .B(n2478), .C(n421), .Y(n1553) );
  NAND2X1 U740 ( .A(\mem<19><5> ), .B(n2477), .Y(n421) );
  OAI21X1 U741 ( .A(n2455), .B(n2478), .C(n422), .Y(n1554) );
  NAND2X1 U742 ( .A(\mem<19><6> ), .B(n2477), .Y(n422) );
  OAI21X1 U743 ( .A(n2456), .B(n2478), .C(n423), .Y(n1555) );
  NAND2X1 U744 ( .A(\mem<19><7> ), .B(n2477), .Y(n423) );
  OAI21X1 U745 ( .A(n2457), .B(n2478), .C(n424), .Y(n1556) );
  NAND2X1 U746 ( .A(\mem<18><0> ), .B(n2477), .Y(n424) );
  OAI21X1 U747 ( .A(n2458), .B(n2478), .C(n425), .Y(n1557) );
  NAND2X1 U748 ( .A(\mem<18><1> ), .B(n2477), .Y(n425) );
  OAI21X1 U749 ( .A(n2459), .B(n2478), .C(n426), .Y(n1558) );
  NAND2X1 U750 ( .A(\mem<18><2> ), .B(n2477), .Y(n426) );
  OAI21X1 U751 ( .A(n2460), .B(n2478), .C(n427), .Y(n1559) );
  NAND2X1 U752 ( .A(\mem<18><3> ), .B(n2477), .Y(n427) );
  OAI21X1 U753 ( .A(n2461), .B(n2477), .C(n428), .Y(n1560) );
  NAND2X1 U754 ( .A(\mem<18><4> ), .B(n2477), .Y(n428) );
  OAI21X1 U755 ( .A(n2462), .B(n2477), .C(n429), .Y(n1561) );
  NAND2X1 U756 ( .A(\mem<18><5> ), .B(n2477), .Y(n429) );
  OAI21X1 U757 ( .A(n2463), .B(n2477), .C(n430), .Y(n1562) );
  NAND2X1 U758 ( .A(\mem<18><6> ), .B(n2478), .Y(n430) );
  OAI21X1 U759 ( .A(n2464), .B(n2477), .C(n431), .Y(n1563) );
  NAND2X1 U760 ( .A(\mem<18><7> ), .B(n2478), .Y(n431) );
  OAI21X1 U762 ( .A(n2449), .B(n2476), .C(n434), .Y(n1564) );
  NAND2X1 U763 ( .A(\mem<17><0> ), .B(n2476), .Y(n434) );
  OAI21X1 U764 ( .A(n2450), .B(n2476), .C(n435), .Y(n1565) );
  NAND2X1 U765 ( .A(\mem<17><1> ), .B(n2476), .Y(n435) );
  OAI21X1 U766 ( .A(n2451), .B(n2476), .C(n436), .Y(n1566) );
  NAND2X1 U767 ( .A(\mem<17><2> ), .B(n2475), .Y(n436) );
  OAI21X1 U768 ( .A(n2452), .B(n2476), .C(n437), .Y(n1567) );
  NAND2X1 U769 ( .A(\mem<17><3> ), .B(n2475), .Y(n437) );
  OAI21X1 U770 ( .A(n2453), .B(n2476), .C(n438), .Y(n1568) );
  NAND2X1 U771 ( .A(\mem<17><4> ), .B(n2475), .Y(n438) );
  OAI21X1 U772 ( .A(n2454), .B(n2476), .C(n439), .Y(n1569) );
  NAND2X1 U773 ( .A(\mem<17><5> ), .B(n2475), .Y(n439) );
  OAI21X1 U774 ( .A(n2455), .B(n2476), .C(n440), .Y(n1570) );
  NAND2X1 U775 ( .A(\mem<17><6> ), .B(n2475), .Y(n440) );
  OAI21X1 U776 ( .A(n2456), .B(n2476), .C(n441), .Y(n1571) );
  NAND2X1 U777 ( .A(\mem<17><7> ), .B(n2475), .Y(n441) );
  OAI21X1 U778 ( .A(n2457), .B(n2476), .C(n442), .Y(n1572) );
  NAND2X1 U779 ( .A(\mem<16><0> ), .B(n2475), .Y(n442) );
  OAI21X1 U780 ( .A(n2458), .B(n2476), .C(n443), .Y(n1573) );
  NAND2X1 U781 ( .A(\mem<16><1> ), .B(n2475), .Y(n443) );
  OAI21X1 U782 ( .A(n2459), .B(n2476), .C(n444), .Y(n1574) );
  NAND2X1 U783 ( .A(\mem<16><2> ), .B(n2475), .Y(n444) );
  OAI21X1 U784 ( .A(n2460), .B(n2476), .C(n445), .Y(n1575) );
  NAND2X1 U785 ( .A(\mem<16><3> ), .B(n2475), .Y(n445) );
  OAI21X1 U786 ( .A(n2461), .B(n2475), .C(n446), .Y(n1576) );
  NAND2X1 U787 ( .A(\mem<16><4> ), .B(n2475), .Y(n446) );
  OAI21X1 U788 ( .A(n2462), .B(n2475), .C(n447), .Y(n1577) );
  NAND2X1 U789 ( .A(\mem<16><5> ), .B(n2475), .Y(n447) );
  OAI21X1 U790 ( .A(n2463), .B(n2475), .C(n448), .Y(n1578) );
  NAND2X1 U791 ( .A(\mem<16><6> ), .B(n2476), .Y(n448) );
  OAI21X1 U792 ( .A(n2464), .B(n2475), .C(n449), .Y(n1579) );
  NAND2X1 U793 ( .A(\mem<16><7> ), .B(n2476), .Y(n449) );
  OAI21X1 U795 ( .A(n2449), .B(n2474), .C(n452), .Y(n1580) );
  NAND2X1 U796 ( .A(\mem<15><0> ), .B(n2474), .Y(n452) );
  OAI21X1 U797 ( .A(n2450), .B(n2474), .C(n453), .Y(n1581) );
  NAND2X1 U798 ( .A(\mem<15><1> ), .B(n2474), .Y(n453) );
  OAI21X1 U799 ( .A(n2451), .B(n2474), .C(n454), .Y(n1582) );
  NAND2X1 U800 ( .A(\mem<15><2> ), .B(n2473), .Y(n454) );
  OAI21X1 U801 ( .A(n2452), .B(n2474), .C(n455), .Y(n1583) );
  NAND2X1 U802 ( .A(\mem<15><3> ), .B(n2473), .Y(n455) );
  OAI21X1 U803 ( .A(n2453), .B(n2474), .C(n456), .Y(n1584) );
  NAND2X1 U804 ( .A(\mem<15><4> ), .B(n2473), .Y(n456) );
  OAI21X1 U805 ( .A(n2454), .B(n2474), .C(n457), .Y(n1585) );
  NAND2X1 U806 ( .A(\mem<15><5> ), .B(n2473), .Y(n457) );
  OAI21X1 U807 ( .A(n2455), .B(n2474), .C(n458), .Y(n1586) );
  NAND2X1 U808 ( .A(\mem<15><6> ), .B(n2473), .Y(n458) );
  OAI21X1 U809 ( .A(n2456), .B(n2474), .C(n459), .Y(n1587) );
  NAND2X1 U810 ( .A(\mem<15><7> ), .B(n2473), .Y(n459) );
  OAI21X1 U811 ( .A(n2457), .B(n2474), .C(n460), .Y(n1588) );
  NAND2X1 U812 ( .A(\mem<14><0> ), .B(n2473), .Y(n460) );
  OAI21X1 U813 ( .A(n2458), .B(n2474), .C(n461), .Y(n1589) );
  NAND2X1 U814 ( .A(\mem<14><1> ), .B(n2473), .Y(n461) );
  OAI21X1 U815 ( .A(n2459), .B(n2474), .C(n462), .Y(n1590) );
  NAND2X1 U816 ( .A(\mem<14><2> ), .B(n2473), .Y(n462) );
  OAI21X1 U817 ( .A(n2460), .B(n2474), .C(n463), .Y(n1591) );
  NAND2X1 U818 ( .A(\mem<14><3> ), .B(n2473), .Y(n463) );
  OAI21X1 U819 ( .A(n2461), .B(n2473), .C(n464), .Y(n1592) );
  NAND2X1 U820 ( .A(\mem<14><4> ), .B(n2473), .Y(n464) );
  OAI21X1 U821 ( .A(n2462), .B(n2473), .C(n465), .Y(n1593) );
  NAND2X1 U822 ( .A(\mem<14><5> ), .B(n2473), .Y(n465) );
  OAI21X1 U823 ( .A(n2463), .B(n2473), .C(n466), .Y(n1594) );
  NAND2X1 U824 ( .A(\mem<14><6> ), .B(n2474), .Y(n466) );
  OAI21X1 U825 ( .A(n2464), .B(n2473), .C(n467), .Y(n1595) );
  NAND2X1 U826 ( .A(\mem<14><7> ), .B(n2474), .Y(n467) );
  OAI21X1 U828 ( .A(n2449), .B(n2472), .C(n470), .Y(n1596) );
  NAND2X1 U829 ( .A(\mem<13><0> ), .B(n2472), .Y(n470) );
  OAI21X1 U830 ( .A(n2450), .B(n2472), .C(n471), .Y(n1597) );
  NAND2X1 U831 ( .A(\mem<13><1> ), .B(n2472), .Y(n471) );
  OAI21X1 U832 ( .A(n2451), .B(n2472), .C(n472), .Y(n1598) );
  NAND2X1 U833 ( .A(\mem<13><2> ), .B(n2471), .Y(n472) );
  OAI21X1 U834 ( .A(n2452), .B(n2472), .C(n473), .Y(n1599) );
  NAND2X1 U835 ( .A(\mem<13><3> ), .B(n2471), .Y(n473) );
  OAI21X1 U836 ( .A(n2453), .B(n2472), .C(n474), .Y(n1600) );
  NAND2X1 U837 ( .A(\mem<13><4> ), .B(n2471), .Y(n474) );
  OAI21X1 U838 ( .A(n2454), .B(n2472), .C(n475), .Y(n1601) );
  NAND2X1 U839 ( .A(\mem<13><5> ), .B(n2471), .Y(n475) );
  OAI21X1 U840 ( .A(n2455), .B(n2472), .C(n476), .Y(n1602) );
  NAND2X1 U841 ( .A(\mem<13><6> ), .B(n2471), .Y(n476) );
  OAI21X1 U842 ( .A(n2456), .B(n2472), .C(n477), .Y(n1603) );
  NAND2X1 U843 ( .A(\mem<13><7> ), .B(n2471), .Y(n477) );
  OAI21X1 U844 ( .A(n2457), .B(n2472), .C(n478), .Y(n1604) );
  NAND2X1 U845 ( .A(\mem<12><0> ), .B(n2471), .Y(n478) );
  OAI21X1 U846 ( .A(n2458), .B(n2472), .C(n479), .Y(n1605) );
  NAND2X1 U847 ( .A(\mem<12><1> ), .B(n2471), .Y(n479) );
  OAI21X1 U848 ( .A(n2459), .B(n2472), .C(n480), .Y(n1606) );
  NAND2X1 U849 ( .A(\mem<12><2> ), .B(n2471), .Y(n480) );
  OAI21X1 U850 ( .A(n2460), .B(n2472), .C(n481), .Y(n1607) );
  NAND2X1 U851 ( .A(\mem<12><3> ), .B(n2471), .Y(n481) );
  OAI21X1 U852 ( .A(n2461), .B(n2471), .C(n482), .Y(n1608) );
  NAND2X1 U853 ( .A(\mem<12><4> ), .B(n2471), .Y(n482) );
  OAI21X1 U854 ( .A(n2462), .B(n2471), .C(n483), .Y(n1609) );
  NAND2X1 U855 ( .A(\mem<12><5> ), .B(n2471), .Y(n483) );
  OAI21X1 U856 ( .A(n2463), .B(n2471), .C(n484), .Y(n1610) );
  NAND2X1 U857 ( .A(\mem<12><6> ), .B(n2472), .Y(n484) );
  OAI21X1 U858 ( .A(n2464), .B(n2471), .C(n485), .Y(n1611) );
  NAND2X1 U859 ( .A(\mem<12><7> ), .B(n2472), .Y(n485) );
  OAI21X1 U861 ( .A(n2449), .B(n2470), .C(n488), .Y(n1612) );
  NAND2X1 U862 ( .A(\mem<11><0> ), .B(n2470), .Y(n488) );
  OAI21X1 U863 ( .A(n2450), .B(n2470), .C(n489), .Y(n1613) );
  NAND2X1 U864 ( .A(\mem<11><1> ), .B(n2470), .Y(n489) );
  OAI21X1 U865 ( .A(n2451), .B(n2470), .C(n490), .Y(n1614) );
  NAND2X1 U866 ( .A(\mem<11><2> ), .B(n2470), .Y(n490) );
  OAI21X1 U867 ( .A(n2452), .B(n2470), .C(n491), .Y(n1615) );
  NAND2X1 U868 ( .A(\mem<11><3> ), .B(n2470), .Y(n491) );
  OAI21X1 U869 ( .A(n2453), .B(n2470), .C(n492), .Y(n1616) );
  NAND2X1 U870 ( .A(\mem<11><4> ), .B(n2470), .Y(n492) );
  OAI21X1 U871 ( .A(n2454), .B(n2470), .C(n493), .Y(n1617) );
  NAND2X1 U872 ( .A(\mem<11><5> ), .B(n2470), .Y(n493) );
  OAI21X1 U873 ( .A(n2455), .B(n2470), .C(n494), .Y(n1618) );
  NAND2X1 U874 ( .A(\mem<11><6> ), .B(n2470), .Y(n494) );
  OAI21X1 U875 ( .A(n2456), .B(n2470), .C(n495), .Y(n1619) );
  NAND2X1 U876 ( .A(\mem<11><7> ), .B(n2470), .Y(n495) );
  OAI21X1 U877 ( .A(n2457), .B(n2470), .C(n496), .Y(n1620) );
  NAND2X1 U878 ( .A(\mem<10><0> ), .B(n2470), .Y(n496) );
  OAI21X1 U879 ( .A(n2458), .B(n2470), .C(n497), .Y(n1621) );
  NAND2X1 U880 ( .A(\mem<10><1> ), .B(n2470), .Y(n497) );
  OAI21X1 U881 ( .A(n2459), .B(n2470), .C(n498), .Y(n1622) );
  NAND2X1 U882 ( .A(\mem<10><2> ), .B(n2470), .Y(n498) );
  OAI21X1 U883 ( .A(n2460), .B(n2470), .C(n499), .Y(n1623) );
  NAND2X1 U884 ( .A(\mem<10><3> ), .B(n2470), .Y(n499) );
  OAI21X1 U885 ( .A(n2461), .B(n2470), .C(n500), .Y(n1624) );
  NAND2X1 U886 ( .A(\mem<10><4> ), .B(n2470), .Y(n500) );
  OAI21X1 U887 ( .A(n2462), .B(n2470), .C(n501), .Y(n1625) );
  NAND2X1 U888 ( .A(\mem<10><5> ), .B(n2470), .Y(n501) );
  OAI21X1 U889 ( .A(n2463), .B(n2470), .C(n502), .Y(n1626) );
  NAND2X1 U890 ( .A(\mem<10><6> ), .B(n2470), .Y(n502) );
  OAI21X1 U891 ( .A(n2464), .B(n2470), .C(n503), .Y(n1627) );
  NAND2X1 U892 ( .A(\mem<10><7> ), .B(n2470), .Y(n503) );
  OAI21X1 U894 ( .A(n2449), .B(n2469), .C(n506), .Y(n1628) );
  NAND2X1 U895 ( .A(\mem<9><0> ), .B(n2469), .Y(n506) );
  OAI21X1 U896 ( .A(n2450), .B(n2469), .C(n507), .Y(n1629) );
  NAND2X1 U897 ( .A(\mem<9><1> ), .B(n2469), .Y(n507) );
  OAI21X1 U898 ( .A(n2451), .B(n2469), .C(n508), .Y(n1630) );
  NAND2X1 U899 ( .A(\mem<9><2> ), .B(n2469), .Y(n508) );
  OAI21X1 U900 ( .A(n2452), .B(n2469), .C(n509), .Y(n1631) );
  NAND2X1 U901 ( .A(\mem<9><3> ), .B(n2469), .Y(n509) );
  OAI21X1 U902 ( .A(n2453), .B(n2469), .C(n510), .Y(n1632) );
  NAND2X1 U903 ( .A(\mem<9><4> ), .B(n2469), .Y(n510) );
  OAI21X1 U904 ( .A(n2454), .B(n2469), .C(n511), .Y(n1633) );
  NAND2X1 U905 ( .A(\mem<9><5> ), .B(n2469), .Y(n511) );
  OAI21X1 U906 ( .A(n2455), .B(n2469), .C(n512), .Y(n1634) );
  NAND2X1 U907 ( .A(\mem<9><6> ), .B(n2469), .Y(n512) );
  OAI21X1 U908 ( .A(n2456), .B(n2469), .C(n513), .Y(n1635) );
  NAND2X1 U909 ( .A(\mem<9><7> ), .B(n2469), .Y(n513) );
  OAI21X1 U910 ( .A(n2457), .B(n2469), .C(n514), .Y(n1636) );
  NAND2X1 U911 ( .A(\mem<8><0> ), .B(n2469), .Y(n514) );
  OAI21X1 U912 ( .A(n2458), .B(n2469), .C(n515), .Y(n1637) );
  NAND2X1 U913 ( .A(\mem<8><1> ), .B(n2469), .Y(n515) );
  OAI21X1 U914 ( .A(n2459), .B(n2469), .C(n516), .Y(n1638) );
  NAND2X1 U915 ( .A(\mem<8><2> ), .B(n2469), .Y(n516) );
  OAI21X1 U916 ( .A(n2460), .B(n2469), .C(n517), .Y(n1639) );
  NAND2X1 U917 ( .A(\mem<8><3> ), .B(n2469), .Y(n517) );
  OAI21X1 U918 ( .A(n2461), .B(n2469), .C(n518), .Y(n1640) );
  NAND2X1 U919 ( .A(\mem<8><4> ), .B(n2469), .Y(n518) );
  OAI21X1 U920 ( .A(n2462), .B(n2469), .C(n519), .Y(n1641) );
  NAND2X1 U921 ( .A(\mem<8><5> ), .B(n2469), .Y(n519) );
  OAI21X1 U922 ( .A(n2463), .B(n2469), .C(n520), .Y(n1642) );
  NAND2X1 U923 ( .A(\mem<8><6> ), .B(n2469), .Y(n520) );
  OAI21X1 U924 ( .A(n2464), .B(n2469), .C(n521), .Y(n1643) );
  NAND2X1 U925 ( .A(\mem<8><7> ), .B(n2469), .Y(n521) );
  OAI21X1 U927 ( .A(n2449), .B(n2468), .C(n524), .Y(n1644) );
  NAND2X1 U928 ( .A(\mem<7><0> ), .B(n2468), .Y(n524) );
  OAI21X1 U929 ( .A(n2450), .B(n2468), .C(n525), .Y(n1645) );
  NAND2X1 U930 ( .A(\mem<7><1> ), .B(n2468), .Y(n525) );
  OAI21X1 U931 ( .A(n2451), .B(n2468), .C(n526), .Y(n1646) );
  NAND2X1 U932 ( .A(\mem<7><2> ), .B(n2468), .Y(n526) );
  OAI21X1 U933 ( .A(n2452), .B(n2468), .C(n527), .Y(n1647) );
  NAND2X1 U934 ( .A(\mem<7><3> ), .B(n2468), .Y(n527) );
  OAI21X1 U935 ( .A(n2453), .B(n2468), .C(n528), .Y(n1648) );
  NAND2X1 U936 ( .A(\mem<7><4> ), .B(n2468), .Y(n528) );
  OAI21X1 U937 ( .A(n2454), .B(n2468), .C(n529), .Y(n1649) );
  NAND2X1 U938 ( .A(\mem<7><5> ), .B(n2468), .Y(n529) );
  OAI21X1 U939 ( .A(n2455), .B(n2468), .C(n530), .Y(n1650) );
  NAND2X1 U940 ( .A(\mem<7><6> ), .B(n2468), .Y(n530) );
  OAI21X1 U941 ( .A(n2456), .B(n2468), .C(n531), .Y(n1651) );
  NAND2X1 U942 ( .A(\mem<7><7> ), .B(n2468), .Y(n531) );
  OAI21X1 U943 ( .A(n2457), .B(n2468), .C(n532), .Y(n1652) );
  NAND2X1 U944 ( .A(\mem<6><0> ), .B(n2468), .Y(n532) );
  OAI21X1 U945 ( .A(n2458), .B(n2468), .C(n533), .Y(n1653) );
  NAND2X1 U946 ( .A(\mem<6><1> ), .B(n2468), .Y(n533) );
  OAI21X1 U947 ( .A(n2459), .B(n2468), .C(n534), .Y(n1654) );
  NAND2X1 U948 ( .A(\mem<6><2> ), .B(n2468), .Y(n534) );
  OAI21X1 U949 ( .A(n2460), .B(n2468), .C(n535), .Y(n1655) );
  NAND2X1 U950 ( .A(\mem<6><3> ), .B(n2468), .Y(n535) );
  OAI21X1 U951 ( .A(n2461), .B(n2468), .C(n536), .Y(n1656) );
  NAND2X1 U952 ( .A(\mem<6><4> ), .B(n2468), .Y(n536) );
  OAI21X1 U953 ( .A(n2462), .B(n2468), .C(n537), .Y(n1657) );
  NAND2X1 U954 ( .A(\mem<6><5> ), .B(n2468), .Y(n537) );
  OAI21X1 U955 ( .A(n2463), .B(n2468), .C(n538), .Y(n1658) );
  NAND2X1 U956 ( .A(\mem<6><6> ), .B(n2468), .Y(n538) );
  OAI21X1 U957 ( .A(n2464), .B(n2468), .C(n539), .Y(n1659) );
  NAND2X1 U958 ( .A(\mem<6><7> ), .B(n2468), .Y(n539) );
  OAI21X1 U960 ( .A(n2449), .B(n2467), .C(n542), .Y(n1660) );
  NAND2X1 U961 ( .A(\mem<5><0> ), .B(n2467), .Y(n542) );
  OAI21X1 U962 ( .A(n2450), .B(n2467), .C(n543), .Y(n1661) );
  NAND2X1 U963 ( .A(\mem<5><1> ), .B(n2467), .Y(n543) );
  OAI21X1 U964 ( .A(n2451), .B(n2467), .C(n544), .Y(n1662) );
  NAND2X1 U965 ( .A(\mem<5><2> ), .B(n2467), .Y(n544) );
  OAI21X1 U966 ( .A(n2452), .B(n2467), .C(n545), .Y(n1663) );
  NAND2X1 U967 ( .A(\mem<5><3> ), .B(n2467), .Y(n545) );
  OAI21X1 U968 ( .A(n2453), .B(n2467), .C(n546), .Y(n1664) );
  NAND2X1 U969 ( .A(\mem<5><4> ), .B(n2467), .Y(n546) );
  OAI21X1 U970 ( .A(n2454), .B(n2467), .C(n547), .Y(n1665) );
  NAND2X1 U971 ( .A(\mem<5><5> ), .B(n2467), .Y(n547) );
  OAI21X1 U972 ( .A(n2455), .B(n2467), .C(n548), .Y(n1666) );
  NAND2X1 U973 ( .A(\mem<5><6> ), .B(n2467), .Y(n548) );
  OAI21X1 U974 ( .A(n2456), .B(n2467), .C(n549), .Y(n1667) );
  NAND2X1 U975 ( .A(\mem<5><7> ), .B(n2467), .Y(n549) );
  OAI21X1 U976 ( .A(n2457), .B(n2467), .C(n550), .Y(n1668) );
  NAND2X1 U977 ( .A(\mem<4><0> ), .B(n2467), .Y(n550) );
  OAI21X1 U978 ( .A(n2458), .B(n2467), .C(n551), .Y(n1669) );
  NAND2X1 U979 ( .A(\mem<4><1> ), .B(n2467), .Y(n551) );
  OAI21X1 U980 ( .A(n2459), .B(n2467), .C(n552), .Y(n1670) );
  NAND2X1 U981 ( .A(\mem<4><2> ), .B(n2467), .Y(n552) );
  OAI21X1 U982 ( .A(n2460), .B(n2467), .C(n553), .Y(n1671) );
  NAND2X1 U983 ( .A(\mem<4><3> ), .B(n2467), .Y(n553) );
  OAI21X1 U984 ( .A(n2461), .B(n2467), .C(n554), .Y(n1672) );
  NAND2X1 U985 ( .A(\mem<4><4> ), .B(n2467), .Y(n554) );
  OAI21X1 U986 ( .A(n2462), .B(n2467), .C(n555), .Y(n1673) );
  NAND2X1 U987 ( .A(\mem<4><5> ), .B(n2467), .Y(n555) );
  OAI21X1 U988 ( .A(n2463), .B(n2467), .C(n556), .Y(n1674) );
  NAND2X1 U989 ( .A(\mem<4><6> ), .B(n2467), .Y(n556) );
  OAI21X1 U990 ( .A(n2464), .B(n2467), .C(n557), .Y(n1675) );
  NAND2X1 U991 ( .A(\mem<4><7> ), .B(n2467), .Y(n557) );
  OAI21X1 U993 ( .A(n2449), .B(n2466), .C(n560), .Y(n1676) );
  NAND2X1 U994 ( .A(\mem<3><0> ), .B(n2466), .Y(n560) );
  OAI21X1 U995 ( .A(n2450), .B(n2466), .C(n561), .Y(n1677) );
  NAND2X1 U996 ( .A(\mem<3><1> ), .B(n2466), .Y(n561) );
  OAI21X1 U997 ( .A(n2451), .B(n2466), .C(n562), .Y(n1678) );
  NAND2X1 U998 ( .A(\mem<3><2> ), .B(n2466), .Y(n562) );
  OAI21X1 U999 ( .A(n2452), .B(n2466), .C(n563), .Y(n1679) );
  NAND2X1 U1000 ( .A(\mem<3><3> ), .B(n2466), .Y(n563) );
  OAI21X1 U1001 ( .A(n2453), .B(n2466), .C(n564), .Y(n1680) );
  NAND2X1 U1002 ( .A(\mem<3><4> ), .B(n2466), .Y(n564) );
  OAI21X1 U1003 ( .A(n2454), .B(n2466), .C(n565), .Y(n1681) );
  NAND2X1 U1004 ( .A(\mem<3><5> ), .B(n2466), .Y(n565) );
  OAI21X1 U1005 ( .A(n2455), .B(n2466), .C(n566), .Y(n1682) );
  NAND2X1 U1006 ( .A(\mem<3><6> ), .B(n2466), .Y(n566) );
  OAI21X1 U1007 ( .A(n2456), .B(n2466), .C(n567), .Y(n1683) );
  NAND2X1 U1008 ( .A(\mem<3><7> ), .B(n2466), .Y(n567) );
  OAI21X1 U1009 ( .A(n2457), .B(n2466), .C(n568), .Y(n1684) );
  NAND2X1 U1010 ( .A(\mem<2><0> ), .B(n2466), .Y(n568) );
  OAI21X1 U1011 ( .A(n2458), .B(n2466), .C(n569), .Y(n1685) );
  NAND2X1 U1012 ( .A(\mem<2><1> ), .B(n2466), .Y(n569) );
  OAI21X1 U1013 ( .A(n2459), .B(n2466), .C(n570), .Y(n1686) );
  NAND2X1 U1014 ( .A(\mem<2><2> ), .B(n2466), .Y(n570) );
  OAI21X1 U1015 ( .A(n2460), .B(n2466), .C(n571), .Y(n1687) );
  NAND2X1 U1016 ( .A(\mem<2><3> ), .B(n2466), .Y(n571) );
  OAI21X1 U1017 ( .A(n2461), .B(n2466), .C(n572), .Y(n1688) );
  NAND2X1 U1018 ( .A(\mem<2><4> ), .B(n2466), .Y(n572) );
  OAI21X1 U1019 ( .A(n2462), .B(n2466), .C(n573), .Y(n1689) );
  NAND2X1 U1020 ( .A(\mem<2><5> ), .B(n2466), .Y(n573) );
  OAI21X1 U1021 ( .A(n2463), .B(n2466), .C(n574), .Y(n1690) );
  NAND2X1 U1022 ( .A(\mem<2><6> ), .B(n2466), .Y(n574) );
  OAI21X1 U1023 ( .A(n2464), .B(n2466), .C(n575), .Y(n1691) );
  NAND2X1 U1024 ( .A(\mem<2><7> ), .B(n2466), .Y(n575) );
  OAI21X1 U1026 ( .A(n2449), .B(n2465), .C(n578), .Y(n1692) );
  NAND2X1 U1027 ( .A(\mem<1><0> ), .B(n2465), .Y(n578) );
  OAI21X1 U1029 ( .A(n2450), .B(n2465), .C(n579), .Y(n1693) );
  NAND2X1 U1030 ( .A(\mem<1><1> ), .B(n2465), .Y(n579) );
  OAI21X1 U1032 ( .A(n2451), .B(n2465), .C(n580), .Y(n1694) );
  NAND2X1 U1033 ( .A(\mem<1><2> ), .B(n2465), .Y(n580) );
  OAI21X1 U1035 ( .A(n2452), .B(n2465), .C(n581), .Y(n1695) );
  NAND2X1 U1036 ( .A(\mem<1><3> ), .B(n2465), .Y(n581) );
  OAI21X1 U1038 ( .A(n2453), .B(n2465), .C(n582), .Y(n1696) );
  NAND2X1 U1039 ( .A(\mem<1><4> ), .B(n2465), .Y(n582) );
  OAI21X1 U1041 ( .A(n2454), .B(n2465), .C(n583), .Y(n1697) );
  NAND2X1 U1042 ( .A(\mem<1><5> ), .B(n2465), .Y(n583) );
  OAI21X1 U1044 ( .A(n2455), .B(n2465), .C(n584), .Y(n1698) );
  NAND2X1 U1045 ( .A(\mem<1><6> ), .B(n2465), .Y(n584) );
  OAI21X1 U1047 ( .A(n2456), .B(n2465), .C(n585), .Y(n1699) );
  NAND2X1 U1048 ( .A(\mem<1><7> ), .B(n2465), .Y(n585) );
  OAI21X1 U1050 ( .A(n2457), .B(n2465), .C(n586), .Y(n1700) );
  NAND2X1 U1051 ( .A(\mem<0><0> ), .B(n2465), .Y(n586) );
  OAI21X1 U1053 ( .A(n2458), .B(n2465), .C(n587), .Y(n1701) );
  NAND2X1 U1054 ( .A(\mem<0><1> ), .B(n2465), .Y(n587) );
  OAI21X1 U1056 ( .A(n2459), .B(n2465), .C(n588), .Y(n1702) );
  NAND2X1 U1057 ( .A(\mem<0><2> ), .B(n2465), .Y(n588) );
  OAI21X1 U1059 ( .A(n2460), .B(n2465), .C(n589), .Y(n1703) );
  NAND2X1 U1060 ( .A(\mem<0><3> ), .B(n2465), .Y(n589) );
  OAI21X1 U1062 ( .A(n2461), .B(n2465), .C(n590), .Y(n1704) );
  NAND2X1 U1063 ( .A(\mem<0><4> ), .B(n2465), .Y(n590) );
  OAI21X1 U1065 ( .A(n2462), .B(n2465), .C(n591), .Y(n1705) );
  NAND2X1 U1066 ( .A(\mem<0><5> ), .B(n2465), .Y(n591) );
  OAI21X1 U1068 ( .A(n2463), .B(n2465), .C(n592), .Y(n1706) );
  NAND2X1 U1069 ( .A(\mem<0><6> ), .B(n2465), .Y(n592) );
  OAI21X1 U1071 ( .A(n2464), .B(n2465), .C(n593), .Y(n1707) );
  NAND2X1 U1072 ( .A(\mem<0><7> ), .B(n2465), .Y(n593) );
  NOR3X1 U1074 ( .A(n2546), .B(n2533), .C(n2548), .Y(n36) );
  OAI21X1 U1076 ( .A(n2533), .B(n2579), .C(n598), .Y(n1162) );
  NAND2X1 U1077 ( .A(n2535), .B(\rand_pat<1> ), .Y(n598) );
  OAI21X1 U1079 ( .A(n2533), .B(n2578), .C(n600), .Y(n1163) );
  NAND2X1 U1080 ( .A(\rand_pat<2> ), .B(n2535), .Y(n600) );
  OAI21X1 U1082 ( .A(n2533), .B(n2577), .C(n602), .Y(n1164) );
  NAND2X1 U1083 ( .A(\rand_pat<3> ), .B(n2535), .Y(n602) );
  OAI21X1 U1085 ( .A(n2533), .B(n2576), .C(n604), .Y(n1165) );
  NAND2X1 U1086 ( .A(\rand_pat<4> ), .B(n2535), .Y(n604) );
  OAI21X1 U1088 ( .A(n2534), .B(n2575), .C(n606), .Y(n1166) );
  NAND2X1 U1089 ( .A(\rand_pat<5> ), .B(n2535), .Y(n606) );
  OAI21X1 U1091 ( .A(n2534), .B(n2574), .C(n608), .Y(n1167) );
  NAND2X1 U1092 ( .A(\rand_pat<6> ), .B(n2535), .Y(n608) );
  OAI21X1 U1094 ( .A(n2534), .B(n2573), .C(n610), .Y(n1168) );
  NAND2X1 U1095 ( .A(\rand_pat<7> ), .B(n2535), .Y(n610) );
  OAI21X1 U1097 ( .A(n2534), .B(n2572), .C(n612), .Y(n1169) );
  NAND2X1 U1098 ( .A(\rand_pat<8> ), .B(n2535), .Y(n612) );
  OAI21X1 U1100 ( .A(n2534), .B(n2571), .C(n614), .Y(n1170) );
  NAND2X1 U1101 ( .A(\rand_pat<9> ), .B(n2535), .Y(n614) );
  OAI21X1 U1103 ( .A(n2534), .B(n2570), .C(n616), .Y(n1171) );
  NAND2X1 U1104 ( .A(\rand_pat<10> ), .B(n2535), .Y(n616) );
  OAI21X1 U1106 ( .A(n2534), .B(n2569), .C(n618), .Y(n1172) );
  NAND2X1 U1107 ( .A(\rand_pat<11> ), .B(n2535), .Y(n618) );
  OAI21X1 U1109 ( .A(n2534), .B(n2568), .C(n620), .Y(n1173) );
  NAND2X1 U1110 ( .A(\rand_pat<12> ), .B(n2535), .Y(n620) );
  OAI21X1 U1112 ( .A(n2534), .B(n2567), .C(n622), .Y(n1174) );
  NAND2X1 U1113 ( .A(\rand_pat<13> ), .B(n2535), .Y(n622) );
  OAI21X1 U1115 ( .A(n2534), .B(n2566), .C(n624), .Y(n1175) );
  NAND2X1 U1116 ( .A(\rand_pat<14> ), .B(n2535), .Y(n624) );
  OAI21X1 U1118 ( .A(n2534), .B(n2565), .C(n626), .Y(n1176) );
  NAND2X1 U1119 ( .A(\rand_pat<15> ), .B(n2535), .Y(n626) );
  OAI21X1 U1121 ( .A(n2534), .B(n2564), .C(n628), .Y(n1177) );
  NAND2X1 U1122 ( .A(\rand_pat<16> ), .B(n2535), .Y(n628) );
  OAI21X1 U1124 ( .A(n2534), .B(n2563), .C(n630), .Y(n1178) );
  NAND2X1 U1125 ( .A(\rand_pat<17> ), .B(n2535), .Y(n630) );
  OAI21X1 U1127 ( .A(n2534), .B(n2562), .C(n632), .Y(n1179) );
  NAND2X1 U1128 ( .A(\rand_pat<18> ), .B(n2535), .Y(n632) );
  OAI21X1 U1130 ( .A(n2534), .B(n2561), .C(n634), .Y(n1180) );
  NAND2X1 U1131 ( .A(\rand_pat<19> ), .B(n2535), .Y(n634) );
  OAI21X1 U1133 ( .A(n2534), .B(n2560), .C(n636), .Y(n1181) );
  NAND2X1 U1134 ( .A(\rand_pat<20> ), .B(n2535), .Y(n636) );
  OAI21X1 U1136 ( .A(n2534), .B(n2559), .C(n638), .Y(n1182) );
  NAND2X1 U1137 ( .A(\rand_pat<21> ), .B(n2535), .Y(n638) );
  OAI21X1 U1139 ( .A(n2534), .B(n2558), .C(n640), .Y(n1183) );
  NAND2X1 U1140 ( .A(\rand_pat<22> ), .B(n2535), .Y(n640) );
  OAI21X1 U1142 ( .A(n2534), .B(n2557), .C(n642), .Y(n1184) );
  NAND2X1 U1143 ( .A(\rand_pat<23> ), .B(n2535), .Y(n642) );
  OAI21X1 U1145 ( .A(n2533), .B(n2556), .C(n644), .Y(n1185) );
  NAND2X1 U1146 ( .A(\rand_pat<24> ), .B(n2535), .Y(n644) );
  OAI21X1 U1148 ( .A(n2533), .B(n2555), .C(n646), .Y(n1186) );
  NAND2X1 U1149 ( .A(\rand_pat<25> ), .B(n2535), .Y(n646) );
  OAI21X1 U1151 ( .A(n2533), .B(n2554), .C(n648), .Y(n1187) );
  NAND2X1 U1152 ( .A(\rand_pat<26> ), .B(n2535), .Y(n648) );
  OAI21X1 U1154 ( .A(n2533), .B(n2553), .C(n650), .Y(n1188) );
  NAND2X1 U1155 ( .A(\rand_pat<27> ), .B(n2535), .Y(n650) );
  OAI21X1 U1157 ( .A(n2533), .B(n2552), .C(n652), .Y(n1189) );
  NAND2X1 U1158 ( .A(\rand_pat<28> ), .B(n2535), .Y(n652) );
  OAI21X1 U1160 ( .A(n2533), .B(n2551), .C(n654), .Y(n1190) );
  NAND2X1 U1161 ( .A(\rand_pat<29> ), .B(n2535), .Y(n654) );
  OAI21X1 U1163 ( .A(n2533), .B(n2550), .C(n656), .Y(n1191) );
  NAND2X1 U1164 ( .A(\rand_pat<30> ), .B(n2534), .Y(n656) );
  OAI21X1 U1166 ( .A(n2533), .B(n2549), .C(n658), .Y(n1192) );
  NAND2X1 U1167 ( .A(\rand_pat<31> ), .B(n2535), .Y(n658) );
  OAI21X1 U1168 ( .A(n2533), .B(n2580), .C(n660), .Y(n1193) );
  NAND2X1 U1169 ( .A(n2535), .B(\rand_pat<0> ), .Y(n660) );
  AOI21X1 U1171 ( .A(n2548), .B(n2547), .C(\rand_pat<0> ), .Y(n2581) );
  OAI21X1 U1172 ( .A(n662), .B(n2448), .C(n1099), .Y(\DataOut<9> ) );
  NOR3X1 U1174 ( .A(n666), .B(n739), .C(n915), .Y(n662) );
  AOI22X1 U1177 ( .A(n674), .B(\mem<34><1> ), .C(n675), .D(\mem<32><1> ), .Y(
        n673) );
  AOI22X1 U1178 ( .A(n676), .B(\mem<38><1> ), .C(n677), .D(\mem<36><1> ), .Y(
        n672) );
  AOI22X1 U1179 ( .A(n678), .B(\mem<42><1> ), .C(n679), .D(\mem<40><1> ), .Y(
        n670) );
  AOI22X1 U1180 ( .A(n680), .B(\mem<46><1> ), .C(n681), .D(\mem<44><1> ), .Y(
        n669) );
  AOI22X1 U1183 ( .A(n687), .B(\mem<58><1> ), .C(n688), .D(\mem<56><1> ), .Y(
        n686) );
  AOI22X1 U1184 ( .A(n689), .B(\mem<62><1> ), .C(n690), .D(\mem<60><1> ), .Y(
        n685) );
  AOI22X1 U1185 ( .A(n691), .B(\mem<50><1> ), .C(n692), .D(\mem<48><1> ), .Y(
        n683) );
  AOI22X1 U1186 ( .A(n693), .B(\mem<54><1> ), .C(n694), .D(\mem<52><1> ), .Y(
        n682) );
  AOI22X1 U1190 ( .A(n702), .B(\mem<2><1> ), .C(n703), .D(\mem<0><1> ), .Y(
        n701) );
  AOI22X1 U1191 ( .A(n704), .B(\mem<6><1> ), .C(n705), .D(\mem<4><1> ), .Y(
        n700) );
  AOI22X1 U1192 ( .A(n706), .B(\mem<10><1> ), .C(n707), .D(\mem<8><1> ), .Y(
        n698) );
  AOI22X1 U1193 ( .A(n708), .B(\mem<14><1> ), .C(n709), .D(\mem<12><1> ), .Y(
        n697) );
  AOI22X1 U1196 ( .A(n715), .B(\mem<18><1> ), .C(n716), .D(\mem<16><1> ), .Y(
        n714) );
  AOI22X1 U1197 ( .A(n717), .B(\mem<22><1> ), .C(n718), .D(\mem<20><1> ), .Y(
        n713) );
  AOI22X1 U1198 ( .A(n719), .B(\mem<26><1> ), .C(n720), .D(\mem<24><1> ), .Y(
        n711) );
  AOI22X1 U1199 ( .A(n721), .B(\mem<30><1> ), .C(n722), .D(\mem<28><1> ), .Y(
        n710) );
  OAI21X1 U1200 ( .A(n723), .B(n2448), .C(n1079), .Y(\DataOut<8> ) );
  NOR3X1 U1202 ( .A(n725), .B(n727), .C(n902), .Y(n723) );
  AOI22X1 U1205 ( .A(n674), .B(\mem<34><0> ), .C(n675), .D(\mem<32><0> ), .Y(
        n732) );
  AOI22X1 U1206 ( .A(n676), .B(\mem<38><0> ), .C(n677), .D(\mem<36><0> ), .Y(
        n731) );
  AOI22X1 U1207 ( .A(n678), .B(\mem<42><0> ), .C(n679), .D(\mem<40><0> ), .Y(
        n729) );
  AOI22X1 U1208 ( .A(n680), .B(\mem<46><0> ), .C(n681), .D(\mem<44><0> ), .Y(
        n728) );
  AOI22X1 U1211 ( .A(n687), .B(\mem<58><0> ), .C(n688), .D(\mem<56><0> ), .Y(
        n737) );
  AOI22X1 U1212 ( .A(n689), .B(\mem<62><0> ), .C(n690), .D(\mem<60><0> ), .Y(
        n736) );
  AOI22X1 U1213 ( .A(n691), .B(\mem<50><0> ), .C(n692), .D(\mem<48><0> ), .Y(
        n734) );
  AOI22X1 U1214 ( .A(n693), .B(\mem<54><0> ), .C(n694), .D(\mem<52><0> ), .Y(
        n733) );
  AOI22X1 U1218 ( .A(n702), .B(\mem<2><0> ), .C(n703), .D(\mem<0><0> ), .Y(
        n744) );
  AOI22X1 U1219 ( .A(n704), .B(\mem<6><0> ), .C(n705), .D(\mem<4><0> ), .Y(
        n743) );
  AOI22X1 U1220 ( .A(n706), .B(\mem<10><0> ), .C(n707), .D(\mem<8><0> ), .Y(
        n741) );
  AOI22X1 U1221 ( .A(n708), .B(\mem<14><0> ), .C(n709), .D(\mem<12><0> ), .Y(
        n740) );
  AOI22X1 U1224 ( .A(n715), .B(\mem<18><0> ), .C(n716), .D(\mem<16><0> ), .Y(
        n749) );
  AOI22X1 U1225 ( .A(n717), .B(\mem<22><0> ), .C(n718), .D(\mem<20><0> ), .Y(
        n748) );
  AOI22X1 U1226 ( .A(n719), .B(\mem<26><0> ), .C(n720), .D(\mem<24><0> ), .Y(
        n746) );
  AOI22X1 U1227 ( .A(n721), .B(\mem<30><0> ), .C(n722), .D(\mem<28><0> ), .Y(
        n745) );
  OAI21X1 U1228 ( .A(n750), .B(n2447), .C(n1065), .Y(\DataOut<7> ) );
  NOR3X1 U1230 ( .A(n754), .B(n724), .C(n890), .Y(n750) );
  AOI22X1 U1233 ( .A(\mem<29><7> ), .B(n342), .C(\mem<31><7> ), .D(n324), .Y(
        n761) );
  AOI22X1 U1234 ( .A(\mem<25><7> ), .B(n378), .C(\mem<27><7> ), .D(n360), .Y(
        n760) );
  AOI22X1 U1235 ( .A(\mem<21><7> ), .B(n414), .C(\mem<23><7> ), .D(n396), .Y(
        n758) );
  AOI22X1 U1236 ( .A(\mem<17><7> ), .B(n450), .C(\mem<19><7> ), .D(n432), .Y(
        n757) );
  AOI22X1 U1239 ( .A(\mem<13><7> ), .B(n486), .C(\mem<15><7> ), .D(n468), .Y(
        n766) );
  AOI22X1 U1240 ( .A(\mem<9><7> ), .B(n522), .C(\mem<11><7> ), .D(n504), .Y(
        n765) );
  AOI22X1 U1241 ( .A(\mem<5><7> ), .B(n558), .C(\mem<7><7> ), .D(n540), .Y(
        n763) );
  AOI22X1 U1242 ( .A(\mem<1><7> ), .B(n594), .C(\mem<3><7> ), .D(n576), .Y(
        n762) );
  AOI22X1 U1246 ( .A(\mem<61><7> ), .B(n54), .C(\mem<63><7> ), .D(n35), .Y(
        n773) );
  AOI22X1 U1247 ( .A(\mem<57><7> ), .B(n90), .C(\mem<59><7> ), .D(n72), .Y(
        n772) );
  AOI22X1 U1248 ( .A(\mem<53><7> ), .B(n126), .C(\mem<55><7> ), .D(n108), .Y(
        n770) );
  AOI22X1 U1249 ( .A(\mem<49><7> ), .B(n162), .C(\mem<51><7> ), .D(n144), .Y(
        n769) );
  AOI22X1 U1252 ( .A(\mem<45><7> ), .B(n198), .C(\mem<47><7> ), .D(n180), .Y(
        n778) );
  AOI22X1 U1253 ( .A(\mem<41><7> ), .B(n234), .C(\mem<43><7> ), .D(n216), .Y(
        n777) );
  AOI22X1 U1254 ( .A(\mem<37><7> ), .B(n270), .C(\mem<39><7> ), .D(n252), .Y(
        n775) );
  AOI22X1 U1255 ( .A(\mem<33><7> ), .B(n306), .C(\mem<35><7> ), .D(n288), .Y(
        n774) );
  OAI21X1 U1256 ( .A(n779), .B(n2447), .C(n1053), .Y(\DataOut<6> ) );
  NOR3X1 U1258 ( .A(n781), .B(n695), .C(n876), .Y(n779) );
  AOI22X1 U1261 ( .A(\mem<29><6> ), .B(n342), .C(\mem<31><6> ), .D(n324), .Y(
        n788) );
  AOI22X1 U1262 ( .A(\mem<25><6> ), .B(n378), .C(\mem<27><6> ), .D(n360), .Y(
        n787) );
  AOI22X1 U1263 ( .A(\mem<21><6> ), .B(n414), .C(\mem<23><6> ), .D(n396), .Y(
        n785) );
  AOI22X1 U1264 ( .A(\mem<17><6> ), .B(n450), .C(\mem<19><6> ), .D(n432), .Y(
        n784) );
  AOI22X1 U1267 ( .A(\mem<13><6> ), .B(n486), .C(\mem<15><6> ), .D(n468), .Y(
        n793) );
  AOI22X1 U1268 ( .A(\mem<9><6> ), .B(n522), .C(\mem<11><6> ), .D(n504), .Y(
        n792) );
  AOI22X1 U1269 ( .A(\mem<5><6> ), .B(n558), .C(\mem<7><6> ), .D(n540), .Y(
        n790) );
  AOI22X1 U1270 ( .A(\mem<1><6> ), .B(n594), .C(\mem<3><6> ), .D(n576), .Y(
        n789) );
  AOI22X1 U1274 ( .A(\mem<61><6> ), .B(n54), .C(\mem<63><6> ), .D(n35), .Y(
        n800) );
  AOI22X1 U1275 ( .A(\mem<57><6> ), .B(n90), .C(\mem<59><6> ), .D(n72), .Y(
        n799) );
  AOI22X1 U1276 ( .A(\mem<53><6> ), .B(n126), .C(\mem<55><6> ), .D(n108), .Y(
        n797) );
  AOI22X1 U1277 ( .A(\mem<49><6> ), .B(n162), .C(\mem<51><6> ), .D(n144), .Y(
        n796) );
  AOI22X1 U1280 ( .A(\mem<45><6> ), .B(n198), .C(\mem<47><6> ), .D(n180), .Y(
        n805) );
  AOI22X1 U1281 ( .A(\mem<41><6> ), .B(n234), .C(\mem<43><6> ), .D(n216), .Y(
        n804) );
  AOI22X1 U1282 ( .A(\mem<37><6> ), .B(n270), .C(\mem<39><6> ), .D(n252), .Y(
        n802) );
  AOI22X1 U1283 ( .A(\mem<33><6> ), .B(n306), .C(\mem<35><6> ), .D(n288), .Y(
        n801) );
  OAI21X1 U1284 ( .A(n806), .B(n2447), .C(n1050), .Y(\DataOut<5> ) );
  NOR3X1 U1286 ( .A(n808), .B(n667), .C(n864), .Y(n806) );
  AOI22X1 U1289 ( .A(\mem<29><5> ), .B(n342), .C(\mem<31><5> ), .D(n324), .Y(
        n815) );
  AOI22X1 U1290 ( .A(\mem<25><5> ), .B(n378), .C(\mem<27><5> ), .D(n360), .Y(
        n814) );
  AOI22X1 U1291 ( .A(\mem<21><5> ), .B(n414), .C(\mem<23><5> ), .D(n396), .Y(
        n812) );
  AOI22X1 U1292 ( .A(\mem<17><5> ), .B(n450), .C(\mem<19><5> ), .D(n432), .Y(
        n811) );
  AOI22X1 U1295 ( .A(\mem<13><5> ), .B(n486), .C(\mem<15><5> ), .D(n468), .Y(
        n820) );
  AOI22X1 U1296 ( .A(\mem<9><5> ), .B(n522), .C(\mem<11><5> ), .D(n504), .Y(
        n819) );
  AOI22X1 U1297 ( .A(\mem<5><5> ), .B(n558), .C(\mem<7><5> ), .D(n540), .Y(
        n817) );
  AOI22X1 U1298 ( .A(\mem<1><5> ), .B(n594), .C(\mem<3><5> ), .D(n576), .Y(
        n816) );
  AOI22X1 U1302 ( .A(\mem<61><5> ), .B(n54), .C(\mem<63><5> ), .D(n35), .Y(
        n827) );
  AOI22X1 U1303 ( .A(\mem<57><5> ), .B(n90), .C(\mem<59><5> ), .D(n72), .Y(
        n826) );
  AOI22X1 U1304 ( .A(\mem<53><5> ), .B(n126), .C(\mem<55><5> ), .D(n108), .Y(
        n824) );
  AOI22X1 U1305 ( .A(\mem<49><5> ), .B(n162), .C(\mem<51><5> ), .D(n144), .Y(
        n823) );
  AOI22X1 U1308 ( .A(\mem<45><5> ), .B(n198), .C(\mem<47><5> ), .D(n180), .Y(
        n832) );
  AOI22X1 U1309 ( .A(\mem<41><5> ), .B(n234), .C(\mem<43><5> ), .D(n216), .Y(
        n831) );
  AOI22X1 U1310 ( .A(\mem<37><5> ), .B(n270), .C(\mem<39><5> ), .D(n252), .Y(
        n829) );
  AOI22X1 U1311 ( .A(\mem<33><5> ), .B(n306), .C(\mem<35><5> ), .D(n288), .Y(
        n828) );
  OAI21X1 U1312 ( .A(n833), .B(n2447), .C(n1037), .Y(\DataOut<4> ) );
  NOR3X1 U1314 ( .A(n835), .B(n664), .C(n861), .Y(n833) );
  AOI22X1 U1317 ( .A(\mem<29><4> ), .B(n342), .C(\mem<31><4> ), .D(n324), .Y(
        n842) );
  AOI22X1 U1318 ( .A(\mem<25><4> ), .B(n378), .C(\mem<27><4> ), .D(n360), .Y(
        n841) );
  AOI22X1 U1319 ( .A(\mem<21><4> ), .B(n414), .C(\mem<23><4> ), .D(n396), .Y(
        n839) );
  AOI22X1 U1320 ( .A(\mem<17><4> ), .B(n450), .C(\mem<19><4> ), .D(n432), .Y(
        n838) );
  AOI22X1 U1323 ( .A(\mem<13><4> ), .B(n486), .C(\mem<15><4> ), .D(n468), .Y(
        n847) );
  AOI22X1 U1324 ( .A(\mem<9><4> ), .B(n522), .C(\mem<11><4> ), .D(n504), .Y(
        n846) );
  AOI22X1 U1325 ( .A(\mem<5><4> ), .B(n558), .C(\mem<7><4> ), .D(n540), .Y(
        n844) );
  AOI22X1 U1326 ( .A(\mem<1><4> ), .B(n594), .C(\mem<3><4> ), .D(n576), .Y(
        n843) );
  AOI22X1 U1330 ( .A(\mem<61><4> ), .B(n54), .C(\mem<63><4> ), .D(n35), .Y(
        n854) );
  AOI22X1 U1331 ( .A(\mem<57><4> ), .B(n90), .C(\mem<59><4> ), .D(n72), .Y(
        n853) );
  AOI22X1 U1332 ( .A(\mem<53><4> ), .B(n126), .C(\mem<55><4> ), .D(n108), .Y(
        n851) );
  AOI22X1 U1333 ( .A(\mem<49><4> ), .B(n162), .C(\mem<51><4> ), .D(n144), .Y(
        n850) );
  AOI22X1 U1336 ( .A(\mem<45><4> ), .B(n198), .C(\mem<47><4> ), .D(n180), .Y(
        n859) );
  AOI22X1 U1337 ( .A(\mem<41><4> ), .B(n234), .C(\mem<43><4> ), .D(n216), .Y(
        n858) );
  AOI22X1 U1338 ( .A(\mem<37><4> ), .B(n270), .C(\mem<39><4> ), .D(n252), .Y(
        n856) );
  AOI22X1 U1339 ( .A(\mem<33><4> ), .B(n306), .C(\mem<35><4> ), .D(n288), .Y(
        n855) );
  OAI21X1 U1340 ( .A(n860), .B(n2447), .C(n1025), .Y(\DataOut<3> ) );
  NOR3X1 U1342 ( .A(n862), .B(n659), .C(n848), .Y(n860) );
  AOI22X1 U1345 ( .A(\mem<29><3> ), .B(n342), .C(\mem<31><3> ), .D(n324), .Y(
        n869) );
  AOI22X1 U1346 ( .A(\mem<25><3> ), .B(n378), .C(\mem<27><3> ), .D(n360), .Y(
        n868) );
  AOI22X1 U1347 ( .A(\mem<21><3> ), .B(n414), .C(\mem<23><3> ), .D(n396), .Y(
        n866) );
  AOI22X1 U1348 ( .A(\mem<17><3> ), .B(n450), .C(\mem<19><3> ), .D(n432), .Y(
        n865) );
  AOI22X1 U1351 ( .A(\mem<13><3> ), .B(n486), .C(\mem<15><3> ), .D(n468), .Y(
        n874) );
  AOI22X1 U1352 ( .A(\mem<9><3> ), .B(n522), .C(\mem<11><3> ), .D(n504), .Y(
        n873) );
  AOI22X1 U1353 ( .A(\mem<5><3> ), .B(n558), .C(\mem<7><3> ), .D(n540), .Y(
        n871) );
  AOI22X1 U1354 ( .A(\mem<1><3> ), .B(n594), .C(\mem<3><3> ), .D(n576), .Y(
        n870) );
  AOI22X1 U1358 ( .A(\mem<61><3> ), .B(n54), .C(\mem<63><3> ), .D(n35), .Y(
        n881) );
  AOI22X1 U1359 ( .A(\mem<57><3> ), .B(n90), .C(\mem<59><3> ), .D(n72), .Y(
        n880) );
  AOI22X1 U1360 ( .A(\mem<53><3> ), .B(n126), .C(\mem<55><3> ), .D(n108), .Y(
        n878) );
  AOI22X1 U1361 ( .A(\mem<49><3> ), .B(n162), .C(\mem<51><3> ), .D(n144), .Y(
        n877) );
  AOI22X1 U1364 ( .A(\mem<45><3> ), .B(n198), .C(\mem<47><3> ), .D(n180), .Y(
        n886) );
  AOI22X1 U1365 ( .A(\mem<41><3> ), .B(n234), .C(\mem<43><3> ), .D(n216), .Y(
        n885) );
  AOI22X1 U1366 ( .A(\mem<37><3> ), .B(n270), .C(\mem<39><3> ), .D(n252), .Y(
        n883) );
  AOI22X1 U1367 ( .A(\mem<33><3> ), .B(n306), .C(\mem<35><3> ), .D(n288), .Y(
        n882) );
  OAI21X1 U1368 ( .A(n887), .B(n2447), .C(n1011), .Y(\DataOut<2> ) );
  NOR3X1 U1370 ( .A(n889), .B(n655), .C(n836), .Y(n887) );
  AOI22X1 U1373 ( .A(\mem<29><2> ), .B(n342), .C(\mem<31><2> ), .D(n324), .Y(
        n896) );
  AOI22X1 U1374 ( .A(\mem<25><2> ), .B(n378), .C(\mem<27><2> ), .D(n360), .Y(
        n895) );
  AOI22X1 U1375 ( .A(\mem<21><2> ), .B(n414), .C(\mem<23><2> ), .D(n396), .Y(
        n893) );
  AOI22X1 U1376 ( .A(\mem<17><2> ), .B(n450), .C(\mem<19><2> ), .D(n432), .Y(
        n892) );
  AOI22X1 U1379 ( .A(\mem<13><2> ), .B(n486), .C(\mem<15><2> ), .D(n468), .Y(
        n901) );
  AOI22X1 U1380 ( .A(\mem<9><2> ), .B(n522), .C(\mem<11><2> ), .D(n504), .Y(
        n900) );
  AOI22X1 U1381 ( .A(\mem<5><2> ), .B(n558), .C(\mem<7><2> ), .D(n540), .Y(
        n898) );
  AOI22X1 U1382 ( .A(\mem<1><2> ), .B(n594), .C(\mem<3><2> ), .D(n576), .Y(
        n897) );
  AOI22X1 U1386 ( .A(\mem<61><2> ), .B(n54), .C(\mem<63><2> ), .D(n35), .Y(
        n908) );
  AOI22X1 U1387 ( .A(\mem<57><2> ), .B(n90), .C(\mem<59><2> ), .D(n72), .Y(
        n907) );
  AOI22X1 U1388 ( .A(\mem<53><2> ), .B(n126), .C(\mem<55><2> ), .D(n108), .Y(
        n905) );
  AOI22X1 U1389 ( .A(\mem<49><2> ), .B(n162), .C(\mem<51><2> ), .D(n144), .Y(
        n904) );
  AOI22X1 U1392 ( .A(\mem<45><2> ), .B(n198), .C(\mem<47><2> ), .D(n180), .Y(
        n913) );
  AOI22X1 U1393 ( .A(\mem<41><2> ), .B(n234), .C(\mem<43><2> ), .D(n216), .Y(
        n912) );
  AOI22X1 U1394 ( .A(\mem<37><2> ), .B(n270), .C(\mem<39><2> ), .D(n252), .Y(
        n910) );
  AOI22X1 U1395 ( .A(\mem<33><2> ), .B(n306), .C(\mem<35><2> ), .D(n288), .Y(
        n909) );
  OAI21X1 U1396 ( .A(n914), .B(n2447), .C(n999), .Y(\DataOut<1> ) );
  NOR3X1 U1398 ( .A(n916), .B(n651), .C(n822), .Y(n914) );
  AOI22X1 U1401 ( .A(\mem<29><1> ), .B(n342), .C(\mem<31><1> ), .D(n324), .Y(
        n923) );
  AOI22X1 U1402 ( .A(\mem<25><1> ), .B(n378), .C(\mem<27><1> ), .D(n360), .Y(
        n922) );
  AOI22X1 U1403 ( .A(\mem<21><1> ), .B(n414), .C(\mem<23><1> ), .D(n396), .Y(
        n920) );
  AOI22X1 U1404 ( .A(\mem<17><1> ), .B(n450), .C(\mem<19><1> ), .D(n432), .Y(
        n919) );
  AOI22X1 U1407 ( .A(\mem<13><1> ), .B(n486), .C(\mem<15><1> ), .D(n468), .Y(
        n928) );
  AOI22X1 U1408 ( .A(\mem<9><1> ), .B(n522), .C(\mem<11><1> ), .D(n504), .Y(
        n927) );
  AOI22X1 U1409 ( .A(\mem<5><1> ), .B(n558), .C(\mem<7><1> ), .D(n540), .Y(
        n925) );
  AOI22X1 U1410 ( .A(\mem<1><1> ), .B(n594), .C(\mem<3><1> ), .D(n576), .Y(
        n924) );
  AOI22X1 U1414 ( .A(\mem<61><1> ), .B(n54), .C(\mem<63><1> ), .D(n35), .Y(
        n935) );
  AOI22X1 U1415 ( .A(\mem<57><1> ), .B(n90), .C(\mem<59><1> ), .D(n72), .Y(
        n934) );
  AOI22X1 U1416 ( .A(\mem<53><1> ), .B(n126), .C(\mem<55><1> ), .D(n108), .Y(
        n932) );
  AOI22X1 U1417 ( .A(\mem<49><1> ), .B(n162), .C(\mem<51><1> ), .D(n144), .Y(
        n931) );
  AOI22X1 U1420 ( .A(\mem<45><1> ), .B(n198), .C(\mem<47><1> ), .D(n180), .Y(
        n940) );
  AOI22X1 U1421 ( .A(\mem<41><1> ), .B(n234), .C(\mem<43><1> ), .D(n216), .Y(
        n939) );
  AOI22X1 U1422 ( .A(\mem<37><1> ), .B(n270), .C(\mem<39><1> ), .D(n252), .Y(
        n937) );
  AOI22X1 U1423 ( .A(\mem<33><1> ), .B(n306), .C(\mem<35><1> ), .D(n288), .Y(
        n936) );
  OAI21X1 U1424 ( .A(n941), .B(n2448), .C(n996), .Y(\DataOut<15> ) );
  NOR3X1 U1426 ( .A(n943), .B(n647), .C(n810), .Y(n941) );
  AOI22X1 U1429 ( .A(n674), .B(\mem<34><7> ), .C(n675), .D(\mem<32><7> ), .Y(
        n950) );
  AOI22X1 U1430 ( .A(n676), .B(\mem<38><7> ), .C(n677), .D(\mem<36><7> ), .Y(
        n949) );
  AOI22X1 U1431 ( .A(n678), .B(\mem<42><7> ), .C(n679), .D(\mem<40><7> ), .Y(
        n947) );
  AOI22X1 U1432 ( .A(n680), .B(\mem<46><7> ), .C(n681), .D(\mem<44><7> ), .Y(
        n946) );
  AOI22X1 U1435 ( .A(n687), .B(\mem<58><7> ), .C(n688), .D(\mem<56><7> ), .Y(
        n955) );
  AOI22X1 U1436 ( .A(n689), .B(\mem<62><7> ), .C(n690), .D(\mem<60><7> ), .Y(
        n954) );
  AOI22X1 U1437 ( .A(n691), .B(\mem<50><7> ), .C(n692), .D(\mem<48><7> ), .Y(
        n952) );
  AOI22X1 U1438 ( .A(n693), .B(\mem<54><7> ), .C(n694), .D(\mem<52><7> ), .Y(
        n951) );
  AOI22X1 U1442 ( .A(n702), .B(\mem<2><7> ), .C(n703), .D(\mem<0><7> ), .Y(
        n962) );
  AOI22X1 U1443 ( .A(n704), .B(\mem<6><7> ), .C(n705), .D(\mem<4><7> ), .Y(
        n961) );
  AOI22X1 U1444 ( .A(n706), .B(\mem<10><7> ), .C(n707), .D(\mem<8><7> ), .Y(
        n959) );
  AOI22X1 U1445 ( .A(n708), .B(\mem<14><7> ), .C(n709), .D(\mem<12><7> ), .Y(
        n958) );
  AOI22X1 U1448 ( .A(n715), .B(\mem<18><7> ), .C(n716), .D(\mem<16><7> ), .Y(
        n967) );
  AOI22X1 U1449 ( .A(n717), .B(\mem<22><7> ), .C(n718), .D(\mem<20><7> ), .Y(
        n966) );
  AOI22X1 U1450 ( .A(n719), .B(\mem<26><7> ), .C(n720), .D(\mem<24><7> ), .Y(
        n964) );
  AOI22X1 U1451 ( .A(n721), .B(\mem<30><7> ), .C(n722), .D(\mem<28><7> ), .Y(
        n963) );
  OAI21X1 U1452 ( .A(n968), .B(n2448), .C(n983), .Y(\DataOut<14> ) );
  NOR3X1 U1454 ( .A(n970), .B(n643), .C(n807), .Y(n968) );
  AOI22X1 U1457 ( .A(n674), .B(\mem<34><6> ), .C(n675), .D(\mem<32><6> ), .Y(
        n977) );
  AOI22X1 U1458 ( .A(n676), .B(\mem<38><6> ), .C(n677), .D(\mem<36><6> ), .Y(
        n976) );
  AOI22X1 U1459 ( .A(n678), .B(\mem<42><6> ), .C(n679), .D(\mem<40><6> ), .Y(
        n974) );
  AOI22X1 U1460 ( .A(n680), .B(\mem<46><6> ), .C(n681), .D(\mem<44><6> ), .Y(
        n973) );
  AOI22X1 U1463 ( .A(n687), .B(\mem<58><6> ), .C(n688), .D(\mem<56><6> ), .Y(
        n982) );
  AOI22X1 U1464 ( .A(n689), .B(\mem<62><6> ), .C(n690), .D(\mem<60><6> ), .Y(
        n981) );
  AOI22X1 U1465 ( .A(n691), .B(\mem<50><6> ), .C(n692), .D(\mem<48><6> ), .Y(
        n979) );
  AOI22X1 U1466 ( .A(n693), .B(\mem<54><6> ), .C(n694), .D(\mem<52><6> ), .Y(
        n978) );
  AOI22X1 U1470 ( .A(n702), .B(\mem<2><6> ), .C(n703), .D(\mem<0><6> ), .Y(
        n989) );
  AOI22X1 U1471 ( .A(n704), .B(\mem<6><6> ), .C(n705), .D(\mem<4><6> ), .Y(
        n988) );
  AOI22X1 U1472 ( .A(n706), .B(\mem<10><6> ), .C(n707), .D(\mem<8><6> ), .Y(
        n986) );
  AOI22X1 U1473 ( .A(n708), .B(\mem<14><6> ), .C(n709), .D(\mem<12><6> ), .Y(
        n985) );
  AOI22X1 U1476 ( .A(n715), .B(\mem<18><6> ), .C(n716), .D(\mem<16><6> ), .Y(
        n994) );
  AOI22X1 U1477 ( .A(n717), .B(\mem<22><6> ), .C(n718), .D(\mem<20><6> ), .Y(
        n993) );
  AOI22X1 U1478 ( .A(n719), .B(\mem<26><6> ), .C(n720), .D(\mem<24><6> ), .Y(
        n991) );
  AOI22X1 U1479 ( .A(n721), .B(\mem<30><6> ), .C(n722), .D(\mem<28><6> ), .Y(
        n990) );
  OAI21X1 U1480 ( .A(n995), .B(n2448), .C(n971), .Y(\DataOut<13> ) );
  NOR3X1 U1482 ( .A(n997), .B(n639), .C(n794), .Y(n995) );
  AOI22X1 U1485 ( .A(n674), .B(\mem<34><5> ), .C(n675), .D(\mem<32><5> ), .Y(
        n1004) );
  AOI22X1 U1486 ( .A(n676), .B(\mem<38><5> ), .C(n677), .D(\mem<36><5> ), .Y(
        n1003) );
  AOI22X1 U1487 ( .A(n678), .B(\mem<42><5> ), .C(n679), .D(\mem<40><5> ), .Y(
        n1001) );
  AOI22X1 U1488 ( .A(n680), .B(\mem<46><5> ), .C(n681), .D(\mem<44><5> ), .Y(
        n1000) );
  AOI22X1 U1491 ( .A(n687), .B(\mem<58><5> ), .C(n688), .D(\mem<56><5> ), .Y(
        n1009) );
  AOI22X1 U1492 ( .A(n689), .B(\mem<62><5> ), .C(n690), .D(\mem<60><5> ), .Y(
        n1008) );
  AOI22X1 U1493 ( .A(n691), .B(\mem<50><5> ), .C(n692), .D(\mem<48><5> ), .Y(
        n1006) );
  AOI22X1 U1494 ( .A(n693), .B(\mem<54><5> ), .C(n694), .D(\mem<52><5> ), .Y(
        n1005) );
  AOI22X1 U1498 ( .A(n702), .B(\mem<2><5> ), .C(n703), .D(\mem<0><5> ), .Y(
        n1016) );
  AOI22X1 U1499 ( .A(n704), .B(\mem<6><5> ), .C(n705), .D(\mem<4><5> ), .Y(
        n1015) );
  AOI22X1 U1500 ( .A(n706), .B(\mem<10><5> ), .C(n707), .D(\mem<8><5> ), .Y(
        n1013) );
  AOI22X1 U1501 ( .A(n708), .B(\mem<14><5> ), .C(n709), .D(\mem<12><5> ), .Y(
        n1012) );
  AOI22X1 U1504 ( .A(n715), .B(\mem<18><5> ), .C(n716), .D(\mem<16><5> ), .Y(
        n1021) );
  AOI22X1 U1505 ( .A(n717), .B(\mem<22><5> ), .C(n718), .D(\mem<20><5> ), .Y(
        n1020) );
  AOI22X1 U1506 ( .A(n719), .B(\mem<26><5> ), .C(n720), .D(\mem<24><5> ), .Y(
        n1018) );
  AOI22X1 U1507 ( .A(n721), .B(\mem<30><5> ), .C(n722), .D(\mem<28><5> ), .Y(
        n1017) );
  OAI21X1 U1508 ( .A(n1022), .B(n2448), .C(n957), .Y(\DataOut<12> ) );
  NOR3X1 U1510 ( .A(n1024), .B(n635), .C(n782), .Y(n1022) );
  AOI22X1 U1513 ( .A(n674), .B(\mem<34><4> ), .C(n675), .D(\mem<32><4> ), .Y(
        n1031) );
  AOI22X1 U1514 ( .A(n676), .B(\mem<38><4> ), .C(n677), .D(\mem<36><4> ), .Y(
        n1030) );
  AOI22X1 U1515 ( .A(n678), .B(\mem<42><4> ), .C(n679), .D(\mem<40><4> ), .Y(
        n1028) );
  AOI22X1 U1516 ( .A(n680), .B(\mem<46><4> ), .C(n681), .D(\mem<44><4> ), .Y(
        n1027) );
  AOI22X1 U1519 ( .A(n687), .B(\mem<58><4> ), .C(n688), .D(\mem<56><4> ), .Y(
        n1036) );
  AOI22X1 U1520 ( .A(n689), .B(\mem<62><4> ), .C(n690), .D(\mem<60><4> ), .Y(
        n1035) );
  AOI22X1 U1521 ( .A(n691), .B(\mem<50><4> ), .C(n692), .D(\mem<48><4> ), .Y(
        n1033) );
  AOI22X1 U1522 ( .A(n693), .B(\mem<54><4> ), .C(n694), .D(\mem<52><4> ), .Y(
        n1032) );
  AOI22X1 U1526 ( .A(n702), .B(\mem<2><4> ), .C(n703), .D(\mem<0><4> ), .Y(
        n1043) );
  AOI22X1 U1527 ( .A(n704), .B(\mem<6><4> ), .C(n705), .D(\mem<4><4> ), .Y(
        n1042) );
  AOI22X1 U1528 ( .A(n706), .B(\mem<10><4> ), .C(n707), .D(\mem<8><4> ), .Y(
        n1040) );
  AOI22X1 U1529 ( .A(n708), .B(\mem<14><4> ), .C(n709), .D(\mem<12><4> ), .Y(
        n1039) );
  AOI22X1 U1532 ( .A(n715), .B(\mem<18><4> ), .C(n716), .D(\mem<16><4> ), .Y(
        n1048) );
  AOI22X1 U1533 ( .A(n717), .B(\mem<22><4> ), .C(n718), .D(\mem<20><4> ), .Y(
        n1047) );
  AOI22X1 U1534 ( .A(n719), .B(\mem<26><4> ), .C(n720), .D(\mem<24><4> ), .Y(
        n1045) );
  AOI22X1 U1535 ( .A(n721), .B(\mem<30><4> ), .C(n722), .D(\mem<28><4> ), .Y(
        n1044) );
  OAI21X1 U1536 ( .A(n1049), .B(n2448), .C(n945), .Y(\DataOut<11> ) );
  NOR3X1 U1538 ( .A(n1051), .B(n631), .C(n768), .Y(n1049) );
  AOI22X1 U1541 ( .A(n674), .B(\mem<34><3> ), .C(n675), .D(\mem<32><3> ), .Y(
        n1058) );
  AOI22X1 U1542 ( .A(n676), .B(\mem<38><3> ), .C(n677), .D(\mem<36><3> ), .Y(
        n1057) );
  AOI22X1 U1543 ( .A(n678), .B(\mem<42><3> ), .C(n679), .D(\mem<40><3> ), .Y(
        n1055) );
  AOI22X1 U1544 ( .A(n680), .B(\mem<46><3> ), .C(n681), .D(\mem<44><3> ), .Y(
        n1054) );
  AOI22X1 U1547 ( .A(n687), .B(\mem<58><3> ), .C(n688), .D(\mem<56><3> ), .Y(
        n1063) );
  AOI22X1 U1548 ( .A(n689), .B(\mem<62><3> ), .C(n690), .D(\mem<60><3> ), .Y(
        n1062) );
  AOI22X1 U1549 ( .A(n691), .B(\mem<50><3> ), .C(n692), .D(\mem<48><3> ), .Y(
        n1060) );
  AOI22X1 U1550 ( .A(n693), .B(\mem<54><3> ), .C(n694), .D(\mem<52><3> ), .Y(
        n1059) );
  AOI22X1 U1554 ( .A(n702), .B(\mem<2><3> ), .C(n703), .D(\mem<0><3> ), .Y(
        n1070) );
  AOI22X1 U1555 ( .A(n704), .B(\mem<6><3> ), .C(n705), .D(\mem<4><3> ), .Y(
        n1069) );
  AOI22X1 U1556 ( .A(n706), .B(\mem<10><3> ), .C(n707), .D(\mem<8><3> ), .Y(
        n1067) );
  AOI22X1 U1557 ( .A(n708), .B(\mem<14><3> ), .C(n709), .D(\mem<12><3> ), .Y(
        n1066) );
  AOI22X1 U1560 ( .A(n715), .B(\mem<18><3> ), .C(n716), .D(\mem<16><3> ), .Y(
        n1075) );
  AOI22X1 U1561 ( .A(n717), .B(\mem<22><3> ), .C(n718), .D(\mem<20><3> ), .Y(
        n1074) );
  AOI22X1 U1562 ( .A(n719), .B(\mem<26><3> ), .C(n720), .D(\mem<24><3> ), .Y(
        n1072) );
  AOI22X1 U1563 ( .A(n721), .B(\mem<30><3> ), .C(n722), .D(\mem<28><3> ), .Y(
        n1071) );
  OAI21X1 U1564 ( .A(n1076), .B(n2448), .C(n942), .Y(\DataOut<10> ) );
  NOR3X1 U1567 ( .A(n1078), .B(n627), .C(n756), .Y(n1076) );
  AOI22X1 U1570 ( .A(n674), .B(\mem<34><2> ), .C(n675), .D(\mem<32><2> ), .Y(
        n1085) );
  AOI22X1 U1573 ( .A(n676), .B(\mem<38><2> ), .C(n677), .D(\mem<36><2> ), .Y(
        n1084) );
  AOI22X1 U1576 ( .A(n678), .B(\mem<42><2> ), .C(n679), .D(\mem<40><2> ), .Y(
        n1082) );
  AOI22X1 U1579 ( .A(n680), .B(\mem<46><2> ), .C(n681), .D(\mem<44><2> ), .Y(
        n1081) );
  AOI22X1 U1584 ( .A(n687), .B(\mem<58><2> ), .C(n688), .D(\mem<56><2> ), .Y(
        n1096) );
  AOI22X1 U1587 ( .A(n689), .B(\mem<62><2> ), .C(n690), .D(\mem<60><2> ), .Y(
        n1095) );
  AOI22X1 U1590 ( .A(n691), .B(\mem<50><2> ), .C(n692), .D(\mem<48><2> ), .Y(
        n1093) );
  AOI22X1 U1593 ( .A(n693), .B(\mem<54><2> ), .C(n694), .D(\mem<52><2> ), .Y(
        n1092) );
  AOI22X1 U1599 ( .A(n702), .B(\mem<2><2> ), .C(n703), .D(\mem<0><2> ), .Y(
        n1105) );
  AOI22X1 U1602 ( .A(n704), .B(\mem<6><2> ), .C(n705), .D(\mem<4><2> ), .Y(
        n1104) );
  AOI22X1 U1605 ( .A(n706), .B(\mem<10><2> ), .C(n707), .D(\mem<8><2> ), .Y(
        n1102) );
  AOI22X1 U1608 ( .A(n708), .B(\mem<14><2> ), .C(n709), .D(\mem<12><2> ), .Y(
        n1101) );
  AOI22X1 U1613 ( .A(n715), .B(\mem<18><2> ), .C(n716), .D(\mem<16><2> ), .Y(
        n1112) );
  AOI22X1 U1616 ( .A(n717), .B(\mem<22><2> ), .C(n718), .D(\mem<20><2> ), .Y(
        n1111) );
  AOI22X1 U1619 ( .A(n719), .B(\mem<26><2> ), .C(n720), .D(\mem<24><2> ), .Y(
        n1109) );
  AOI22X1 U1622 ( .A(n721), .B(\mem<30><2> ), .C(n722), .D(\mem<28><2> ), .Y(
        n1108) );
  OAI21X1 U1625 ( .A(n1115), .B(n2447), .C(n929), .Y(\DataOut<0> ) );
  NAND2X1 U1628 ( .A(err), .B(n2548), .Y(n663) );
  NOR2X1 U1629 ( .A(n2527), .B(n2546), .Y(err) );
  NAND3X1 U1631 ( .A(n2527), .B(n2548), .C(Done), .Y(n751) );
  AOI21X1 U1632 ( .A(n2548), .B(n2547), .C(n2549), .Y(Done) );
  NOR3X1 U1636 ( .A(n1118), .B(n623), .C(n753), .Y(n1115) );
  AOI22X1 U1639 ( .A(\mem<29><0> ), .B(n342), .C(\mem<31><0> ), .D(n324), .Y(
        n1125) );
  AOI22X1 U1642 ( .A(\mem<25><0> ), .B(n378), .C(\mem<27><0> ), .D(n360), .Y(
        n1124) );
  NOR3X1 U1645 ( .A(n2529), .B(N258), .C(n2530), .Y(n1114) );
  AOI22X1 U1646 ( .A(\mem<21><0> ), .B(n414), .C(\mem<23><0> ), .D(n396), .Y(
        n1122) );
  AOI22X1 U1649 ( .A(\mem<17><0> ), .B(n450), .C(\mem<19><0> ), .D(n432), .Y(
        n1121) );
  NOR3X1 U1652 ( .A(N256), .B(N258), .C(n2530), .Y(n1113) );
  AOI22X1 U1655 ( .A(\mem<13><0> ), .B(n486), .C(\mem<15><0> ), .D(n468), .Y(
        n1136) );
  AOI22X1 U1658 ( .A(\mem<9><0> ), .B(n522), .C(\mem<11><0> ), .D(n504), .Y(
        n1135) );
  NOR3X1 U1661 ( .A(N257), .B(N258), .C(n2529), .Y(n1107) );
  AOI22X1 U1662 ( .A(\mem<5><0> ), .B(n558), .C(\mem<7><0> ), .D(n540), .Y(
        n1133) );
  AOI22X1 U1665 ( .A(\mem<1><0> ), .B(n594), .C(\mem<3><0> ), .D(n576), .Y(
        n1132) );
  NOR3X1 U1668 ( .A(N257), .B(N258), .C(N256), .Y(n1106) );
  AOI22X1 U1672 ( .A(\mem<61><0> ), .B(n54), .C(\mem<63><0> ), .D(n35), .Y(
        n1143) );
  AOI22X1 U1675 ( .A(\mem<57><0> ), .B(n90), .C(\mem<59><0> ), .D(n72), .Y(
        n1142) );
  NOR3X1 U1678 ( .A(n2530), .B(n2529), .C(n2543), .Y(n1097) );
  AOI22X1 U1679 ( .A(\mem<53><0> ), .B(n126), .C(\mem<55><0> ), .D(n108), .Y(
        n1140) );
  AOI22X1 U1682 ( .A(\mem<49><0> ), .B(n162), .C(\mem<51><0> ), .D(n144), .Y(
        n1139) );
  NOR3X1 U1685 ( .A(n2530), .B(N256), .C(n2543), .Y(n1098) );
  AOI22X1 U1689 ( .A(\mem<45><0> ), .B(n198), .C(\mem<47><0> ), .D(n180), .Y(
        n1149) );
  AOI22X1 U1692 ( .A(\mem<41><0> ), .B(n234), .C(\mem<43><0> ), .D(n216), .Y(
        n1148) );
  NOR3X1 U1695 ( .A(n2529), .B(N257), .C(n2543), .Y(n1091) );
  AOI22X1 U1697 ( .A(\mem<37><0> ), .B(n270), .C(\mem<39><0> ), .D(n252), .Y(
        n1146) );
  NAND3X1 U1700 ( .A(n2544), .B(n2527), .C(n1090), .Y(n1150) );
  NAND3X1 U1704 ( .A(n2544), .B(n2527), .C(n1089), .Y(n1152) );
  AOI22X1 U1706 ( .A(\mem<33><0> ), .B(n306), .C(\mem<35><0> ), .D(n288), .Y(
        n1145) );
  NAND3X1 U1709 ( .A(n2544), .B(n2527), .C(n2446), .Y(n1154) );
  NOR2X1 U1710 ( .A(n2528), .B(N255), .Y(n1088) );
  NAND3X1 U1714 ( .A(n2544), .B(n2527), .C(n2445), .Y(n1155) );
  NOR2X1 U1715 ( .A(N254), .B(N255), .Y(n1087) );
  NAND3X1 U1718 ( .A(n1157), .B(n1158), .C(n1159), .Y(n1156) );
  NOR3X1 U1719 ( .A(n2545), .B(\Addr<6> ), .C(\Addr<15> ), .Y(n1159) );
  NOR3X1 U1721 ( .A(\Addr<7> ), .B(\Addr<9> ), .C(\Addr<8> ), .Y(n1161) );
  NOR3X1 U1722 ( .A(\Addr<12> ), .B(\Addr<14> ), .C(\Addr<13> ), .Y(n1158) );
  NOR2X1 U1723 ( .A(\Addr<11> ), .B(\Addr<10> ), .Y(n1157) );
  NOR3X1 U1724 ( .A(N256), .B(N257), .C(n2543), .Y(n1086) );
  AND2X2 U1176 ( .A(n672), .B(n673), .Y(n671) );
  AND2X2 U1182 ( .A(n685), .B(n686), .Y(n684) );
  AND2X2 U1189 ( .A(n700), .B(n701), .Y(n699) );
  AND2X2 U1195 ( .A(n713), .B(n714), .Y(n712) );
  AND2X2 U1204 ( .A(n731), .B(n732), .Y(n730) );
  AND2X2 U1210 ( .A(n736), .B(n737), .Y(n735) );
  AND2X2 U1217 ( .A(n743), .B(n744), .Y(n742) );
  AND2X2 U1223 ( .A(n748), .B(n749), .Y(n747) );
  AND2X2 U1232 ( .A(n760), .B(n761), .Y(n759) );
  AND2X2 U1238 ( .A(n765), .B(n766), .Y(n764) );
  AND2X2 U1245 ( .A(n772), .B(n773), .Y(n771) );
  AND2X2 U1251 ( .A(n777), .B(n778), .Y(n776) );
  AND2X2 U1260 ( .A(n787), .B(n788), .Y(n786) );
  AND2X2 U1266 ( .A(n792), .B(n793), .Y(n791) );
  AND2X2 U1273 ( .A(n799), .B(n800), .Y(n798) );
  AND2X2 U1279 ( .A(n804), .B(n805), .Y(n803) );
  AND2X2 U1288 ( .A(n814), .B(n815), .Y(n813) );
  AND2X2 U1294 ( .A(n819), .B(n820), .Y(n818) );
  AND2X2 U1301 ( .A(n826), .B(n827), .Y(n825) );
  AND2X2 U1307 ( .A(n831), .B(n832), .Y(n830) );
  AND2X2 U1316 ( .A(n841), .B(n842), .Y(n840) );
  AND2X2 U1322 ( .A(n846), .B(n847), .Y(n845) );
  AND2X2 U1329 ( .A(n853), .B(n854), .Y(n852) );
  AND2X2 U1335 ( .A(n858), .B(n859), .Y(n857) );
  AND2X2 U1344 ( .A(n868), .B(n869), .Y(n867) );
  AND2X2 U1350 ( .A(n873), .B(n874), .Y(n872) );
  AND2X2 U1357 ( .A(n880), .B(n881), .Y(n879) );
  AND2X2 U1363 ( .A(n885), .B(n886), .Y(n884) );
  AND2X2 U1372 ( .A(n895), .B(n896), .Y(n894) );
  AND2X2 U1378 ( .A(n900), .B(n901), .Y(n899) );
  AND2X2 U1385 ( .A(n907), .B(n908), .Y(n906) );
  AND2X2 U1391 ( .A(n912), .B(n913), .Y(n911) );
  AND2X2 U1400 ( .A(n922), .B(n923), .Y(n921) );
  AND2X2 U1406 ( .A(n927), .B(n928), .Y(n926) );
  AND2X2 U1413 ( .A(n934), .B(n935), .Y(n933) );
  AND2X2 U1419 ( .A(n939), .B(n940), .Y(n938) );
  AND2X2 U1428 ( .A(n949), .B(n950), .Y(n948) );
  AND2X2 U1434 ( .A(n954), .B(n955), .Y(n953) );
  AND2X2 U1441 ( .A(n961), .B(n962), .Y(n960) );
  AND2X2 U1447 ( .A(n966), .B(n967), .Y(n965) );
  AND2X2 U1456 ( .A(n976), .B(n977), .Y(n975) );
  AND2X2 U1462 ( .A(n981), .B(n982), .Y(n980) );
  AND2X2 U1469 ( .A(n988), .B(n989), .Y(n987) );
  AND2X2 U1475 ( .A(n993), .B(n994), .Y(n992) );
  AND2X2 U1484 ( .A(n1003), .B(n1004), .Y(n1002) );
  AND2X2 U1490 ( .A(n1008), .B(n1009), .Y(n1007) );
  AND2X2 U1497 ( .A(n1015), .B(n1016), .Y(n1014) );
  AND2X2 U1503 ( .A(n1020), .B(n1021), .Y(n1019) );
  AND2X2 U1512 ( .A(n1030), .B(n1031), .Y(n1029) );
  AND2X2 U1518 ( .A(n1035), .B(n1036), .Y(n1034) );
  AND2X2 U1525 ( .A(n1042), .B(n1043), .Y(n1041) );
  AND2X2 U1531 ( .A(n1047), .B(n1048), .Y(n1046) );
  AND2X2 U1540 ( .A(n1057), .B(n1058), .Y(n1056) );
  AND2X2 U1546 ( .A(n1062), .B(n1063), .Y(n1061) );
  AND2X2 U1553 ( .A(n1069), .B(n1070), .Y(n1068) );
  AND2X2 U1559 ( .A(n1074), .B(n1075), .Y(n1073) );
  AND2X2 U1569 ( .A(n1084), .B(n1085), .Y(n1083) );
  AND2X2 U1583 ( .A(n1095), .B(n1096), .Y(n1094) );
  AND2X2 U1598 ( .A(n1104), .B(n1105), .Y(n1103) );
  AND2X2 U1612 ( .A(n1111), .B(n1112), .Y(n1110) );
  AND2X2 U1638 ( .A(n1124), .B(n1125), .Y(n1123) );
  AND2X2 U1654 ( .A(n1135), .B(n1136), .Y(n1134) );
  AND2X2 U1671 ( .A(n1142), .B(n1143), .Y(n1141) );
  AND2X2 U1688 ( .A(n1148), .B(n1149), .Y(n1147) );
  INVX1 U35 ( .A(n2536), .Y(n2533) );
  AND2X1 U68 ( .A(n1107), .B(n1090), .Y(n708) );
  AND2X1 U101 ( .A(n1107), .B(n1089), .Y(n709) );
  INVX1 U134 ( .A(Rd), .Y(n2547) );
  INVX1 U167 ( .A(\rand_pat<2> ), .Y(n2579) );
  INVX1 U200 ( .A(n2426), .Y(n2427) );
  INVX1 U233 ( .A(n2425), .Y(n2428) );
  INVX1 U266 ( .A(n2424), .Y(n2431) );
  INVX1 U299 ( .A(n2424), .Y(n2433) );
  AND2X1 U332 ( .A(n1113), .B(n1090), .Y(n717) );
  AND2X1 U365 ( .A(n1113), .B(n1089), .Y(n718) );
  AND2X1 U398 ( .A(n1113), .B(n2446), .Y(n715) );
  AND2X1 U431 ( .A(n1113), .B(n2445), .Y(n716) );
  AND2X1 U464 ( .A(n1114), .B(n2446), .Y(n719) );
  AND2X1 U497 ( .A(n1114), .B(n2445), .Y(n720) );
  AND2X1 U530 ( .A(n1106), .B(n1090), .Y(n704) );
  AND2X1 U563 ( .A(n1106), .B(n1089), .Y(n705) );
  AND2X1 U596 ( .A(n1106), .B(n2446), .Y(n702) );
  AND2X1 U629 ( .A(n1106), .B(n2445), .Y(n703) );
  AND2X1 U662 ( .A(n1107), .B(n2446), .Y(n706) );
  AND2X1 U695 ( .A(n1107), .B(n2445), .Y(n707) );
  INVX1 U728 ( .A(N258), .Y(n2543) );
  INVX1 U761 ( .A(n1161), .Y(n2545) );
  INVX1 U794 ( .A(n2423), .Y(n2440) );
  INVX1 U827 ( .A(n2425), .Y(n2429) );
  INVX1 U860 ( .A(n2425), .Y(n2430) );
  INVX1 U893 ( .A(n2424), .Y(n2432) );
  INVX1 U926 ( .A(n2424), .Y(n2442) );
  INVX1 U959 ( .A(n2425), .Y(n2444) );
  INVX1 U992 ( .A(n2426), .Y(n2437) );
  AND2X1 U1025 ( .A(n1086), .B(n1090), .Y(n676) );
  AND2X1 U1028 ( .A(n1086), .B(n1089), .Y(n677) );
  AND2X1 U1031 ( .A(n1086), .B(n2446), .Y(n674) );
  AND2X1 U1034 ( .A(n1086), .B(n2445), .Y(n675) );
  AND2X1 U1037 ( .A(n1091), .B(n2446), .Y(n678) );
  AND2X1 U1040 ( .A(n1091), .B(n2445), .Y(n679) );
  AND2X1 U1043 ( .A(n1114), .B(n1090), .Y(n721) );
  AND2X1 U1046 ( .A(n1114), .B(n1089), .Y(n722) );
  AND2X1 U1049 ( .A(n2446), .B(n1097), .Y(n687) );
  AND2X1 U1052 ( .A(n2445), .B(n1097), .Y(n688) );
  AND2X1 U1055 ( .A(n1097), .B(n1090), .Y(n689) );
  AND2X1 U1058 ( .A(n1089), .B(n1097), .Y(n690) );
  AND2X1 U1061 ( .A(n1098), .B(n2446), .Y(n691) );
  AND2X1 U1064 ( .A(n1098), .B(n2445), .Y(n692) );
  AND2X1 U1067 ( .A(N255), .B(N254), .Y(n1090) );
  AND2X1 U1070 ( .A(N255), .B(n2528), .Y(n1089) );
  AND2X1 U1073 ( .A(n1091), .B(n1090), .Y(n680) );
  AND2X1 U1075 ( .A(n1091), .B(n1089), .Y(n681) );
  INVX1 U1078 ( .A(n2447), .Y(n2538) );
  AND2X1 U1081 ( .A(n1098), .B(n1090), .Y(n693) );
  AND2X1 U1084 ( .A(n1098), .B(n1089), .Y(n694) );
  OR2X1 U1087 ( .A(n1), .B(n289), .Y(n1118) );
  OR2X1 U1090 ( .A(n27), .B(n541), .Y(n916) );
  OR2X1 U1093 ( .A(n31), .B(n577), .Y(n889) );
  OR2X1 U1096 ( .A(n37), .B(n596), .Y(n862) );
  OR2X1 U1099 ( .A(n73), .B(n599), .Y(n835) );
  OR2X1 U1102 ( .A(n109), .B(n603), .Y(n808) );
  OR2X1 U1105 ( .A(n145), .B(n607), .Y(n781) );
  INVX1 U1108 ( .A(n2448), .Y(n2537) );
  OR2X1 U1111 ( .A(n181), .B(n611), .Y(n754) );
  OR2X1 U1114 ( .A(n217), .B(n615), .Y(n725) );
  OR2X1 U1117 ( .A(n253), .B(n619), .Y(n666) );
  OR2X1 U1120 ( .A(n3), .B(n325), .Y(n1078) );
  OR2X1 U1123 ( .A(n7), .B(n361), .Y(n1051) );
  OR2X1 U1126 ( .A(n11), .B(n397), .Y(n1024) );
  OR2X1 U1129 ( .A(n15), .B(n433), .Y(n997) );
  OR2X1 U1132 ( .A(n19), .B(n469), .Y(n970) );
  OR2X1 U1135 ( .A(n23), .B(n505), .Y(n943) );
  INVX1 U1138 ( .A(\rand_pat<0> ), .Y(n2549) );
  INVX1 U1141 ( .A(\rand_pat<3> ), .Y(n2578) );
  INVX1 U1144 ( .A(\rand_pat<4> ), .Y(n2577) );
  INVX1 U1147 ( .A(\rand_pat<5> ), .Y(n2576) );
  INVX1 U1150 ( .A(\rand_pat<6> ), .Y(n2575) );
  INVX1 U1153 ( .A(\rand_pat<7> ), .Y(n2574) );
  INVX1 U1156 ( .A(\rand_pat<8> ), .Y(n2573) );
  INVX1 U1159 ( .A(\rand_pat<9> ), .Y(n2572) );
  INVX1 U1162 ( .A(\rand_pat<10> ), .Y(n2571) );
  INVX1 U1165 ( .A(\rand_pat<11> ), .Y(n2570) );
  INVX1 U1170 ( .A(\rand_pat<12> ), .Y(n2569) );
  INVX1 U1173 ( .A(\rand_pat<13> ), .Y(n2568) );
  INVX1 U1175 ( .A(\rand_pat<14> ), .Y(n2567) );
  INVX1 U1181 ( .A(\rand_pat<15> ), .Y(n2566) );
  INVX1 U1187 ( .A(\rand_pat<16> ), .Y(n2565) );
  INVX1 U1188 ( .A(\rand_pat<17> ), .Y(n2564) );
  INVX1 U1194 ( .A(\rand_pat<18> ), .Y(n2563) );
  INVX1 U1201 ( .A(\rand_pat<19> ), .Y(n2562) );
  INVX1 U1203 ( .A(\rand_pat<20> ), .Y(n2561) );
  INVX1 U1209 ( .A(\rand_pat<21> ), .Y(n2560) );
  INVX1 U1215 ( .A(\rand_pat<22> ), .Y(n2559) );
  INVX1 U1216 ( .A(\rand_pat<23> ), .Y(n2558) );
  INVX1 U1222 ( .A(\rand_pat<24> ), .Y(n2557) );
  INVX1 U1229 ( .A(\rand_pat<25> ), .Y(n2556) );
  INVX1 U1231 ( .A(\rand_pat<26> ), .Y(n2555) );
  INVX1 U1237 ( .A(\rand_pat<27> ), .Y(n2554) );
  INVX1 U1243 ( .A(\rand_pat<28> ), .Y(n2553) );
  INVX1 U1244 ( .A(\rand_pat<29> ), .Y(n2552) );
  INVX1 U1250 ( .A(\rand_pat<30> ), .Y(n2551) );
  INVX1 U1257 ( .A(\rand_pat<31> ), .Y(n2550) );
  INVX1 U1259 ( .A(\rand_pat<1> ), .Y(n2580) );
  INVX1 U1265 ( .A(n2423), .Y(n2443) );
  INVX1 U1271 ( .A(n2423), .Y(n2441) );
  INVX1 U1272 ( .A(n2423), .Y(n2439) );
  INVX1 U1278 ( .A(n2528), .Y(n2419) );
  INVX1 U1285 ( .A(n2528), .Y(n2418) );
  INVX2 U1287 ( .A(n2527), .Y(n2435) );
  INVX1 U1293 ( .A(n2528), .Y(n2422) );
  INVX1 U1299 ( .A(n2528), .Y(n2420) );
  INVX1 U1300 ( .A(n2528), .Y(n2421) );
  INVX1 U1306 ( .A(n2532), .Y(Stall) );
  INVX1 U1313 ( .A(n2527), .Y(n2526) );
  INVX1 U1315 ( .A(n2412), .Y(n2414) );
  INVX1 U1321 ( .A(n2412), .Y(n2415) );
  INVX1 U1327 ( .A(N254), .Y(n2528) );
  INVX1 U1328 ( .A(n2528), .Y(n2416) );
  INVX1 U1334 ( .A(n2528), .Y(n2417) );
  INVX1 U1341 ( .A(n2423), .Y(n2438) );
  INVX1 U1343 ( .A(n2423), .Y(n2436) );
  INVX1 U1349 ( .A(n2423), .Y(n2434) );
  INVX2 U1355 ( .A(n1881), .Y(n2465) );
  INVX2 U1356 ( .A(n1882), .Y(n2466) );
  INVX2 U1362 ( .A(n1883), .Y(n2467) );
  INVX2 U1369 ( .A(n1884), .Y(n2468) );
  INVX2 U1371 ( .A(n1885), .Y(n2469) );
  INVX2 U1377 ( .A(n1886), .Y(n2470) );
  INVX1 U1383 ( .A(N256), .Y(n2529) );
  INVX1 U1384 ( .A(N255), .Y(n2412) );
  INVX1 U1390 ( .A(n2526), .Y(n2425) );
  INVX1 U1397 ( .A(n2526), .Y(n2424) );
  INVX1 U1399 ( .A(N253), .Y(n2423) );
  INVX1 U1405 ( .A(N257), .Y(n2530) );
  INVX1 U1411 ( .A(n2536), .Y(n2534) );
  INVX1 U1412 ( .A(n36), .Y(n2523) );
  INVX1 U1418 ( .A(n2523), .Y(n2521) );
  INVX1 U1425 ( .A(n2523), .Y(n2522) );
  INVX1 U1427 ( .A(n2529), .Y(n2411) );
  INVX1 U1433 ( .A(n2529), .Y(n2410) );
  INVX1 U1439 ( .A(n2412), .Y(n2413) );
  INVX1 U1440 ( .A(rst), .Y(n2536) );
  INVX1 U1446 ( .A(n2526), .Y(n2426) );
  INVX1 U1453 ( .A(\DataIn<15> ), .Y(n2464) );
  INVX1 U1455 ( .A(\DataIn<14> ), .Y(n2463) );
  INVX1 U1461 ( .A(\DataIn<13> ), .Y(n2462) );
  INVX1 U1467 ( .A(\DataIn<12> ), .Y(n2461) );
  INVX1 U1468 ( .A(\DataIn<11> ), .Y(n2460) );
  INVX1 U1474 ( .A(\DataIn<10> ), .Y(n2459) );
  INVX1 U1481 ( .A(\DataIn<9> ), .Y(n2458) );
  INVX1 U1483 ( .A(\DataIn<8> ), .Y(n2457) );
  INVX1 U1489 ( .A(\DataIn<7> ), .Y(n2456) );
  INVX1 U1495 ( .A(\DataIn<6> ), .Y(n2455) );
  INVX1 U1496 ( .A(\DataIn<5> ), .Y(n2454) );
  INVX1 U1502 ( .A(\DataIn<4> ), .Y(n2453) );
  INVX1 U1509 ( .A(\DataIn<3> ), .Y(n2452) );
  INVX1 U1511 ( .A(\DataIn<2> ), .Y(n2451) );
  INVX1 U1517 ( .A(\DataIn<1> ), .Y(n2450) );
  INVX1 U1523 ( .A(\DataIn<0> ), .Y(n2449) );
  INVX1 U1524 ( .A(n2530), .Y(n2409) );
  BUFX2 U1530 ( .A(n751), .Y(n2447) );
  INVX1 U1537 ( .A(N253), .Y(n2527) );
  BUFX2 U1539 ( .A(n663), .Y(n2448) );
  INVX1 U1545 ( .A(n2581), .Y(n2532) );
  AND2X1 U1551 ( .A(n1113), .B(n2542), .Y(n450) );
  AND2X1 U1552 ( .A(n1106), .B(n2542), .Y(n594) );
  AND2X1 U1558 ( .A(n1086), .B(n2542), .Y(n306) );
  AND2X1 U1565 ( .A(n1098), .B(n2542), .Y(n162) );
  AND2X1 U1566 ( .A(n1114), .B(n2542), .Y(n378) );
  AND2X1 U1568 ( .A(n1107), .B(n2542), .Y(n522) );
  AND2X1 U1571 ( .A(n1091), .B(n2542), .Y(n234) );
  AND2X1 U1572 ( .A(n2542), .B(n1097), .Y(n90) );
  BUFX2 U1574 ( .A(n1087), .Y(n2445) );
  AND2X1 U1575 ( .A(n1113), .B(n2541), .Y(n432) );
  AND2X1 U1577 ( .A(n1106), .B(n2541), .Y(n576) );
  AND2X1 U1578 ( .A(n1086), .B(n2541), .Y(n288) );
  AND2X1 U1580 ( .A(n1098), .B(n2541), .Y(n144) );
  AND2X1 U1581 ( .A(n1114), .B(n2541), .Y(n360) );
  AND2X1 U1582 ( .A(n1107), .B(n2541), .Y(n504) );
  AND2X1 U1585 ( .A(n1091), .B(n2541), .Y(n216) );
  AND2X1 U1586 ( .A(n2541), .B(n1097), .Y(n72) );
  BUFX2 U1588 ( .A(n1088), .Y(n2446) );
  AND2X1 U1589 ( .A(n1113), .B(n2540), .Y(n414) );
  AND2X1 U1591 ( .A(n1106), .B(n2540), .Y(n558) );
  AND2X1 U1592 ( .A(n1114), .B(n2540), .Y(n342) );
  AND2X1 U1594 ( .A(n1107), .B(n2540), .Y(n486) );
  AND2X1 U1595 ( .A(n1086), .B(n2540), .Y(n270) );
  AND2X1 U1596 ( .A(n1098), .B(n2540), .Y(n126) );
  AND2X1 U1597 ( .A(n1091), .B(n2540), .Y(n198) );
  AND2X1 U1600 ( .A(n2540), .B(n1097), .Y(n54) );
  AND2X1 U1601 ( .A(n1113), .B(n2539), .Y(n396) );
  AND2X1 U1603 ( .A(n1106), .B(n2539), .Y(n540) );
  AND2X1 U1604 ( .A(n1114), .B(n2539), .Y(n324) );
  AND2X1 U1606 ( .A(n1107), .B(n2539), .Y(n468) );
  AND2X1 U1607 ( .A(n1086), .B(n2539), .Y(n252) );
  AND2X1 U1609 ( .A(n1098), .B(n2539), .Y(n108) );
  AND2X1 U1610 ( .A(n1091), .B(n2539), .Y(n180) );
  AND2X1 U1611 ( .A(n1097), .B(n2539), .Y(n35) );
  OR2X1 U1614 ( .A(n1117), .B(n2), .Y(n1) );
  OR2X1 U1615 ( .A(n1100), .B(n1116), .Y(n2) );
  OR2X1 U1617 ( .A(n1126), .B(n5), .Y(n3) );
  OR2X1 U1618 ( .A(n1119), .B(n1120), .Y(n5) );
  OR2X1 U1620 ( .A(n1129), .B(n9), .Y(n7) );
  OR2X1 U1621 ( .A(n1127), .B(n1128), .Y(n9) );
  OR2X1 U1623 ( .A(n1137), .B(n13), .Y(n11) );
  OR2X1 U1624 ( .A(n1130), .B(n1131), .Y(n13) );
  OR2X1 U1626 ( .A(n1151), .B(n17), .Y(n15) );
  OR2X1 U1627 ( .A(n1138), .B(n1144), .Y(n17) );
  OR2X1 U1630 ( .A(n1194), .B(n21), .Y(n19) );
  OR2X1 U1633 ( .A(n1153), .B(n1160), .Y(n21) );
  OR2X1 U1634 ( .A(n1709), .B(n25), .Y(n23) );
  OR2X1 U1635 ( .A(n1195), .B(n1708), .Y(n25) );
  OR2X1 U1637 ( .A(n1712), .B(n29), .Y(n27) );
  OR2X1 U1640 ( .A(n1710), .B(n1711), .Y(n29) );
  OR2X1 U1641 ( .A(n1715), .B(n33), .Y(n31) );
  OR2X1 U1643 ( .A(n1713), .B(n1714), .Y(n33) );
  OR2X1 U1644 ( .A(n1718), .B(n55), .Y(n37) );
  OR2X1 U1647 ( .A(n1716), .B(n1717), .Y(n55) );
  OR2X1 U1648 ( .A(n1721), .B(n91), .Y(n73) );
  OR2X1 U1650 ( .A(n1719), .B(n1720), .Y(n91) );
  OR2X1 U1651 ( .A(n1724), .B(n127), .Y(n109) );
  OR2X1 U1653 ( .A(n1722), .B(n1723), .Y(n127) );
  OR2X1 U1656 ( .A(n1727), .B(n163), .Y(n145) );
  OR2X1 U1657 ( .A(n1725), .B(n1726), .Y(n163) );
  OR2X1 U1659 ( .A(n1730), .B(n199), .Y(n181) );
  OR2X1 U1660 ( .A(n1728), .B(n1729), .Y(n199) );
  OR2X1 U1663 ( .A(n1733), .B(n235), .Y(n217) );
  OR2X1 U1664 ( .A(n1731), .B(n1732), .Y(n235) );
  OR2X1 U1666 ( .A(n1736), .B(n271), .Y(n253) );
  OR2X1 U1667 ( .A(n1734), .B(n1735), .Y(n271) );
  OR2X1 U1669 ( .A(n1739), .B(n307), .Y(n289) );
  OR2X1 U1670 ( .A(n1737), .B(n1738), .Y(n307) );
  OR2X1 U1673 ( .A(n1742), .B(n343), .Y(n325) );
  OR2X1 U1674 ( .A(n1740), .B(n1741), .Y(n343) );
  OR2X1 U1676 ( .A(n1745), .B(n379), .Y(n361) );
  OR2X1 U1677 ( .A(n1743), .B(n1744), .Y(n379) );
  OR2X1 U1680 ( .A(n1748), .B(n415), .Y(n397) );
  OR2X1 U1681 ( .A(n1746), .B(n1747), .Y(n415) );
  OR2X1 U1683 ( .A(n1751), .B(n451), .Y(n433) );
  OR2X1 U1684 ( .A(n1749), .B(n1750), .Y(n451) );
  OR2X1 U1686 ( .A(n1754), .B(n487), .Y(n469) );
  OR2X1 U1687 ( .A(n1752), .B(n1753), .Y(n487) );
  OR2X1 U1690 ( .A(n1757), .B(n523), .Y(n505) );
  OR2X1 U1691 ( .A(n1755), .B(n1756), .Y(n523) );
  OR2X1 U1693 ( .A(n1760), .B(n559), .Y(n541) );
  OR2X1 U1694 ( .A(n1758), .B(n1759), .Y(n559) );
  OR2X1 U1696 ( .A(n1763), .B(n595), .Y(n577) );
  OR2X1 U1698 ( .A(n1761), .B(n1762), .Y(n595) );
  OR2X1 U1699 ( .A(n1766), .B(n597), .Y(n596) );
  OR2X1 U1701 ( .A(n1764), .B(n1765), .Y(n597) );
  OR2X1 U1702 ( .A(n1769), .B(n601), .Y(n599) );
  OR2X1 U1703 ( .A(n1767), .B(n1768), .Y(n601) );
  OR2X1 U1705 ( .A(n1772), .B(n605), .Y(n603) );
  OR2X1 U1707 ( .A(n1770), .B(n1771), .Y(n605) );
  OR2X1 U1708 ( .A(n1775), .B(n609), .Y(n607) );
  OR2X1 U1711 ( .A(n1773), .B(n1774), .Y(n609) );
  OR2X1 U1712 ( .A(n1778), .B(n613), .Y(n611) );
  OR2X1 U1713 ( .A(n1776), .B(n1777), .Y(n613) );
  OR2X1 U1716 ( .A(n1781), .B(n617), .Y(n615) );
  OR2X1 U1717 ( .A(n1779), .B(n1780), .Y(n617) );
  OR2X1 U1720 ( .A(n1784), .B(n621), .Y(n619) );
  OR2X1 U1725 ( .A(n1782), .B(n1783), .Y(n621) );
  OR2X1 U1726 ( .A(n1787), .B(n625), .Y(n623) );
  OR2X1 U1727 ( .A(n1785), .B(n1786), .Y(n625) );
  OR2X1 U1728 ( .A(n1790), .B(n629), .Y(n627) );
  OR2X1 U1729 ( .A(n1788), .B(n1789), .Y(n629) );
  OR2X1 U1730 ( .A(n1793), .B(n633), .Y(n631) );
  OR2X1 U1731 ( .A(n1791), .B(n1792), .Y(n633) );
  OR2X1 U1732 ( .A(n1796), .B(n637), .Y(n635) );
  OR2X1 U1733 ( .A(n1794), .B(n1795), .Y(n637) );
  OR2X1 U1734 ( .A(n1799), .B(n641), .Y(n639) );
  OR2X1 U1735 ( .A(n1797), .B(n1798), .Y(n641) );
  OR2X1 U1736 ( .A(n1802), .B(n645), .Y(n643) );
  OR2X1 U1737 ( .A(n1800), .B(n1801), .Y(n645) );
  OR2X1 U1738 ( .A(n1805), .B(n649), .Y(n647) );
  OR2X1 U1739 ( .A(n1803), .B(n1804), .Y(n649) );
  OR2X1 U1740 ( .A(n1808), .B(n653), .Y(n651) );
  OR2X1 U1741 ( .A(n1806), .B(n1807), .Y(n653) );
  OR2X1 U1742 ( .A(n1811), .B(n657), .Y(n655) );
  OR2X1 U1743 ( .A(n1809), .B(n1810), .Y(n657) );
  OR2X1 U1744 ( .A(n1814), .B(n661), .Y(n659) );
  OR2X1 U1745 ( .A(n1812), .B(n1813), .Y(n661) );
  OR2X1 U1746 ( .A(n1817), .B(n665), .Y(n664) );
  OR2X1 U1747 ( .A(n1815), .B(n1816), .Y(n665) );
  OR2X1 U1748 ( .A(n1820), .B(n668), .Y(n667) );
  OR2X1 U1749 ( .A(n1818), .B(n1819), .Y(n668) );
  OR2X1 U1750 ( .A(n1823), .B(n696), .Y(n695) );
  OR2X1 U1751 ( .A(n1821), .B(n1822), .Y(n696) );
  OR2X1 U1752 ( .A(n1826), .B(n726), .Y(n724) );
  OR2X1 U1753 ( .A(n1824), .B(n1825), .Y(n726) );
  OR2X1 U1754 ( .A(n1829), .B(n738), .Y(n727) );
  OR2X1 U1755 ( .A(n1827), .B(n1828), .Y(n738) );
  OR2X1 U1756 ( .A(n1832), .B(n752), .Y(n739) );
  OR2X1 U1757 ( .A(n1830), .B(n1831), .Y(n752) );
  OR2X1 U1758 ( .A(n1835), .B(n755), .Y(n753) );
  OR2X1 U1759 ( .A(n1833), .B(n1834), .Y(n755) );
  OR2X1 U1760 ( .A(n1838), .B(n767), .Y(n756) );
  OR2X1 U1761 ( .A(n1836), .B(n1837), .Y(n767) );
  OR2X1 U1762 ( .A(n1841), .B(n780), .Y(n768) );
  OR2X1 U1763 ( .A(n1839), .B(n1840), .Y(n780) );
  OR2X1 U1764 ( .A(n1844), .B(n783), .Y(n782) );
  OR2X1 U1765 ( .A(n1842), .B(n1843), .Y(n783) );
  OR2X1 U1766 ( .A(n1847), .B(n795), .Y(n794) );
  OR2X1 U1767 ( .A(n1845), .B(n1846), .Y(n795) );
  OR2X1 U1768 ( .A(n1850), .B(n809), .Y(n807) );
  OR2X1 U1769 ( .A(n1848), .B(n1849), .Y(n809) );
  OR2X1 U1770 ( .A(n1853), .B(n821), .Y(n810) );
  OR2X1 U1771 ( .A(n1851), .B(n1852), .Y(n821) );
  OR2X1 U1772 ( .A(n1856), .B(n834), .Y(n822) );
  OR2X1 U1773 ( .A(n1854), .B(n1855), .Y(n834) );
  OR2X1 U1774 ( .A(n1859), .B(n837), .Y(n836) );
  OR2X1 U1775 ( .A(n1857), .B(n1858), .Y(n837) );
  OR2X1 U1776 ( .A(n1862), .B(n849), .Y(n848) );
  OR2X1 U1777 ( .A(n1860), .B(n1861), .Y(n849) );
  OR2X1 U1778 ( .A(n1865), .B(n863), .Y(n861) );
  OR2X1 U1779 ( .A(n1863), .B(n1864), .Y(n863) );
  OR2X1 U1780 ( .A(n1868), .B(n875), .Y(n864) );
  OR2X1 U1781 ( .A(n1866), .B(n1867), .Y(n875) );
  OR2X1 U1782 ( .A(n1871), .B(n888), .Y(n876) );
  OR2X1 U1783 ( .A(n1869), .B(n1870), .Y(n888) );
  OR2X1 U1784 ( .A(n1874), .B(n891), .Y(n890) );
  OR2X1 U1785 ( .A(n1872), .B(n1873), .Y(n891) );
  OR2X1 U1786 ( .A(n1877), .B(n903), .Y(n902) );
  OR2X1 U1787 ( .A(n1875), .B(n1876), .Y(n903) );
  OR2X1 U1788 ( .A(n1880), .B(n917), .Y(n915) );
  OR2X1 U1789 ( .A(n1878), .B(n1879), .Y(n917) );
  AND2X1 U1790 ( .A(N266), .B(n2537), .Y(n918) );
  INVX1 U1791 ( .A(n918), .Y(n929) );
  AND2X1 U1792 ( .A(N264), .B(n2538), .Y(n930) );
  INVX1 U1793 ( .A(n930), .Y(n942) );
  AND2X1 U1794 ( .A(N263), .B(n2538), .Y(n944) );
  INVX1 U1795 ( .A(n944), .Y(n945) );
  AND2X1 U1796 ( .A(N262), .B(n2538), .Y(n956) );
  INVX1 U1797 ( .A(n956), .Y(n957) );
  AND2X1 U1798 ( .A(N261), .B(n2538), .Y(n969) );
  INVX1 U1799 ( .A(n969), .Y(n971) );
  AND2X1 U1800 ( .A(N260), .B(n2538), .Y(n972) );
  INVX1 U1801 ( .A(n972), .Y(n983) );
  AND2X1 U1802 ( .A(N259), .B(n2538), .Y(n984) );
  INVX1 U1803 ( .A(n984), .Y(n996) );
  AND2X1 U1804 ( .A(N265), .B(n2537), .Y(n998) );
  INVX1 U1805 ( .A(n998), .Y(n999) );
  AND2X1 U1806 ( .A(N264), .B(n2537), .Y(n1010) );
  INVX1 U1807 ( .A(n1010), .Y(n1011) );
  AND2X1 U1808 ( .A(N263), .B(n2537), .Y(n1023) );
  INVX1 U1809 ( .A(n1023), .Y(n1025) );
  AND2X1 U1810 ( .A(N262), .B(n2537), .Y(n1026) );
  INVX1 U1811 ( .A(n1026), .Y(n1037) );
  AND2X1 U1812 ( .A(N261), .B(n2537), .Y(n1038) );
  INVX1 U1813 ( .A(n1038), .Y(n1050) );
  AND2X1 U1814 ( .A(N260), .B(n2537), .Y(n1052) );
  INVX1 U1815 ( .A(n1052), .Y(n1053) );
  AND2X1 U1816 ( .A(N259), .B(n2537), .Y(n1064) );
  INVX1 U1817 ( .A(n1064), .Y(n1065) );
  AND2X1 U1818 ( .A(N266), .B(n2538), .Y(n1077) );
  INVX1 U1819 ( .A(n1077), .Y(n1079) );
  AND2X1 U1820 ( .A(N265), .B(n2538), .Y(n1080) );
  INVX1 U1821 ( .A(n1080), .Y(n1099) );
  INVX1 U1822 ( .A(n2536), .Y(n2535) );
  INVX1 U1823 ( .A(n1887), .Y(n2471) );
  INVX1 U1824 ( .A(n1887), .Y(n2472) );
  INVX1 U1825 ( .A(n1888), .Y(n2473) );
  INVX1 U1826 ( .A(n1888), .Y(n2474) );
  INVX1 U1827 ( .A(n1889), .Y(n2475) );
  INVX1 U1828 ( .A(n1889), .Y(n2476) );
  INVX1 U1829 ( .A(n1890), .Y(n2477) );
  INVX1 U1830 ( .A(n1890), .Y(n2478) );
  INVX1 U1831 ( .A(n1891), .Y(n2479) );
  INVX1 U1832 ( .A(n1891), .Y(n2480) );
  INVX1 U1833 ( .A(n1892), .Y(n2481) );
  INVX1 U1834 ( .A(n1892), .Y(n2482) );
  INVX1 U1835 ( .A(n1893), .Y(n2483) );
  INVX1 U1836 ( .A(n1893), .Y(n2484) );
  INVX1 U1837 ( .A(n1894), .Y(n2485) );
  INVX1 U1838 ( .A(n1894), .Y(n2486) );
  INVX1 U1839 ( .A(n1895), .Y(n2487) );
  INVX1 U1840 ( .A(n1895), .Y(n2488) );
  INVX1 U1841 ( .A(n1896), .Y(n2489) );
  INVX1 U1842 ( .A(n1896), .Y(n2490) );
  INVX1 U1843 ( .A(n1897), .Y(n2491) );
  INVX1 U1844 ( .A(n1897), .Y(n2492) );
  INVX1 U1845 ( .A(n1898), .Y(n2493) );
  INVX1 U1846 ( .A(n1898), .Y(n2494) );
  INVX1 U1847 ( .A(n1899), .Y(n2495) );
  INVX1 U1848 ( .A(n1899), .Y(n2496) );
  INVX1 U1849 ( .A(n1900), .Y(n2497) );
  INVX1 U1850 ( .A(n1900), .Y(n2498) );
  INVX1 U1851 ( .A(n1901), .Y(n2499) );
  INVX1 U1852 ( .A(n1901), .Y(n2500) );
  INVX1 U1853 ( .A(n1902), .Y(n2501) );
  INVX1 U1854 ( .A(n1902), .Y(n2502) );
  INVX1 U1855 ( .A(n1903), .Y(n2503) );
  INVX1 U1856 ( .A(n1903), .Y(n2504) );
  INVX1 U1857 ( .A(n1904), .Y(n2505) );
  INVX1 U1858 ( .A(n1904), .Y(n2506) );
  INVX1 U1859 ( .A(n1905), .Y(n2507) );
  INVX1 U1860 ( .A(n1905), .Y(n2508) );
  INVX1 U1861 ( .A(n1906), .Y(n2509) );
  INVX1 U1862 ( .A(n1906), .Y(n2510) );
  INVX1 U1863 ( .A(n1907), .Y(n2511) );
  INVX1 U1864 ( .A(n1907), .Y(n2512) );
  INVX1 U1865 ( .A(n1908), .Y(n2513) );
  INVX1 U1866 ( .A(n1908), .Y(n2514) );
  INVX1 U1867 ( .A(n1909), .Y(n2515) );
  INVX1 U1868 ( .A(n1909), .Y(n2516) );
  INVX1 U1869 ( .A(n1910), .Y(n2517) );
  INVX1 U1870 ( .A(n1910), .Y(n2518) );
  INVX1 U1871 ( .A(n1911), .Y(n2519) );
  INVX1 U1872 ( .A(n1911), .Y(n2520) );
  INVX1 U1873 ( .A(n1912), .Y(n2524) );
  INVX1 U1874 ( .A(n1912), .Y(n2525) );
  INVX1 U1875 ( .A(n1147), .Y(n1100) );
  INVX1 U1876 ( .A(n1146), .Y(n1116) );
  INVX1 U1877 ( .A(n1145), .Y(n1117) );
  INVX1 U1878 ( .A(n1110), .Y(n1119) );
  INVX1 U1879 ( .A(n1109), .Y(n1120) );
  INVX1 U1880 ( .A(n1108), .Y(n1126) );
  INVX1 U1881 ( .A(n1073), .Y(n1127) );
  INVX1 U1882 ( .A(n1072), .Y(n1128) );
  INVX1 U1883 ( .A(n1071), .Y(n1129) );
  INVX1 U1884 ( .A(n1046), .Y(n1130) );
  INVX1 U1885 ( .A(n1045), .Y(n1131) );
  INVX1 U1886 ( .A(n1044), .Y(n1137) );
  INVX1 U1887 ( .A(n1019), .Y(n1138) );
  INVX1 U1888 ( .A(n1018), .Y(n1144) );
  INVX1 U1889 ( .A(n1017), .Y(n1151) );
  INVX1 U1890 ( .A(n992), .Y(n1153) );
  INVX1 U1891 ( .A(n991), .Y(n1160) );
  INVX1 U1892 ( .A(n990), .Y(n1194) );
  INVX1 U1893 ( .A(n965), .Y(n1195) );
  INVX1 U1894 ( .A(n964), .Y(n1708) );
  INVX1 U1895 ( .A(n963), .Y(n1709) );
  INVX1 U1896 ( .A(n938), .Y(n1710) );
  INVX1 U1897 ( .A(n937), .Y(n1711) );
  INVX1 U1898 ( .A(n936), .Y(n1712) );
  INVX1 U1899 ( .A(n911), .Y(n1713) );
  INVX1 U1900 ( .A(n910), .Y(n1714) );
  INVX1 U1901 ( .A(n909), .Y(n1715) );
  INVX1 U1902 ( .A(n884), .Y(n1716) );
  INVX1 U1903 ( .A(n883), .Y(n1717) );
  INVX1 U1904 ( .A(n882), .Y(n1718) );
  INVX1 U1905 ( .A(n857), .Y(n1719) );
  INVX1 U1906 ( .A(n856), .Y(n1720) );
  INVX1 U1907 ( .A(n855), .Y(n1721) );
  INVX1 U1908 ( .A(n830), .Y(n1722) );
  INVX1 U1909 ( .A(n829), .Y(n1723) );
  INVX1 U1910 ( .A(n828), .Y(n1724) );
  INVX1 U1911 ( .A(n803), .Y(n1725) );
  INVX1 U1912 ( .A(n802), .Y(n1726) );
  INVX1 U1913 ( .A(n801), .Y(n1727) );
  INVX1 U1914 ( .A(n776), .Y(n1728) );
  INVX1 U1915 ( .A(n775), .Y(n1729) );
  INVX1 U1916 ( .A(n774), .Y(n1730) );
  INVX1 U1917 ( .A(n747), .Y(n1731) );
  INVX1 U1918 ( .A(n746), .Y(n1732) );
  INVX1 U1919 ( .A(n745), .Y(n1733) );
  INVX1 U1920 ( .A(n712), .Y(n1734) );
  INVX1 U1921 ( .A(n711), .Y(n1735) );
  INVX1 U1922 ( .A(n710), .Y(n1736) );
  INVX1 U1923 ( .A(n1141), .Y(n1737) );
  INVX1 U1924 ( .A(n1140), .Y(n1738) );
  INVX1 U1925 ( .A(n1139), .Y(n1739) );
  INVX1 U1926 ( .A(n1103), .Y(n1740) );
  INVX1 U1927 ( .A(n1102), .Y(n1741) );
  INVX1 U1928 ( .A(n1101), .Y(n1742) );
  INVX1 U1929 ( .A(n1068), .Y(n1743) );
  INVX1 U1930 ( .A(n1067), .Y(n1744) );
  INVX1 U1931 ( .A(n1066), .Y(n1745) );
  INVX1 U1932 ( .A(n1041), .Y(n1746) );
  INVX1 U1933 ( .A(n1040), .Y(n1747) );
  INVX1 U1934 ( .A(n1039), .Y(n1748) );
  INVX1 U1935 ( .A(n1014), .Y(n1749) );
  INVX1 U1936 ( .A(n1013), .Y(n1750) );
  INVX1 U1937 ( .A(n1012), .Y(n1751) );
  INVX1 U1938 ( .A(n987), .Y(n1752) );
  INVX1 U1939 ( .A(n986), .Y(n1753) );
  INVX1 U1940 ( .A(n985), .Y(n1754) );
  INVX1 U1941 ( .A(n960), .Y(n1755) );
  INVX1 U1942 ( .A(n959), .Y(n1756) );
  INVX1 U1943 ( .A(n958), .Y(n1757) );
  INVX1 U1944 ( .A(n933), .Y(n1758) );
  INVX1 U1945 ( .A(n932), .Y(n1759) );
  INVX1 U1946 ( .A(n931), .Y(n1760) );
  INVX1 U1947 ( .A(n906), .Y(n1761) );
  INVX1 U1948 ( .A(n905), .Y(n1762) );
  INVX1 U1949 ( .A(n904), .Y(n1763) );
  INVX1 U1950 ( .A(n879), .Y(n1764) );
  INVX1 U1951 ( .A(n878), .Y(n1765) );
  INVX1 U1952 ( .A(n877), .Y(n1766) );
  INVX1 U1953 ( .A(n852), .Y(n1767) );
  INVX1 U1954 ( .A(n851), .Y(n1768) );
  INVX1 U1955 ( .A(n850), .Y(n1769) );
  INVX1 U1956 ( .A(n825), .Y(n1770) );
  INVX1 U1957 ( .A(n824), .Y(n1771) );
  INVX1 U1958 ( .A(n823), .Y(n1772) );
  INVX1 U1959 ( .A(n798), .Y(n1773) );
  INVX1 U1960 ( .A(n797), .Y(n1774) );
  INVX1 U1961 ( .A(n796), .Y(n1775) );
  INVX1 U1962 ( .A(n771), .Y(n1776) );
  INVX1 U1963 ( .A(n770), .Y(n1777) );
  INVX1 U1964 ( .A(n769), .Y(n1778) );
  INVX1 U1965 ( .A(n742), .Y(n1779) );
  INVX1 U1966 ( .A(n741), .Y(n1780) );
  INVX1 U1967 ( .A(n740), .Y(n1781) );
  INVX1 U1968 ( .A(n699), .Y(n1782) );
  INVX1 U1969 ( .A(n698), .Y(n1783) );
  INVX1 U1970 ( .A(n697), .Y(n1784) );
  INVX1 U1971 ( .A(n1155), .Y(n2542) );
  INVX1 U1972 ( .A(n1154), .Y(n2541) );
  INVX1 U1973 ( .A(n1152), .Y(n2540) );
  INVX1 U1974 ( .A(n1150), .Y(n2539) );
  INVX1 U1975 ( .A(n1156), .Y(n2544) );
  INVX1 U1976 ( .A(n1134), .Y(n1785) );
  INVX1 U1977 ( .A(n1133), .Y(n1786) );
  INVX1 U1978 ( .A(n1132), .Y(n1787) );
  INVX1 U1979 ( .A(n1094), .Y(n1788) );
  INVX1 U1980 ( .A(n1093), .Y(n1789) );
  INVX1 U1981 ( .A(n1092), .Y(n1790) );
  INVX1 U1982 ( .A(n1061), .Y(n1791) );
  INVX1 U1983 ( .A(n1060), .Y(n1792) );
  INVX1 U1984 ( .A(n1059), .Y(n1793) );
  INVX1 U1985 ( .A(n1034), .Y(n1794) );
  INVX1 U1986 ( .A(n1033), .Y(n1795) );
  INVX1 U1987 ( .A(n1032), .Y(n1796) );
  INVX1 U1988 ( .A(n1007), .Y(n1797) );
  INVX1 U1989 ( .A(n1006), .Y(n1798) );
  INVX1 U1990 ( .A(n1005), .Y(n1799) );
  INVX1 U1991 ( .A(n980), .Y(n1800) );
  INVX1 U1992 ( .A(n979), .Y(n1801) );
  INVX1 U1993 ( .A(n978), .Y(n1802) );
  INVX1 U1994 ( .A(n953), .Y(n1803) );
  INVX1 U1995 ( .A(n952), .Y(n1804) );
  INVX1 U1996 ( .A(n951), .Y(n1805) );
  INVX1 U1997 ( .A(n926), .Y(n1806) );
  INVX1 U1998 ( .A(n925), .Y(n1807) );
  INVX1 U1999 ( .A(n924), .Y(n1808) );
  INVX1 U2000 ( .A(n899), .Y(n1809) );
  INVX1 U2001 ( .A(n898), .Y(n1810) );
  INVX1 U2002 ( .A(n897), .Y(n1811) );
  INVX1 U2003 ( .A(n872), .Y(n1812) );
  INVX1 U2004 ( .A(n871), .Y(n1813) );
  INVX1 U2005 ( .A(n870), .Y(n1814) );
  INVX1 U2006 ( .A(n845), .Y(n1815) );
  INVX1 U2007 ( .A(n844), .Y(n1816) );
  INVX1 U2008 ( .A(n843), .Y(n1817) );
  INVX1 U2009 ( .A(n818), .Y(n1818) );
  INVX1 U2010 ( .A(n817), .Y(n1819) );
  INVX1 U2011 ( .A(n816), .Y(n1820) );
  INVX1 U2012 ( .A(n791), .Y(n1821) );
  INVX1 U2013 ( .A(n790), .Y(n1822) );
  INVX1 U2014 ( .A(n789), .Y(n1823) );
  INVX1 U2015 ( .A(n764), .Y(n1824) );
  INVX1 U2016 ( .A(n763), .Y(n1825) );
  INVX1 U2017 ( .A(n762), .Y(n1826) );
  INVX1 U2018 ( .A(n735), .Y(n1827) );
  INVX1 U2019 ( .A(n734), .Y(n1828) );
  INVX1 U2020 ( .A(n733), .Y(n1829) );
  INVX1 U2021 ( .A(n684), .Y(n1830) );
  INVX1 U2022 ( .A(n683), .Y(n1831) );
  INVX1 U2023 ( .A(n682), .Y(n1832) );
  INVX1 U2024 ( .A(n1123), .Y(n1833) );
  INVX1 U2025 ( .A(n1122), .Y(n1834) );
  INVX1 U2026 ( .A(n1121), .Y(n1835) );
  INVX1 U2027 ( .A(n1083), .Y(n1836) );
  INVX1 U2028 ( .A(n1082), .Y(n1837) );
  INVX1 U2029 ( .A(n1081), .Y(n1838) );
  INVX1 U2030 ( .A(n1056), .Y(n1839) );
  INVX1 U2031 ( .A(n1055), .Y(n1840) );
  INVX1 U2032 ( .A(n1054), .Y(n1841) );
  INVX1 U2033 ( .A(n1029), .Y(n1842) );
  INVX1 U2034 ( .A(n1028), .Y(n1843) );
  INVX1 U2035 ( .A(n1027), .Y(n1844) );
  INVX1 U2036 ( .A(n1002), .Y(n1845) );
  INVX1 U2037 ( .A(n1001), .Y(n1846) );
  INVX1 U2038 ( .A(n1000), .Y(n1847) );
  INVX1 U2039 ( .A(n975), .Y(n1848) );
  INVX1 U2040 ( .A(n974), .Y(n1849) );
  INVX1 U2041 ( .A(n973), .Y(n1850) );
  INVX1 U2042 ( .A(n948), .Y(n1851) );
  INVX1 U2043 ( .A(n947), .Y(n1852) );
  INVX1 U2044 ( .A(n946), .Y(n1853) );
  INVX1 U2045 ( .A(n921), .Y(n1854) );
  INVX1 U2046 ( .A(n920), .Y(n1855) );
  INVX1 U2047 ( .A(n919), .Y(n1856) );
  INVX1 U2048 ( .A(n894), .Y(n1857) );
  INVX1 U2049 ( .A(n893), .Y(n1858) );
  INVX1 U2050 ( .A(n892), .Y(n1859) );
  INVX1 U2051 ( .A(n867), .Y(n1860) );
  INVX1 U2052 ( .A(n866), .Y(n1861) );
  INVX1 U2053 ( .A(n865), .Y(n1862) );
  INVX1 U2054 ( .A(n840), .Y(n1863) );
  INVX1 U2055 ( .A(n839), .Y(n1864) );
  INVX1 U2056 ( .A(n838), .Y(n1865) );
  INVX1 U2057 ( .A(n813), .Y(n1866) );
  INVX1 U2058 ( .A(n812), .Y(n1867) );
  INVX1 U2059 ( .A(n811), .Y(n1868) );
  INVX1 U2060 ( .A(n786), .Y(n1869) );
  INVX1 U2061 ( .A(n785), .Y(n1870) );
  INVX1 U2062 ( .A(n784), .Y(n1871) );
  INVX1 U2063 ( .A(n759), .Y(n1872) );
  INVX1 U2064 ( .A(n758), .Y(n1873) );
  INVX1 U2065 ( .A(n757), .Y(n1874) );
  INVX1 U2066 ( .A(n730), .Y(n1875) );
  INVX1 U2067 ( .A(n729), .Y(n1876) );
  INVX1 U2068 ( .A(n728), .Y(n1877) );
  INVX1 U2069 ( .A(n671), .Y(n1878) );
  INVX1 U2070 ( .A(n670), .Y(n1879) );
  INVX1 U2071 ( .A(n669), .Y(n1880) );
  INVX1 U2072 ( .A(Done), .Y(n2546) );
  AND2X1 U2073 ( .A(n594), .B(n2522), .Y(n1881) );
  AND2X1 U2074 ( .A(n576), .B(n2521), .Y(n1882) );
  AND2X1 U2075 ( .A(n558), .B(n2521), .Y(n1883) );
  AND2X1 U2076 ( .A(n540), .B(n2522), .Y(n1884) );
  AND2X1 U2077 ( .A(n522), .B(n2522), .Y(n1885) );
  AND2X1 U2078 ( .A(n504), .B(n2521), .Y(n1886) );
  AND2X1 U2079 ( .A(n486), .B(n2522), .Y(n1887) );
  AND2X1 U2080 ( .A(n468), .B(n2522), .Y(n1888) );
  AND2X1 U2081 ( .A(n450), .B(n2522), .Y(n1889) );
  AND2X1 U2082 ( .A(n432), .B(n2522), .Y(n1890) );
  AND2X1 U2083 ( .A(n414), .B(n2522), .Y(n1891) );
  AND2X1 U2084 ( .A(n396), .B(n2522), .Y(n1892) );
  AND2X1 U2085 ( .A(n378), .B(n2522), .Y(n1893) );
  AND2X1 U2086 ( .A(n360), .B(n2522), .Y(n1894) );
  AND2X1 U2087 ( .A(n342), .B(n2522), .Y(n1895) );
  AND2X1 U2088 ( .A(n324), .B(n2522), .Y(n1896) );
  AND2X1 U2089 ( .A(n306), .B(n2522), .Y(n1897) );
  AND2X1 U2090 ( .A(n288), .B(n2522), .Y(n1898) );
  AND2X1 U2091 ( .A(n270), .B(n2522), .Y(n1899) );
  AND2X1 U2092 ( .A(n252), .B(n2521), .Y(n1900) );
  AND2X1 U2093 ( .A(n234), .B(n2521), .Y(n1901) );
  AND2X1 U2094 ( .A(n216), .B(n2521), .Y(n1902) );
  AND2X1 U2095 ( .A(n198), .B(n2521), .Y(n1903) );
  AND2X1 U2096 ( .A(n180), .B(n2521), .Y(n1904) );
  AND2X1 U2097 ( .A(n162), .B(n2521), .Y(n1905) );
  AND2X1 U2098 ( .A(n144), .B(n2521), .Y(n1906) );
  AND2X1 U2099 ( .A(n126), .B(n2521), .Y(n1907) );
  AND2X1 U2100 ( .A(n108), .B(n2521), .Y(n1908) );
  AND2X1 U2101 ( .A(n90), .B(n2521), .Y(n1909) );
  AND2X1 U2102 ( .A(n72), .B(n2521), .Y(n1910) );
  AND2X1 U2103 ( .A(n54), .B(n2521), .Y(n1911) );
  AND2X1 U2104 ( .A(n35), .B(n2521), .Y(n1912) );
  MUX2X1 U2105 ( .B(n1914), .A(n1915), .S(n2416), .Y(n1913) );
  MUX2X1 U2106 ( .B(n1917), .A(n1918), .S(n2416), .Y(n1916) );
  MUX2X1 U2107 ( .B(n1920), .A(n1921), .S(n2417), .Y(n1919) );
  MUX2X1 U2108 ( .B(n1923), .A(n1924), .S(n2416), .Y(n1922) );
  MUX2X1 U2109 ( .B(n1926), .A(n1927), .S(n2411), .Y(n1925) );
  MUX2X1 U2110 ( .B(n1929), .A(n1930), .S(n2417), .Y(n1928) );
  MUX2X1 U2111 ( .B(n1932), .A(n1933), .S(n2416), .Y(n1931) );
  MUX2X1 U2112 ( .B(n1935), .A(n1936), .S(n2417), .Y(n1934) );
  MUX2X1 U2113 ( .B(n1938), .A(n1939), .S(n2417), .Y(n1937) );
  MUX2X1 U2114 ( .B(n1941), .A(n1942), .S(n2411), .Y(n1940) );
  MUX2X1 U2115 ( .B(n1944), .A(n1945), .S(n2416), .Y(n1943) );
  MUX2X1 U2116 ( .B(n1947), .A(n1948), .S(n2416), .Y(n1946) );
  MUX2X1 U2117 ( .B(n1950), .A(n1951), .S(n2416), .Y(n1949) );
  MUX2X1 U2118 ( .B(n1953), .A(n1954), .S(n2416), .Y(n1952) );
  MUX2X1 U2119 ( .B(n1956), .A(n1957), .S(n2411), .Y(n1955) );
  MUX2X1 U2120 ( .B(n1959), .A(n1960), .S(n2416), .Y(n1958) );
  MUX2X1 U2121 ( .B(n1962), .A(n1963), .S(n2416), .Y(n1961) );
  MUX2X1 U2122 ( .B(n1965), .A(n1966), .S(n2416), .Y(n1964) );
  MUX2X1 U2123 ( .B(n1968), .A(n1969), .S(n2416), .Y(n1967) );
  MUX2X1 U2124 ( .B(n1971), .A(n1972), .S(n2411), .Y(n1970) );
  MUX2X1 U2125 ( .B(n1973), .A(n1974), .S(N258), .Y(N266) );
  MUX2X1 U2126 ( .B(n1976), .A(n1977), .S(n2416), .Y(n1975) );
  MUX2X1 U2127 ( .B(n1979), .A(n1980), .S(n2416), .Y(n1978) );
  MUX2X1 U2128 ( .B(n1982), .A(n1983), .S(n2416), .Y(n1981) );
  MUX2X1 U2129 ( .B(n1985), .A(n1986), .S(n2416), .Y(n1984) );
  MUX2X1 U2130 ( .B(n1988), .A(n1989), .S(n2411), .Y(n1987) );
  MUX2X1 U2131 ( .B(n1991), .A(n1992), .S(n2417), .Y(n1990) );
  MUX2X1 U2132 ( .B(n1994), .A(n1995), .S(n2417), .Y(n1993) );
  MUX2X1 U2133 ( .B(n1997), .A(n1998), .S(n2417), .Y(n1996) );
  MUX2X1 U2134 ( .B(n2000), .A(n2001), .S(n2417), .Y(n1999) );
  MUX2X1 U2135 ( .B(n2003), .A(n2004), .S(n2411), .Y(n2002) );
  MUX2X1 U2136 ( .B(n2006), .A(n2007), .S(n2417), .Y(n2005) );
  MUX2X1 U2137 ( .B(n2009), .A(n2010), .S(n2417), .Y(n2008) );
  MUX2X1 U2138 ( .B(n2012), .A(n2013), .S(n2417), .Y(n2011) );
  MUX2X1 U2139 ( .B(n2015), .A(n2016), .S(n2417), .Y(n2014) );
  MUX2X1 U2140 ( .B(n2018), .A(n2019), .S(n2411), .Y(n2017) );
  MUX2X1 U2141 ( .B(n2021), .A(n2022), .S(n2417), .Y(n2020) );
  MUX2X1 U2142 ( .B(n2024), .A(n2025), .S(n2417), .Y(n2023) );
  MUX2X1 U2143 ( .B(n2027), .A(n2028), .S(n2417), .Y(n2026) );
  MUX2X1 U2144 ( .B(n2030), .A(n2031), .S(n2417), .Y(n2029) );
  MUX2X1 U2145 ( .B(n2033), .A(n2034), .S(n2411), .Y(n2032) );
  MUX2X1 U2146 ( .B(n2035), .A(n2036), .S(N258), .Y(N265) );
  MUX2X1 U2147 ( .B(n2038), .A(n2039), .S(n2421), .Y(n2037) );
  MUX2X1 U2148 ( .B(n2041), .A(n2042), .S(n2417), .Y(n2040) );
  MUX2X1 U2149 ( .B(n2044), .A(n2045), .S(n2419), .Y(n2043) );
  MUX2X1 U2150 ( .B(n2047), .A(n2048), .S(n2422), .Y(n2046) );
  MUX2X1 U2151 ( .B(n2050), .A(n2051), .S(n2411), .Y(n2049) );
  MUX2X1 U2152 ( .B(n2053), .A(n2054), .S(n2416), .Y(n2052) );
  MUX2X1 U2153 ( .B(n2056), .A(n2057), .S(n2418), .Y(n2055) );
  MUX2X1 U2154 ( .B(n2059), .A(n2060), .S(n2418), .Y(n2058) );
  MUX2X1 U2155 ( .B(n2062), .A(n2063), .S(n2420), .Y(n2061) );
  MUX2X1 U2156 ( .B(n2065), .A(n2066), .S(n2411), .Y(n2064) );
  MUX2X1 U2157 ( .B(n2068), .A(n2069), .S(n2418), .Y(n2067) );
  MUX2X1 U2158 ( .B(n2071), .A(n2072), .S(n2420), .Y(n2070) );
  MUX2X1 U2159 ( .B(n2074), .A(n2075), .S(n2420), .Y(n2073) );
  MUX2X1 U2160 ( .B(n2077), .A(n2078), .S(n2416), .Y(n2076) );
  MUX2X1 U2161 ( .B(n2080), .A(n2081), .S(n2411), .Y(n2079) );
  MUX2X1 U2162 ( .B(n2083), .A(n2084), .S(n2418), .Y(n2082) );
  MUX2X1 U2163 ( .B(n2086), .A(n2087), .S(n2418), .Y(n2085) );
  MUX2X1 U2164 ( .B(n2089), .A(n2090), .S(n2418), .Y(n2088) );
  MUX2X1 U2165 ( .B(n2092), .A(n2093), .S(n2418), .Y(n2091) );
  MUX2X1 U2166 ( .B(n2095), .A(n2096), .S(n2411), .Y(n2094) );
  MUX2X1 U2167 ( .B(n2097), .A(n2098), .S(N258), .Y(N264) );
  MUX2X1 U2168 ( .B(n2100), .A(n2101), .S(n2418), .Y(n2099) );
  MUX2X1 U2169 ( .B(n2103), .A(n2104), .S(n2418), .Y(n2102) );
  MUX2X1 U2170 ( .B(n2106), .A(n2107), .S(n2418), .Y(n2105) );
  MUX2X1 U2171 ( .B(n2109), .A(n2110), .S(n2418), .Y(n2108) );
  MUX2X1 U2172 ( .B(n2112), .A(n2113), .S(n2410), .Y(n2111) );
  MUX2X1 U2173 ( .B(n2115), .A(n2116), .S(n2418), .Y(n2114) );
  MUX2X1 U2174 ( .B(n2118), .A(n2119), .S(n2418), .Y(n2117) );
  MUX2X1 U2175 ( .B(n2121), .A(n2122), .S(n2418), .Y(n2120) );
  MUX2X1 U2176 ( .B(n2124), .A(n2125), .S(n2418), .Y(n2123) );
  MUX2X1 U2177 ( .B(n2127), .A(n2128), .S(n2410), .Y(n2126) );
  MUX2X1 U2178 ( .B(n2130), .A(n2131), .S(n2419), .Y(n2129) );
  MUX2X1 U2179 ( .B(n2133), .A(n2134), .S(n2419), .Y(n2132) );
  MUX2X1 U2180 ( .B(n2136), .A(n2137), .S(n2419), .Y(n2135) );
  MUX2X1 U2181 ( .B(n2139), .A(n2140), .S(n2419), .Y(n2138) );
  MUX2X1 U2182 ( .B(n2142), .A(n2143), .S(n2410), .Y(n2141) );
  MUX2X1 U2183 ( .B(n2145), .A(n2146), .S(n2419), .Y(n2144) );
  MUX2X1 U2184 ( .B(n2148), .A(n2149), .S(n2419), .Y(n2147) );
  MUX2X1 U2185 ( .B(n2151), .A(n2152), .S(n2419), .Y(n2150) );
  MUX2X1 U2186 ( .B(n2154), .A(n2155), .S(n2419), .Y(n2153) );
  MUX2X1 U2187 ( .B(n2157), .A(n2158), .S(n2410), .Y(n2156) );
  MUX2X1 U2188 ( .B(n2159), .A(n2160), .S(N258), .Y(N263) );
  MUX2X1 U2189 ( .B(n2162), .A(n2163), .S(n2419), .Y(n2161) );
  MUX2X1 U2190 ( .B(n2165), .A(n2166), .S(n2419), .Y(n2164) );
  MUX2X1 U2191 ( .B(n2168), .A(n2169), .S(n2419), .Y(n2167) );
  MUX2X1 U2192 ( .B(n2171), .A(n2172), .S(n2419), .Y(n2170) );
  MUX2X1 U2193 ( .B(n2174), .A(n2175), .S(n2410), .Y(n2173) );
  MUX2X1 U2194 ( .B(n2177), .A(n2178), .S(n2420), .Y(n2176) );
  MUX2X1 U2195 ( .B(n2180), .A(n2181), .S(n2420), .Y(n2179) );
  MUX2X1 U2196 ( .B(n2183), .A(n2184), .S(n2420), .Y(n2182) );
  MUX2X1 U2197 ( .B(n2186), .A(n2187), .S(n2420), .Y(n2185) );
  MUX2X1 U2198 ( .B(n2189), .A(n2190), .S(n2410), .Y(n2188) );
  MUX2X1 U2199 ( .B(n2192), .A(n2193), .S(n2420), .Y(n2191) );
  MUX2X1 U2200 ( .B(n2195), .A(n2196), .S(n2420), .Y(n2194) );
  MUX2X1 U2201 ( .B(n2198), .A(n2199), .S(n2420), .Y(n2197) );
  MUX2X1 U2202 ( .B(n2201), .A(n2202), .S(n2420), .Y(n2200) );
  MUX2X1 U2203 ( .B(n2204), .A(n2205), .S(n2410), .Y(n2203) );
  MUX2X1 U2204 ( .B(n2207), .A(n2208), .S(n2420), .Y(n2206) );
  MUX2X1 U2205 ( .B(n2210), .A(n2211), .S(n2420), .Y(n2209) );
  MUX2X1 U2206 ( .B(n2213), .A(n2214), .S(n2420), .Y(n2212) );
  MUX2X1 U2207 ( .B(n2216), .A(n2217), .S(n2420), .Y(n2215) );
  MUX2X1 U2208 ( .B(n2219), .A(n2220), .S(n2410), .Y(n2218) );
  MUX2X1 U2209 ( .B(n2221), .A(n2222), .S(N258), .Y(N262) );
  MUX2X1 U2210 ( .B(n2224), .A(n2225), .S(n2421), .Y(n2223) );
  MUX2X1 U2211 ( .B(n2227), .A(n2228), .S(n2421), .Y(n2226) );
  MUX2X1 U2212 ( .B(n2230), .A(n2231), .S(n2421), .Y(n2229) );
  MUX2X1 U2213 ( .B(n2233), .A(n2234), .S(n2421), .Y(n2232) );
  MUX2X1 U2214 ( .B(n2236), .A(n2237), .S(n2410), .Y(n2235) );
  MUX2X1 U2215 ( .B(n2239), .A(n2240), .S(n2421), .Y(n2238) );
  MUX2X1 U2216 ( .B(n2242), .A(n2243), .S(n2421), .Y(n2241) );
  MUX2X1 U2217 ( .B(n2245), .A(n2246), .S(n2421), .Y(n2244) );
  MUX2X1 U2218 ( .B(n2248), .A(n2249), .S(n2421), .Y(n2247) );
  MUX2X1 U2219 ( .B(n2251), .A(n2252), .S(n2410), .Y(n2250) );
  MUX2X1 U2220 ( .B(n2254), .A(n2255), .S(n2421), .Y(n2253) );
  MUX2X1 U2221 ( .B(n2257), .A(n2258), .S(n2421), .Y(n2256) );
  MUX2X1 U2222 ( .B(n2260), .A(n2261), .S(n2421), .Y(n2259) );
  MUX2X1 U2223 ( .B(n2263), .A(n2264), .S(n2421), .Y(n2262) );
  MUX2X1 U2224 ( .B(n2266), .A(n2267), .S(n2410), .Y(n2265) );
  MUX2X1 U2225 ( .B(n2269), .A(n2270), .S(n2422), .Y(n2268) );
  MUX2X1 U2226 ( .B(n2272), .A(n2273), .S(n2422), .Y(n2271) );
  MUX2X1 U2227 ( .B(n2275), .A(n2276), .S(n2422), .Y(n2274) );
  MUX2X1 U2228 ( .B(n2278), .A(n2279), .S(n2422), .Y(n2277) );
  MUX2X1 U2229 ( .B(n2281), .A(n2282), .S(n2410), .Y(n2280) );
  MUX2X1 U2230 ( .B(n2283), .A(n2284), .S(N258), .Y(N261) );
  MUX2X1 U2231 ( .B(n2286), .A(n2287), .S(n2422), .Y(n2285) );
  MUX2X1 U2232 ( .B(n2289), .A(n2290), .S(n2422), .Y(n2288) );
  MUX2X1 U2233 ( .B(n2292), .A(n2293), .S(n2422), .Y(n2291) );
  MUX2X1 U2234 ( .B(n2295), .A(n2296), .S(n2422), .Y(n2294) );
  MUX2X1 U2235 ( .B(n2298), .A(n2299), .S(n2410), .Y(n2297) );
  MUX2X1 U2236 ( .B(n2301), .A(n2302), .S(n2422), .Y(n2300) );
  MUX2X1 U2237 ( .B(n2304), .A(n2305), .S(n2422), .Y(n2303) );
  MUX2X1 U2238 ( .B(n2307), .A(n2308), .S(n2422), .Y(n2306) );
  MUX2X1 U2239 ( .B(n2310), .A(n2311), .S(n2422), .Y(n2309) );
  MUX2X1 U2240 ( .B(n2313), .A(n2314), .S(n2410), .Y(n2312) );
  MUX2X1 U2241 ( .B(n2316), .A(n2317), .S(n2419), .Y(n2315) );
  MUX2X1 U2242 ( .B(n2319), .A(n2320), .S(n2419), .Y(n2318) );
  MUX2X1 U2243 ( .B(n2322), .A(n2323), .S(n2418), .Y(n2321) );
  MUX2X1 U2244 ( .B(n2325), .A(n2326), .S(n2417), .Y(n2324) );
  MUX2X1 U2245 ( .B(n2328), .A(n2329), .S(n2410), .Y(n2327) );
  MUX2X1 U2246 ( .B(n2331), .A(n2332), .S(n2418), .Y(n2330) );
  MUX2X1 U2247 ( .B(n2334), .A(n2335), .S(n2419), .Y(n2333) );
  MUX2X1 U2248 ( .B(n2337), .A(n2338), .S(n2419), .Y(n2336) );
  MUX2X1 U2249 ( .B(n2340), .A(n2341), .S(n2419), .Y(n2339) );
  MUX2X1 U2250 ( .B(n2343), .A(n2344), .S(n2410), .Y(n2342) );
  MUX2X1 U2251 ( .B(n2345), .A(n2346), .S(N258), .Y(N260) );
  MUX2X1 U2252 ( .B(n2348), .A(n2349), .S(n2418), .Y(n2347) );
  MUX2X1 U2253 ( .B(n2351), .A(n2352), .S(n2418), .Y(n2350) );
  MUX2X1 U2254 ( .B(n2354), .A(n2355), .S(n2422), .Y(n2353) );
  MUX2X1 U2255 ( .B(n2357), .A(n2358), .S(n2421), .Y(n2356) );
  MUX2X1 U2256 ( .B(n2360), .A(n2361), .S(n2411), .Y(n2359) );
  MUX2X1 U2257 ( .B(n2363), .A(n2364), .S(n2422), .Y(n2362) );
  MUX2X1 U2258 ( .B(n2366), .A(n2367), .S(n2422), .Y(n2365) );
  MUX2X1 U2259 ( .B(n2369), .A(n2370), .S(n2420), .Y(n2368) );
  MUX2X1 U2260 ( .B(n2372), .A(n2373), .S(n2420), .Y(n2371) );
  MUX2X1 U2261 ( .B(n2375), .A(n2376), .S(n2411), .Y(n2374) );
  MUX2X1 U2262 ( .B(n2378), .A(n2379), .S(n2422), .Y(n2377) );
  MUX2X1 U2263 ( .B(n2381), .A(n2382), .S(n2421), .Y(n2380) );
  MUX2X1 U2264 ( .B(n2384), .A(n2385), .S(n2421), .Y(n2383) );
  MUX2X1 U2265 ( .B(n2387), .A(n2388), .S(n2421), .Y(n2386) );
  MUX2X1 U2266 ( .B(n2390), .A(n2391), .S(n2411), .Y(n2389) );
  MUX2X1 U2267 ( .B(n2393), .A(n2394), .S(n2422), .Y(n2392) );
  MUX2X1 U2268 ( .B(n2396), .A(n2397), .S(n2421), .Y(n2395) );
  MUX2X1 U2269 ( .B(n2399), .A(n2400), .S(n2420), .Y(n2398) );
  MUX2X1 U2270 ( .B(n2402), .A(n2403), .S(n2420), .Y(n2401) );
  MUX2X1 U2271 ( .B(n2405), .A(n2406), .S(n2411), .Y(n2404) );
  MUX2X1 U2272 ( .B(n2407), .A(n2408), .S(N258), .Y(N259) );
  MUX2X1 U2273 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n2435), .Y(n1915) );
  MUX2X1 U2274 ( .B(\mem<60><0> ), .A(\mem<61><0> ), .S(n2435), .Y(n1914) );
  MUX2X1 U2275 ( .B(\mem<58><0> ), .A(\mem<59><0> ), .S(n2435), .Y(n1918) );
  MUX2X1 U2276 ( .B(\mem<56><0> ), .A(\mem<57><0> ), .S(n2435), .Y(n1917) );
  MUX2X1 U2277 ( .B(n1916), .A(n1913), .S(n2415), .Y(n1927) );
  MUX2X1 U2278 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n2427), .Y(n1921) );
  MUX2X1 U2279 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n2427), .Y(n1920) );
  MUX2X1 U2280 ( .B(\mem<50><0> ), .A(\mem<51><0> ), .S(n2427), .Y(n1924) );
  MUX2X1 U2281 ( .B(\mem<48><0> ), .A(\mem<49><0> ), .S(n2427), .Y(n1923) );
  MUX2X1 U2282 ( .B(n1922), .A(n1919), .S(n2415), .Y(n1926) );
  MUX2X1 U2283 ( .B(\mem<46><0> ), .A(\mem<47><0> ), .S(n2427), .Y(n1930) );
  MUX2X1 U2284 ( .B(\mem<44><0> ), .A(\mem<45><0> ), .S(n2427), .Y(n1929) );
  MUX2X1 U2285 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n2427), .Y(n1933) );
  MUX2X1 U2286 ( .B(\mem<40><0> ), .A(\mem<41><0> ), .S(n2427), .Y(n1932) );
  MUX2X1 U2287 ( .B(n1931), .A(n1928), .S(n2415), .Y(n1942) );
  MUX2X1 U2288 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n2427), .Y(n1936) );
  MUX2X1 U2289 ( .B(\mem<36><0> ), .A(\mem<37><0> ), .S(n2427), .Y(n1935) );
  MUX2X1 U2290 ( .B(\mem<34><0> ), .A(\mem<35><0> ), .S(n2427), .Y(n1939) );
  MUX2X1 U2291 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n2427), .Y(n1938) );
  MUX2X1 U2292 ( .B(n1937), .A(n1934), .S(n2415), .Y(n1941) );
  MUX2X1 U2293 ( .B(n1940), .A(n1925), .S(n2409), .Y(n1974) );
  MUX2X1 U2294 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n2440), .Y(n1945) );
  MUX2X1 U2295 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n2439), .Y(n1944) );
  MUX2X1 U2296 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n2439), .Y(n1948) );
  MUX2X1 U2297 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n2439), .Y(n1947) );
  MUX2X1 U2298 ( .B(n1946), .A(n1943), .S(n2415), .Y(n1957) );
  MUX2X1 U2299 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n2443), .Y(n1951) );
  MUX2X1 U2300 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n2441), .Y(n1950) );
  MUX2X1 U2301 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n2440), .Y(n1954) );
  MUX2X1 U2302 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n2441), .Y(n1953) );
  MUX2X1 U2303 ( .B(n1952), .A(n1949), .S(n2415), .Y(n1956) );
  MUX2X1 U2304 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n2443), .Y(n1960) );
  MUX2X1 U2305 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n2443), .Y(n1959) );
  MUX2X1 U2306 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n2443), .Y(n1963) );
  MUX2X1 U2307 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n2440), .Y(n1962) );
  MUX2X1 U2308 ( .B(n1961), .A(n1958), .S(n2415), .Y(n1972) );
  MUX2X1 U2309 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n2428), .Y(n1966) );
  MUX2X1 U2310 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n2428), .Y(n1965) );
  MUX2X1 U2311 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n2428), .Y(n1969) );
  MUX2X1 U2312 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n2428), .Y(n1968) );
  MUX2X1 U2313 ( .B(n1967), .A(n1964), .S(n2415), .Y(n1971) );
  MUX2X1 U2314 ( .B(n1970), .A(n1955), .S(n2409), .Y(n1973) );
  MUX2X1 U2315 ( .B(\mem<62><1> ), .A(\mem<63><1> ), .S(n2428), .Y(n1977) );
  MUX2X1 U2316 ( .B(\mem<60><1> ), .A(\mem<61><1> ), .S(n2428), .Y(n1976) );
  MUX2X1 U2317 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n2428), .Y(n1980) );
  MUX2X1 U2318 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n2428), .Y(n1979) );
  MUX2X1 U2319 ( .B(n1978), .A(n1975), .S(n2415), .Y(n1989) );
  MUX2X1 U2320 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n2428), .Y(n1983) );
  MUX2X1 U2321 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n2428), .Y(n1982) );
  MUX2X1 U2322 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n2428), .Y(n1986) );
  MUX2X1 U2323 ( .B(\mem<48><1> ), .A(\mem<49><1> ), .S(n2428), .Y(n1985) );
  MUX2X1 U2324 ( .B(n1984), .A(n1981), .S(n2415), .Y(n1988) );
  MUX2X1 U2325 ( .B(\mem<46><1> ), .A(\mem<47><1> ), .S(n2429), .Y(n1992) );
  MUX2X1 U2326 ( .B(\mem<44><1> ), .A(\mem<45><1> ), .S(n2429), .Y(n1991) );
  MUX2X1 U2327 ( .B(\mem<42><1> ), .A(\mem<43><1> ), .S(n2429), .Y(n1995) );
  MUX2X1 U2328 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n2429), .Y(n1994) );
  MUX2X1 U2329 ( .B(n1993), .A(n1990), .S(n2415), .Y(n2004) );
  MUX2X1 U2330 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n2429), .Y(n1998) );
  MUX2X1 U2331 ( .B(\mem<36><1> ), .A(\mem<37><1> ), .S(n2429), .Y(n1997) );
  MUX2X1 U2332 ( .B(\mem<34><1> ), .A(\mem<35><1> ), .S(n2429), .Y(n2001) );
  MUX2X1 U2333 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n2429), .Y(n2000) );
  MUX2X1 U2334 ( .B(n1999), .A(n1996), .S(n2415), .Y(n2003) );
  MUX2X1 U2335 ( .B(n2002), .A(n1987), .S(n2409), .Y(n2036) );
  MUX2X1 U2336 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n2429), .Y(n2007) );
  MUX2X1 U2337 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n2429), .Y(n2006) );
  MUX2X1 U2338 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n2429), .Y(n2010) );
  MUX2X1 U2339 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n2429), .Y(n2009) );
  MUX2X1 U2340 ( .B(n2008), .A(n2005), .S(n2414), .Y(n2019) );
  MUX2X1 U2341 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n2430), .Y(n2013) );
  MUX2X1 U2342 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2430), .Y(n2012) );
  MUX2X1 U2343 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n2430), .Y(n2016) );
  MUX2X1 U2344 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n2430), .Y(n2015) );
  MUX2X1 U2345 ( .B(n2014), .A(n2011), .S(n2414), .Y(n2018) );
  MUX2X1 U2346 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n2430), .Y(n2022) );
  MUX2X1 U2347 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n2430), .Y(n2021) );
  MUX2X1 U2348 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n2430), .Y(n2025) );
  MUX2X1 U2349 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2430), .Y(n2024) );
  MUX2X1 U2350 ( .B(n2023), .A(n2020), .S(n2414), .Y(n2034) );
  MUX2X1 U2351 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n2430), .Y(n2028) );
  MUX2X1 U2352 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n2430), .Y(n2027) );
  MUX2X1 U2353 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n2430), .Y(n2031) );
  MUX2X1 U2354 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n2430), .Y(n2030) );
  MUX2X1 U2355 ( .B(n2029), .A(n2026), .S(n2414), .Y(n2033) );
  MUX2X1 U2356 ( .B(n2032), .A(n2017), .S(n2409), .Y(n2035) );
  MUX2X1 U2357 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n2431), .Y(n2039) );
  MUX2X1 U2358 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n2431), .Y(n2038) );
  MUX2X1 U2359 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n2431), .Y(n2042) );
  MUX2X1 U2360 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n2431), .Y(n2041) );
  MUX2X1 U2361 ( .B(n2040), .A(n2037), .S(n2414), .Y(n2051) );
  MUX2X1 U2362 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n2431), .Y(n2045) );
  MUX2X1 U2363 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n2431), .Y(n2044) );
  MUX2X1 U2364 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n2431), .Y(n2048) );
  MUX2X1 U2365 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n2431), .Y(n2047) );
  MUX2X1 U2366 ( .B(n2046), .A(n2043), .S(n2414), .Y(n2050) );
  MUX2X1 U2367 ( .B(\mem<46><2> ), .A(\mem<47><2> ), .S(n2431), .Y(n2054) );
  MUX2X1 U2368 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n2431), .Y(n2053) );
  MUX2X1 U2369 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n2431), .Y(n2057) );
  MUX2X1 U2370 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n2431), .Y(n2056) );
  MUX2X1 U2371 ( .B(n2055), .A(n2052), .S(n2414), .Y(n2066) );
  MUX2X1 U2372 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n2432), .Y(n2060) );
  MUX2X1 U2373 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n2432), .Y(n2059) );
  MUX2X1 U2374 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n2432), .Y(n2063) );
  MUX2X1 U2375 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n2432), .Y(n2062) );
  MUX2X1 U2376 ( .B(n2061), .A(n2058), .S(n2414), .Y(n2065) );
  MUX2X1 U2377 ( .B(n2064), .A(n2049), .S(n2409), .Y(n2098) );
  MUX2X1 U2378 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2432), .Y(n2069) );
  MUX2X1 U2379 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n2432), .Y(n2068) );
  MUX2X1 U2380 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n2432), .Y(n2072) );
  MUX2X1 U2381 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n2432), .Y(n2071) );
  MUX2X1 U2382 ( .B(n2070), .A(n2067), .S(n2414), .Y(n2081) );
  MUX2X1 U2383 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2432), .Y(n2075) );
  MUX2X1 U2384 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n2432), .Y(n2074) );
  MUX2X1 U2385 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n2432), .Y(n2078) );
  MUX2X1 U2386 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n2432), .Y(n2077) );
  MUX2X1 U2387 ( .B(n2076), .A(n2073), .S(n2414), .Y(n2080) );
  MUX2X1 U2388 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2433), .Y(n2084) );
  MUX2X1 U2389 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n2433), .Y(n2083) );
  MUX2X1 U2390 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n2433), .Y(n2087) );
  MUX2X1 U2391 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n2433), .Y(n2086) );
  MUX2X1 U2392 ( .B(n2085), .A(n2082), .S(n2414), .Y(n2096) );
  MUX2X1 U2393 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n2433), .Y(n2090) );
  MUX2X1 U2394 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n2433), .Y(n2089) );
  MUX2X1 U2395 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n2433), .Y(n2093) );
  MUX2X1 U2396 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2433), .Y(n2092) );
  MUX2X1 U2397 ( .B(n2091), .A(n2088), .S(n2414), .Y(n2095) );
  MUX2X1 U2398 ( .B(n2094), .A(n2079), .S(n2409), .Y(n2097) );
  MUX2X1 U2399 ( .B(\mem<62><3> ), .A(\mem<63><3> ), .S(n2433), .Y(n2101) );
  MUX2X1 U2400 ( .B(\mem<60><3> ), .A(\mem<61><3> ), .S(n2433), .Y(n2100) );
  MUX2X1 U2401 ( .B(\mem<58><3> ), .A(\mem<59><3> ), .S(n2433), .Y(n2104) );
  MUX2X1 U2402 ( .B(\mem<56><3> ), .A(\mem<57><3> ), .S(n2433), .Y(n2103) );
  MUX2X1 U2403 ( .B(n2102), .A(n2099), .S(n2415), .Y(n2113) );
  MUX2X1 U2404 ( .B(\mem<54><3> ), .A(\mem<55><3> ), .S(n2434), .Y(n2107) );
  MUX2X1 U2405 ( .B(\mem<52><3> ), .A(\mem<53><3> ), .S(n2434), .Y(n2106) );
  MUX2X1 U2406 ( .B(\mem<50><3> ), .A(\mem<51><3> ), .S(n2434), .Y(n2110) );
  MUX2X1 U2407 ( .B(\mem<48><3> ), .A(\mem<49><3> ), .S(n2434), .Y(n2109) );
  MUX2X1 U2408 ( .B(n2108), .A(n2105), .S(n2414), .Y(n2112) );
  MUX2X1 U2409 ( .B(\mem<46><3> ), .A(\mem<47><3> ), .S(n2434), .Y(n2116) );
  MUX2X1 U2410 ( .B(\mem<44><3> ), .A(\mem<45><3> ), .S(n2434), .Y(n2115) );
  MUX2X1 U2411 ( .B(\mem<42><3> ), .A(\mem<43><3> ), .S(n2434), .Y(n2119) );
  MUX2X1 U2412 ( .B(\mem<40><3> ), .A(\mem<41><3> ), .S(n2434), .Y(n2118) );
  MUX2X1 U2413 ( .B(n2117), .A(n2114), .S(n2415), .Y(n2128) );
  MUX2X1 U2414 ( .B(\mem<38><3> ), .A(\mem<39><3> ), .S(n2434), .Y(n2122) );
  MUX2X1 U2415 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n2434), .Y(n2121) );
  MUX2X1 U2416 ( .B(\mem<34><3> ), .A(\mem<35><3> ), .S(n2434), .Y(n2125) );
  MUX2X1 U2417 ( .B(\mem<32><3> ), .A(\mem<33><3> ), .S(n2434), .Y(n2124) );
  MUX2X1 U2418 ( .B(n2123), .A(n2120), .S(n2414), .Y(n2127) );
  MUX2X1 U2419 ( .B(n2126), .A(n2111), .S(n2409), .Y(n2160) );
  MUX2X1 U2420 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n2435), .Y(n2131) );
  MUX2X1 U2421 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n2435), .Y(n2130) );
  MUX2X1 U2422 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2435), .Y(n2134) );
  MUX2X1 U2423 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n2435), .Y(n2133) );
  MUX2X1 U2424 ( .B(n2132), .A(n2129), .S(n2414), .Y(n2143) );
  MUX2X1 U2425 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n2435), .Y(n2137) );
  MUX2X1 U2426 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n2435), .Y(n2136) );
  MUX2X1 U2427 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n2435), .Y(n2140) );
  MUX2X1 U2428 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n2435), .Y(n2139) );
  MUX2X1 U2429 ( .B(n2138), .A(n2135), .S(n2415), .Y(n2142) );
  MUX2X1 U2430 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n2435), .Y(n2146) );
  MUX2X1 U2431 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n2435), .Y(n2145) );
  MUX2X1 U2432 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n2435), .Y(n2149) );
  MUX2X1 U2433 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n2435), .Y(n2148) );
  MUX2X1 U2434 ( .B(n2147), .A(n2144), .S(n2414), .Y(n2158) );
  MUX2X1 U2435 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n2435), .Y(n2152) );
  MUX2X1 U2436 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n2435), .Y(n2151) );
  MUX2X1 U2437 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n2435), .Y(n2155) );
  MUX2X1 U2438 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2435), .Y(n2154) );
  MUX2X1 U2439 ( .B(n2153), .A(n2150), .S(n2415), .Y(n2157) );
  MUX2X1 U2440 ( .B(n2156), .A(n2141), .S(n2409), .Y(n2159) );
  MUX2X1 U2441 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n2435), .Y(n2163) );
  MUX2X1 U2442 ( .B(\mem<60><4> ), .A(\mem<61><4> ), .S(n2435), .Y(n2162) );
  MUX2X1 U2443 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n2435), .Y(n2166) );
  MUX2X1 U2444 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n2435), .Y(n2165) );
  MUX2X1 U2445 ( .B(n2164), .A(n2161), .S(n2414), .Y(n2175) );
  MUX2X1 U2446 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n2435), .Y(n2169) );
  MUX2X1 U2447 ( .B(\mem<52><4> ), .A(\mem<53><4> ), .S(n2435), .Y(n2168) );
  MUX2X1 U2448 ( .B(\mem<50><4> ), .A(\mem<51><4> ), .S(n2435), .Y(n2172) );
  MUX2X1 U2449 ( .B(\mem<48><4> ), .A(\mem<49><4> ), .S(n2435), .Y(n2171) );
  MUX2X1 U2450 ( .B(n2170), .A(n2167), .S(n2415), .Y(n2174) );
  MUX2X1 U2451 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n2436), .Y(n2178) );
  MUX2X1 U2452 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n2436), .Y(n2177) );
  MUX2X1 U2453 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n2436), .Y(n2181) );
  MUX2X1 U2454 ( .B(\mem<40><4> ), .A(\mem<41><4> ), .S(n2436), .Y(n2180) );
  MUX2X1 U2455 ( .B(n2179), .A(n2176), .S(n2414), .Y(n2190) );
  MUX2X1 U2456 ( .B(\mem<38><4> ), .A(\mem<39><4> ), .S(n2436), .Y(n2184) );
  MUX2X1 U2457 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n2436), .Y(n2183) );
  MUX2X1 U2458 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n2436), .Y(n2187) );
  MUX2X1 U2459 ( .B(\mem<32><4> ), .A(\mem<33><4> ), .S(n2436), .Y(n2186) );
  MUX2X1 U2460 ( .B(n2185), .A(n2182), .S(n2415), .Y(n2189) );
  MUX2X1 U2461 ( .B(n2188), .A(n2173), .S(n2409), .Y(n2222) );
  MUX2X1 U2462 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n2436), .Y(n2193) );
  MUX2X1 U2463 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n2436), .Y(n2192) );
  MUX2X1 U2464 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n2436), .Y(n2196) );
  MUX2X1 U2465 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n2436), .Y(n2195) );
  MUX2X1 U2466 ( .B(n2194), .A(n2191), .S(n2413), .Y(n2205) );
  MUX2X1 U2467 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n2437), .Y(n2199) );
  MUX2X1 U2468 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2437), .Y(n2198) );
  MUX2X1 U2469 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n2437), .Y(n2202) );
  MUX2X1 U2470 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n2437), .Y(n2201) );
  MUX2X1 U2471 ( .B(n2200), .A(n2197), .S(n2413), .Y(n2204) );
  MUX2X1 U2472 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2437), .Y(n2208) );
  MUX2X1 U2473 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n2437), .Y(n2207) );
  MUX2X1 U2474 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n2437), .Y(n2211) );
  MUX2X1 U2475 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n2437), .Y(n2210) );
  MUX2X1 U2476 ( .B(n2209), .A(n2206), .S(n2413), .Y(n2220) );
  MUX2X1 U2477 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n2437), .Y(n2214) );
  MUX2X1 U2478 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2437), .Y(n2213) );
  MUX2X1 U2479 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n2437), .Y(n2217) );
  MUX2X1 U2480 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n2437), .Y(n2216) );
  MUX2X1 U2481 ( .B(n2215), .A(n2212), .S(n2413), .Y(n2219) );
  MUX2X1 U2482 ( .B(n2218), .A(n2203), .S(n2409), .Y(n2221) );
  MUX2X1 U2483 ( .B(\mem<62><5> ), .A(\mem<63><5> ), .S(n2438), .Y(n2225) );
  MUX2X1 U2484 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n2438), .Y(n2224) );
  MUX2X1 U2485 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n2438), .Y(n2228) );
  MUX2X1 U2486 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n2438), .Y(n2227) );
  MUX2X1 U2487 ( .B(n2226), .A(n2223), .S(n2413), .Y(n2237) );
  MUX2X1 U2488 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n2438), .Y(n2231) );
  MUX2X1 U2489 ( .B(\mem<52><5> ), .A(\mem<53><5> ), .S(n2438), .Y(n2230) );
  MUX2X1 U2490 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n2438), .Y(n2234) );
  MUX2X1 U2491 ( .B(\mem<48><5> ), .A(\mem<49><5> ), .S(n2438), .Y(n2233) );
  MUX2X1 U2492 ( .B(n2232), .A(n2229), .S(n2413), .Y(n2236) );
  MUX2X1 U2493 ( .B(\mem<46><5> ), .A(\mem<47><5> ), .S(n2438), .Y(n2240) );
  MUX2X1 U2494 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n2438), .Y(n2239) );
  MUX2X1 U2495 ( .B(\mem<42><5> ), .A(\mem<43><5> ), .S(n2438), .Y(n2243) );
  MUX2X1 U2496 ( .B(\mem<40><5> ), .A(\mem<41><5> ), .S(n2438), .Y(n2242) );
  MUX2X1 U2497 ( .B(n2241), .A(n2238), .S(n2413), .Y(n2252) );
  MUX2X1 U2498 ( .B(\mem<38><5> ), .A(\mem<39><5> ), .S(n2439), .Y(n2246) );
  MUX2X1 U2499 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n2439), .Y(n2245) );
  MUX2X1 U2500 ( .B(\mem<34><5> ), .A(\mem<35><5> ), .S(n2439), .Y(n2249) );
  MUX2X1 U2501 ( .B(\mem<32><5> ), .A(\mem<33><5> ), .S(n2439), .Y(n2248) );
  MUX2X1 U2502 ( .B(n2247), .A(n2244), .S(n2413), .Y(n2251) );
  MUX2X1 U2503 ( .B(n2250), .A(n2235), .S(n2409), .Y(n2284) );
  MUX2X1 U2504 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n2439), .Y(n2255) );
  MUX2X1 U2505 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n2439), .Y(n2254) );
  MUX2X1 U2506 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n2439), .Y(n2258) );
  MUX2X1 U2507 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n2439), .Y(n2257) );
  MUX2X1 U2508 ( .B(n2256), .A(n2253), .S(n2413), .Y(n2267) );
  MUX2X1 U2509 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n2439), .Y(n2261) );
  MUX2X1 U2510 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n2439), .Y(n2260) );
  MUX2X1 U2511 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n2439), .Y(n2264) );
  MUX2X1 U2512 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n2439), .Y(n2263) );
  MUX2X1 U2513 ( .B(n2262), .A(n2259), .S(n2413), .Y(n2266) );
  MUX2X1 U2514 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n2440), .Y(n2270) );
  MUX2X1 U2515 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n2440), .Y(n2269) );
  MUX2X1 U2516 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n2440), .Y(n2273) );
  MUX2X1 U2517 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n2440), .Y(n2272) );
  MUX2X1 U2518 ( .B(n2271), .A(n2268), .S(n2413), .Y(n2282) );
  MUX2X1 U2519 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n2440), .Y(n2276) );
  MUX2X1 U2520 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n2440), .Y(n2275) );
  MUX2X1 U2521 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n2440), .Y(n2279) );
  MUX2X1 U2522 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n2440), .Y(n2278) );
  MUX2X1 U2523 ( .B(n2277), .A(n2274), .S(n2413), .Y(n2281) );
  MUX2X1 U2524 ( .B(n2280), .A(n2265), .S(n2409), .Y(n2283) );
  MUX2X1 U2525 ( .B(\mem<62><6> ), .A(\mem<63><6> ), .S(n2440), .Y(n2287) );
  MUX2X1 U2526 ( .B(\mem<60><6> ), .A(\mem<61><6> ), .S(n2440), .Y(n2286) );
  MUX2X1 U2527 ( .B(\mem<58><6> ), .A(\mem<59><6> ), .S(n2440), .Y(n2290) );
  MUX2X1 U2528 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n2440), .Y(n2289) );
  MUX2X1 U2529 ( .B(n2288), .A(n2285), .S(n2415), .Y(n2299) );
  MUX2X1 U2530 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n2441), .Y(n2293) );
  MUX2X1 U2531 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n2441), .Y(n2292) );
  MUX2X1 U2532 ( .B(\mem<50><6> ), .A(\mem<51><6> ), .S(n2441), .Y(n2296) );
  MUX2X1 U2533 ( .B(\mem<48><6> ), .A(\mem<49><6> ), .S(n2441), .Y(n2295) );
  MUX2X1 U2534 ( .B(n2294), .A(n2291), .S(n2415), .Y(n2298) );
  MUX2X1 U2535 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n2441), .Y(n2302) );
  MUX2X1 U2536 ( .B(\mem<44><6> ), .A(\mem<45><6> ), .S(n2441), .Y(n2301) );
  MUX2X1 U2537 ( .B(\mem<42><6> ), .A(\mem<43><6> ), .S(n2441), .Y(n2305) );
  MUX2X1 U2538 ( .B(\mem<40><6> ), .A(\mem<41><6> ), .S(n2441), .Y(n2304) );
  MUX2X1 U2539 ( .B(n2303), .A(n2300), .S(n2413), .Y(n2314) );
  MUX2X1 U2540 ( .B(\mem<38><6> ), .A(\mem<39><6> ), .S(n2441), .Y(n2308) );
  MUX2X1 U2541 ( .B(\mem<36><6> ), .A(\mem<37><6> ), .S(n2441), .Y(n2307) );
  MUX2X1 U2542 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n2441), .Y(n2311) );
  MUX2X1 U2543 ( .B(\mem<32><6> ), .A(\mem<33><6> ), .S(n2441), .Y(n2310) );
  MUX2X1 U2544 ( .B(n2309), .A(n2306), .S(n2413), .Y(n2313) );
  MUX2X1 U2545 ( .B(n2312), .A(n2297), .S(n2409), .Y(n2346) );
  MUX2X1 U2546 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n2442), .Y(n2317) );
  MUX2X1 U2547 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n2442), .Y(n2316) );
  MUX2X1 U2548 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n2442), .Y(n2320) );
  MUX2X1 U2549 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n2442), .Y(n2319) );
  MUX2X1 U2550 ( .B(n2318), .A(n2315), .S(n2414), .Y(n2329) );
  MUX2X1 U2551 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n2442), .Y(n2323) );
  MUX2X1 U2552 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n2442), .Y(n2322) );
  MUX2X1 U2553 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n2442), .Y(n2326) );
  MUX2X1 U2554 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n2442), .Y(n2325) );
  MUX2X1 U2555 ( .B(n2324), .A(n2321), .S(n2413), .Y(n2328) );
  MUX2X1 U2556 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n2442), .Y(n2332) );
  MUX2X1 U2557 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n2442), .Y(n2331) );
  MUX2X1 U2558 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n2442), .Y(n2335) );
  MUX2X1 U2559 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n2442), .Y(n2334) );
  MUX2X1 U2560 ( .B(n2333), .A(n2330), .S(n2413), .Y(n2344) );
  MUX2X1 U2561 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n2443), .Y(n2338) );
  MUX2X1 U2562 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n2443), .Y(n2337) );
  MUX2X1 U2563 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n2443), .Y(n2341) );
  MUX2X1 U2564 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n2443), .Y(n2340) );
  MUX2X1 U2565 ( .B(n2339), .A(n2336), .S(n2414), .Y(n2343) );
  MUX2X1 U2566 ( .B(n2342), .A(n2327), .S(n2409), .Y(n2345) );
  MUX2X1 U2567 ( .B(\mem<62><7> ), .A(\mem<63><7> ), .S(n2443), .Y(n2349) );
  MUX2X1 U2568 ( .B(\mem<60><7> ), .A(\mem<61><7> ), .S(n2443), .Y(n2348) );
  MUX2X1 U2569 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n2443), .Y(n2352) );
  MUX2X1 U2570 ( .B(\mem<56><7> ), .A(\mem<57><7> ), .S(n2443), .Y(n2351) );
  MUX2X1 U2571 ( .B(n2350), .A(n2347), .S(n2413), .Y(n2361) );
  MUX2X1 U2572 ( .B(\mem<54><7> ), .A(\mem<55><7> ), .S(n2443), .Y(n2355) );
  MUX2X1 U2573 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n2443), .Y(n2354) );
  MUX2X1 U2574 ( .B(\mem<50><7> ), .A(\mem<51><7> ), .S(n2443), .Y(n2358) );
  MUX2X1 U2575 ( .B(\mem<48><7> ), .A(\mem<49><7> ), .S(n2443), .Y(n2357) );
  MUX2X1 U2576 ( .B(n2356), .A(n2353), .S(n2413), .Y(n2360) );
  MUX2X1 U2577 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n2444), .Y(n2364) );
  MUX2X1 U2578 ( .B(\mem<44><7> ), .A(\mem<45><7> ), .S(n2444), .Y(n2363) );
  MUX2X1 U2579 ( .B(\mem<42><7> ), .A(\mem<43><7> ), .S(n2444), .Y(n2367) );
  MUX2X1 U2580 ( .B(\mem<40><7> ), .A(\mem<41><7> ), .S(n2444), .Y(n2366) );
  MUX2X1 U2581 ( .B(n2365), .A(n2362), .S(n2413), .Y(n2376) );
  MUX2X1 U2582 ( .B(\mem<38><7> ), .A(\mem<39><7> ), .S(n2444), .Y(n2370) );
  MUX2X1 U2583 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n2444), .Y(n2369) );
  MUX2X1 U2584 ( .B(\mem<34><7> ), .A(\mem<35><7> ), .S(n2444), .Y(n2373) );
  MUX2X1 U2585 ( .B(\mem<32><7> ), .A(\mem<33><7> ), .S(n2444), .Y(n2372) );
  MUX2X1 U2586 ( .B(n2371), .A(n2368), .S(n2413), .Y(n2375) );
  MUX2X1 U2587 ( .B(n2374), .A(n2359), .S(n2409), .Y(n2408) );
  MUX2X1 U2588 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n2444), .Y(n2379) );
  MUX2X1 U2589 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n2444), .Y(n2378) );
  MUX2X1 U2590 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n2444), .Y(n2382) );
  MUX2X1 U2591 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n2444), .Y(n2381) );
  MUX2X1 U2592 ( .B(n2380), .A(n2377), .S(n2413), .Y(n2391) );
  MUX2X1 U2593 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n2437), .Y(n2385) );
  MUX2X1 U2594 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n2435), .Y(n2384) );
  MUX2X1 U2595 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n2435), .Y(n2388) );
  MUX2X1 U2596 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n2435), .Y(n2387) );
  MUX2X1 U2597 ( .B(n2386), .A(n2383), .S(n2414), .Y(n2390) );
  MUX2X1 U2598 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n2435), .Y(n2394) );
  MUX2X1 U2599 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n2435), .Y(n2393) );
  MUX2X1 U2600 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n2438), .Y(n2397) );
  MUX2X1 U2601 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n2434), .Y(n2396) );
  MUX2X1 U2602 ( .B(n2395), .A(n2392), .S(n2413), .Y(n2406) );
  MUX2X1 U2603 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n2435), .Y(n2400) );
  MUX2X1 U2604 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n2437), .Y(n2399) );
  MUX2X1 U2605 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n2436), .Y(n2403) );
  MUX2X1 U2606 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n2437), .Y(n2402) );
  MUX2X1 U2607 ( .B(n2401), .A(n2398), .S(n2415), .Y(n2405) );
  MUX2X1 U2608 ( .B(n2404), .A(n2389), .S(n2409), .Y(n2407) );
  INVX2 U2609 ( .A(Wr), .Y(n2548) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module fetch ( .BranchPC({\BranchPC<15> , \BranchPC<14> , \BranchPC<13> , 
        \BranchPC<12> , \BranchPC<11> , \BranchPC<10> , \BranchPC<9> , 
        \BranchPC<8> , \BranchPC<7> , \BranchPC<6> , \BranchPC<5> , 
        \BranchPC<4> , \BranchPC<3> , \BranchPC<2> , \BranchPC<1> , 
        \BranchPC<0> }), BranchJumpTaken, clk, rst, Halt, Rti, Exception, 
        Stall, .Instr({\Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , 
        \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , 
        \Instr<0> }), .IncPC({\IncPC<15> , \IncPC<14> , \IncPC<13> , 
        \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , 
        \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , 
        \IncPC<1> , \IncPC<0> }), Err, CacheHit, InstrMemStall );
  input \BranchPC<15> , \BranchPC<14> , \BranchPC<13> , \BranchPC<12> ,
         \BranchPC<11> , \BranchPC<10> , \BranchPC<9> , \BranchPC<8> ,
         \BranchPC<7> , \BranchPC<6> , \BranchPC<5> , \BranchPC<4> ,
         \BranchPC<3> , \BranchPC<2> , \BranchPC<1> , \BranchPC<0> ,
         BranchJumpTaken, clk, rst, Halt, Rti, Exception, Stall;
  output \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> ,
         \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> ,
         \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> ,
         \Instr<0> , \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> ,
         \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> ,
         \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> ,
         \IncPC<1> , \IncPC<0> , Err, CacheHit, InstrMemStall;
  wire   \pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , \pc<10> , \pc<9> ,
         \pc<8> , \pc<7> , \pc<6> , \pc<5> , \pc<4> , \pc<3> , \pc<2> ,
         \pc<1> , \pc<0> , \nextEPC<15> , \nextEPC<14> , \nextEPC<13> ,
         \nextEPC<12> , \nextEPC<11> , \nextEPC<10> , \nextEPC<9> ,
         \nextEPC<8> , \nextEPC<7> , \nextEPC<6> , \nextEPC<5> , \nextEPC<4> ,
         \nextEPC<3> , \nextEPC<2> , \nextEPC<1> , \nextEPC<0> , \epc<15> ,
         \epc<14> , \epc<13> , \epc<12> , \epc<11> , \epc<10> , \epc<9> ,
         \epc<8> , \epc<7> , \epc<6> , \epc<5> , \epc<4> , \epc<3> , \epc<2> ,
         \epc<1> , \epc<0> , nextExcptState, curExcptState, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n58, n72, n75, n77, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73, n74, n76, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146;
  assign InstrMemStall = 1'b0;
  assign CacheHit = 1'b0;
  assign Err = 1'b0;

  XOR2X1 U25 ( .A(curExcptState), .B(Exception), .Y(n22) );
  OAI21X1 U26 ( .A(n23), .B(n135), .C(n24), .Y(\nextEPC<9> ) );
  NAND2X1 U27 ( .A(\epc<9> ), .B(n23), .Y(n24) );
  OAI21X1 U28 ( .A(n23), .B(n134), .C(n25), .Y(\nextEPC<8> ) );
  NAND2X1 U29 ( .A(\epc<8> ), .B(n23), .Y(n25) );
  OAI21X1 U30 ( .A(n23), .B(n133), .C(n26), .Y(\nextEPC<7> ) );
  NAND2X1 U31 ( .A(\epc<7> ), .B(n23), .Y(n26) );
  OAI21X1 U32 ( .A(n23), .B(n132), .C(n27), .Y(\nextEPC<6> ) );
  NAND2X1 U33 ( .A(\epc<6> ), .B(n23), .Y(n27) );
  OAI21X1 U34 ( .A(n23), .B(n131), .C(n28), .Y(\nextEPC<5> ) );
  NAND2X1 U35 ( .A(\epc<5> ), .B(n23), .Y(n28) );
  OAI21X1 U36 ( .A(n23), .B(n130), .C(n29), .Y(\nextEPC<4> ) );
  NAND2X1 U37 ( .A(\epc<4> ), .B(n23), .Y(n29) );
  OAI21X1 U38 ( .A(n23), .B(n143), .C(n30), .Y(\nextEPC<3> ) );
  NAND2X1 U39 ( .A(\epc<3> ), .B(n23), .Y(n30) );
  OAI21X1 U40 ( .A(n23), .B(n142), .C(n31), .Y(\nextEPC<2> ) );
  NAND2X1 U41 ( .A(\epc<2> ), .B(n23), .Y(n31) );
  OAI21X1 U42 ( .A(n23), .B(n144), .C(n32), .Y(\nextEPC<1> ) );
  NAND2X1 U43 ( .A(\epc<1> ), .B(n23), .Y(n32) );
  OAI21X1 U44 ( .A(n23), .B(n141), .C(n33), .Y(\nextEPC<15> ) );
  NAND2X1 U45 ( .A(\epc<15> ), .B(n23), .Y(n33) );
  OAI21X1 U46 ( .A(n23), .B(n140), .C(n34), .Y(\nextEPC<14> ) );
  NAND2X1 U47 ( .A(\epc<14> ), .B(n23), .Y(n34) );
  OAI21X1 U48 ( .A(n23), .B(n139), .C(n35), .Y(\nextEPC<13> ) );
  NAND2X1 U49 ( .A(\epc<13> ), .B(n23), .Y(n35) );
  OAI21X1 U50 ( .A(n23), .B(n138), .C(n36), .Y(\nextEPC<12> ) );
  NAND2X1 U51 ( .A(\epc<12> ), .B(n23), .Y(n36) );
  OAI21X1 U52 ( .A(n23), .B(n137), .C(n37), .Y(\nextEPC<11> ) );
  NAND2X1 U53 ( .A(\epc<11> ), .B(n23), .Y(n37) );
  OAI21X1 U54 ( .A(n23), .B(n136), .C(n38), .Y(\nextEPC<10> ) );
  NAND2X1 U55 ( .A(\epc<10> ), .B(n23), .Y(n38) );
  OAI21X1 U56 ( .A(n23), .B(n146), .C(n39), .Y(\nextEPC<0> ) );
  NAND2X1 U57 ( .A(\epc<0> ), .B(n23), .Y(n39) );
  AOI22X1 U84 ( .A(\IncPC<1> ), .B(n98), .C(\BranchPC<1> ), .D(n129), .Y(n58)
         );
  AOI22X1 U105 ( .A(\IncPC<0> ), .B(n98), .C(\BranchPC<0> ), .D(n129), .Y(n72)
         );
  NOR2X1 U108 ( .A(Stall), .B(Halt), .Y(n75) );
  NOR2X1 U110 ( .A(n105), .B(Halt), .Y(n77) );
  dff_388 \pc_reg[0]  ( .q(\pc<0> ), .d(n53), .clk(clk), .rst(n105) );
  dff_389 \pc_reg[1]  ( .q(\pc<1> ), .d(n55), .clk(clk), .rst(n105) );
  dff_390 \pc_reg[2]  ( .q(\pc<2> ), .d(n49), .clk(clk), .rst(rst) );
  dff_391 \pc_reg[3]  ( .q(\pc<3> ), .d(n47), .clk(clk), .rst(rst) );
  dff_392 \pc_reg[4]  ( .q(\pc<4> ), .d(n45), .clk(clk), .rst(rst) );
  dff_393 \pc_reg[5]  ( .q(\pc<5> ), .d(n43), .clk(clk), .rst(rst) );
  dff_394 \pc_reg[6]  ( .q(\pc<6> ), .d(n41), .clk(clk), .rst(n105) );
  dff_395 \pc_reg[7]  ( .q(\pc<7> ), .d(n21), .clk(clk), .rst(n105) );
  dff_396 \pc_reg[8]  ( .q(\pc<8> ), .d(n19), .clk(clk), .rst(n105) );
  dff_397 \pc_reg[9]  ( .q(\pc<9> ), .d(n17), .clk(clk), .rst(n105) );
  dff_398 \pc_reg[10]  ( .q(\pc<10> ), .d(n15), .clk(clk), .rst(n105) );
  dff_399 \pc_reg[11]  ( .q(\pc<11> ), .d(n13), .clk(clk), .rst(n105) );
  dff_400 \pc_reg[12]  ( .q(\pc<12> ), .d(n11), .clk(clk), .rst(n105) );
  dff_401 \pc_reg[13]  ( .q(\pc<13> ), .d(n9), .clk(clk), .rst(n105) );
  dff_402 \pc_reg[14]  ( .q(\pc<14> ), .d(n7), .clk(clk), .rst(n105) );
  dff_403 \pc_reg[15]  ( .q(\pc<15> ), .d(n5), .clk(clk), .rst(n105) );
  dff_372 \epc_reg[0]  ( .q(\epc<0> ), .d(\nextEPC<0> ), .clk(clk), .rst(n105)
         );
  dff_373 \epc_reg[1]  ( .q(\epc<1> ), .d(\nextEPC<1> ), .clk(clk), .rst(n105)
         );
  dff_374 \epc_reg[2]  ( .q(\epc<2> ), .d(\nextEPC<2> ), .clk(clk), .rst(n105)
         );
  dff_375 \epc_reg[3]  ( .q(\epc<3> ), .d(\nextEPC<3> ), .clk(clk), .rst(n105)
         );
  dff_376 \epc_reg[4]  ( .q(\epc<4> ), .d(\nextEPC<4> ), .clk(clk), .rst(n105)
         );
  dff_377 \epc_reg[5]  ( .q(\epc<5> ), .d(\nextEPC<5> ), .clk(clk), .rst(n105)
         );
  dff_378 \epc_reg[6]  ( .q(\epc<6> ), .d(\nextEPC<6> ), .clk(clk), .rst(n105)
         );
  dff_379 \epc_reg[7]  ( .q(\epc<7> ), .d(\nextEPC<7> ), .clk(clk), .rst(n105)
         );
  dff_380 \epc_reg[8]  ( .q(\epc<8> ), .d(\nextEPC<8> ), .clk(clk), .rst(n105)
         );
  dff_381 \epc_reg[9]  ( .q(\epc<9> ), .d(\nextEPC<9> ), .clk(clk), .rst(n105)
         );
  dff_382 \epc_reg[10]  ( .q(\epc<10> ), .d(\nextEPC<10> ), .clk(clk), .rst(
        n105) );
  dff_383 \epc_reg[11]  ( .q(\epc<11> ), .d(\nextEPC<11> ), .clk(clk), .rst(
        n105) );
  dff_384 \epc_reg[12]  ( .q(\epc<12> ), .d(\nextEPC<12> ), .clk(clk), .rst(
        n105) );
  dff_385 \epc_reg[13]  ( .q(\epc<13> ), .d(\nextEPC<13> ), .clk(clk), .rst(
        n105) );
  dff_386 \epc_reg[14]  ( .q(\epc<14> ), .d(\nextEPC<14> ), .clk(clk), .rst(
        n105) );
  dff_387 \epc_reg[15]  ( .q(\epc<15> ), .d(\nextEPC<15> ), .clk(clk), .rst(
        n105) );
  dff_404 excpt_reg ( .q(curExcptState), .d(nextExcptState), .clk(clk), .rst(
        n105) );
  memory2c instr_mem ( .data_out({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , 
        \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , 
        \Instr<1> , \Instr<0> }), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .addr({
        \pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , \pc<10> , \pc<9> , 
        \pc<8> , \pc<7> , \pc<6> , \pc<5> , n103, n101, n99, \pc<1> , \pc<0> }), .enable(1'b1), .wr(1'b0), .createdump(1'b0), .clk(clk), .rst(n105) );
  cla16_2 pc_inc ( .A({\pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , 
        \pc<10> , \pc<9> , \pc<8> , \pc<7> , \pc<6> , \pc<5> , n103, n101, n99, 
        \pc<1> , \pc<0> }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .Cin(1'b0), .S({
        \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> , 
        \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> , 
        \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> }), .Cout() );
  INVX1 U6 ( .A(\pc<2> ), .Y(n100) );
  INVX1 U7 ( .A(\pc<4> ), .Y(n104) );
  AND2X1 U8 ( .A(\BranchPC<2> ), .B(n129), .Y(n95) );
  AND2X1 U9 ( .A(\BranchPC<3> ), .B(n129), .Y(n93) );
  AND2X1 U10 ( .A(\BranchPC<4> ), .B(n129), .Y(n91) );
  AND2X1 U11 ( .A(\BranchPC<5> ), .B(n129), .Y(n89) );
  AND2X1 U12 ( .A(\BranchPC<6> ), .B(n129), .Y(n87) );
  AND2X1 U13 ( .A(\BranchPC<8> ), .B(n129), .Y(n83) );
  AND2X1 U14 ( .A(\BranchPC<9> ), .B(n129), .Y(n81) );
  INVX1 U15 ( .A(\IncPC<3> ), .Y(n143) );
  INVX1 U16 ( .A(\IncPC<6> ), .Y(n132) );
  INVX1 U17 ( .A(\IncPC<7> ), .Y(n133) );
  INVX1 U18 ( .A(\IncPC<9> ), .Y(n135) );
  INVX1 U19 ( .A(\IncPC<10> ), .Y(n136) );
  INVX1 U20 ( .A(\IncPC<11> ), .Y(n137) );
  INVX1 U21 ( .A(\IncPC<12> ), .Y(n138) );
  INVX1 U22 ( .A(\IncPC<13> ), .Y(n139) );
  INVX1 U23 ( .A(\IncPC<14> ), .Y(n140) );
  INVX1 U24 ( .A(\IncPC<15> ), .Y(n141) );
  INVX1 U58 ( .A(Rti), .Y(n145) );
  INVX1 U59 ( .A(Halt), .Y(n107) );
  INVX2 U60 ( .A(rst), .Y(n106) );
  INVX1 U61 ( .A(\pc<3> ), .Y(n102) );
  INVX1 U62 ( .A(\IncPC<0> ), .Y(n146) );
  INVX1 U63 ( .A(\IncPC<1> ), .Y(n144) );
  INVX1 U64 ( .A(\IncPC<2> ), .Y(n142) );
  INVX1 U65 ( .A(\IncPC<4> ), .Y(n130) );
  INVX1 U66 ( .A(\IncPC<5> ), .Y(n131) );
  INVX1 U67 ( .A(\IncPC<8> ), .Y(n134) );
  AND2X1 U68 ( .A(n22), .B(n145), .Y(nextExcptState) );
  INVX2 U69 ( .A(n100), .Y(n99) );
  AND2X1 U70 ( .A(curExcptState), .B(n145), .Y(n23) );
  AND2X1 U71 ( .A(\BranchPC<11> ), .B(n129), .Y(n76) );
  AND2X1 U72 ( .A(\BranchPC<12> ), .B(n129), .Y(n73) );
  AND2X1 U73 ( .A(\BranchPC<14> ), .B(n129), .Y(n70) );
  AND2X1 U74 ( .A(\BranchPC<15> ), .B(n129), .Y(n68) );
  AND2X1 U75 ( .A(\BranchPC<10> ), .B(n129), .Y(n79) );
  AND2X1 U76 ( .A(\BranchPC<7> ), .B(n129), .Y(n85) );
  AND2X2 U77 ( .A(n113), .B(n69), .Y(n4) );
  INVX1 U78 ( .A(n4), .Y(n5) );
  AND2X2 U79 ( .A(n114), .B(n71), .Y(n6) );
  INVX1 U80 ( .A(n6), .Y(n7) );
  AND2X2 U81 ( .A(n115), .B(n51), .Y(n8) );
  INVX1 U82 ( .A(n8), .Y(n9) );
  AND2X2 U83 ( .A(n116), .B(n74), .Y(n10) );
  INVX1 U85 ( .A(n10), .Y(n11) );
  AND2X2 U86 ( .A(n117), .B(n78), .Y(n12) );
  INVX1 U87 ( .A(n12), .Y(n13) );
  AND2X2 U88 ( .A(n118), .B(n80), .Y(n14) );
  INVX1 U89 ( .A(n14), .Y(n15) );
  AND2X2 U90 ( .A(n119), .B(n82), .Y(n16) );
  INVX1 U91 ( .A(n16), .Y(n17) );
  AND2X2 U92 ( .A(n120), .B(n84), .Y(n18) );
  INVX1 U93 ( .A(n18), .Y(n19) );
  AND2X2 U94 ( .A(n121), .B(n86), .Y(n20) );
  INVX1 U95 ( .A(n20), .Y(n21) );
  AND2X2 U96 ( .A(n122), .B(n88), .Y(n40) );
  INVX1 U97 ( .A(n40), .Y(n41) );
  AND2X2 U98 ( .A(n123), .B(n90), .Y(n42) );
  INVX1 U99 ( .A(n42), .Y(n43) );
  AND2X2 U100 ( .A(n124), .B(n92), .Y(n44) );
  INVX1 U101 ( .A(n44), .Y(n45) );
  AND2X2 U102 ( .A(n125), .B(n94), .Y(n46) );
  INVX1 U103 ( .A(n46), .Y(n47) );
  AND2X2 U104 ( .A(n126), .B(n96), .Y(n48) );
  INVX1 U106 ( .A(n48), .Y(n49) );
  AND2X2 U107 ( .A(n129), .B(\BranchPC<13> ), .Y(n50) );
  INVX1 U109 ( .A(n50), .Y(n51) );
  AND2X2 U111 ( .A(n65), .B(n57), .Y(n52) );
  INVX1 U112 ( .A(n52), .Y(n53) );
  AND2X2 U113 ( .A(n67), .B(n60), .Y(n54) );
  INVX1 U114 ( .A(n54), .Y(n55) );
  AND2X2 U115 ( .A(\pc<0> ), .B(n128), .Y(n56) );
  INVX1 U116 ( .A(n56), .Y(n57) );
  AND2X2 U117 ( .A(\pc<1> ), .B(n128), .Y(n59) );
  INVX1 U118 ( .A(n59), .Y(n60) );
  BUFX2 U119 ( .A(n108), .Y(n61) );
  BUFX2 U120 ( .A(BranchJumpTaken), .Y(n62) );
  BUFX2 U121 ( .A(n111), .Y(n63) );
  INVX1 U122 ( .A(n72), .Y(n64) );
  INVX1 U123 ( .A(n64), .Y(n65) );
  INVX1 U124 ( .A(n58), .Y(n66) );
  INVX1 U125 ( .A(n66), .Y(n67) );
  INVX1 U126 ( .A(n68), .Y(n69) );
  INVX1 U127 ( .A(n70), .Y(n71) );
  INVX1 U128 ( .A(n73), .Y(n74) );
  INVX1 U129 ( .A(n76), .Y(n78) );
  INVX1 U130 ( .A(n79), .Y(n80) );
  INVX1 U131 ( .A(n81), .Y(n82) );
  INVX1 U132 ( .A(n83), .Y(n84) );
  INVX1 U133 ( .A(n85), .Y(n86) );
  INVX1 U134 ( .A(n87), .Y(n88) );
  INVX1 U135 ( .A(n89), .Y(n90) );
  INVX1 U136 ( .A(n91), .Y(n92) );
  INVX1 U137 ( .A(n93), .Y(n94) );
  INVX1 U138 ( .A(n95), .Y(n96) );
  INVX1 U139 ( .A(n109), .Y(n129) );
  INVX1 U140 ( .A(n62), .Y(n110) );
  INVX1 U141 ( .A(n61), .Y(n128) );
  BUFX4 U142 ( .A(n127), .Y(n97) );
  BUFX4 U143 ( .A(n127), .Y(n98) );
  INVX8 U144 ( .A(n102), .Y(n101) );
  INVX8 U145 ( .A(n104), .Y(n103) );
  INVX8 U146 ( .A(n106), .Y(n105) );
  NAND3X1 U147 ( .A(n62), .B(n107), .C(n106), .Y(n109) );
  NAND3X1 U148 ( .A(n77), .B(Stall), .C(n110), .Y(n108) );
  AND2X2 U149 ( .A(n61), .B(n109), .Y(n112) );
  NAND3X1 U150 ( .A(n105), .B(n110), .C(n75), .Y(n111) );
  AND2X2 U151 ( .A(n112), .B(n63), .Y(n127) );
  AOI22X1 U152 ( .A(\pc<15> ), .B(n128), .C(\IncPC<15> ), .D(n97), .Y(n113) );
  AOI22X1 U153 ( .A(\pc<14> ), .B(n128), .C(\IncPC<14> ), .D(n97), .Y(n114) );
  AOI22X1 U154 ( .A(\pc<13> ), .B(n128), .C(\IncPC<13> ), .D(n97), .Y(n115) );
  AOI22X1 U155 ( .A(\pc<12> ), .B(n128), .C(\IncPC<12> ), .D(n97), .Y(n116) );
  AOI22X1 U156 ( .A(\pc<11> ), .B(n128), .C(\IncPC<11> ), .D(n97), .Y(n117) );
  AOI22X1 U157 ( .A(\pc<10> ), .B(n128), .C(\IncPC<10> ), .D(n97), .Y(n118) );
  AOI22X1 U158 ( .A(\pc<9> ), .B(n128), .C(\IncPC<9> ), .D(n97), .Y(n119) );
  AOI22X1 U159 ( .A(\pc<8> ), .B(n128), .C(\IncPC<8> ), .D(n97), .Y(n120) );
  AOI22X1 U160 ( .A(\pc<7> ), .B(n128), .C(\IncPC<7> ), .D(n98), .Y(n121) );
  AOI22X1 U161 ( .A(\pc<6> ), .B(n128), .C(\IncPC<6> ), .D(n98), .Y(n122) );
  AOI22X1 U162 ( .A(\pc<5> ), .B(n128), .C(\IncPC<5> ), .D(n98), .Y(n123) );
  AOI22X1 U163 ( .A(n103), .B(n128), .C(\IncPC<4> ), .D(n98), .Y(n124) );
  AOI22X1 U164 ( .A(n101), .B(n128), .C(\IncPC<3> ), .D(n98), .Y(n125) );
  AOI22X1 U165 ( .A(n99), .B(n128), .C(\IncPC<2> ), .D(n98), .Y(n126) );
endmodule


module pipe_fd ( Stall, Flush, rst, clk, .Instr({\Instr<15> , \Instr<14> , 
        \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , 
        \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , 
        \Instr<2> , \Instr<1> , \Instr<0> }), .IncPC({\IncPC<15> , \IncPC<14> , 
        \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , 
        \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , 
        \IncPC<2> , \IncPC<1> , \IncPC<0> }), .Instr_Out({\Instr_Out<15> , 
        \Instr_Out<14> , \Instr_Out<13> , \Instr_Out<12> , \Instr_Out<11> , 
        \Instr_Out<10> , \Instr_Out<9> , \Instr_Out<8> , \Instr_Out<7> , 
        \Instr_Out<6> , \Instr_Out<5> , \Instr_Out<4> , \Instr_Out<3> , 
        \Instr_Out<2> , \Instr_Out<1> , \Instr_Out<0> }), .IncPC_Out({
        \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> , \IncPC_Out<12> , 
        \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> , \IncPC_Out<8> , 
        \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> , \IncPC_Out<4> , 
        \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> , \IncPC_Out<0> }), 
        CPUActive );
  input Stall, Flush, rst, clk, \Instr<15> , \Instr<14> , \Instr<13> ,
         \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> ,
         \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> ,
         \Instr<2> , \Instr<1> , \Instr<0> , \IncPC<15> , \IncPC<14> ,
         \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> ,
         \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> ,
         \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> ;
  output \Instr_Out<15> , \Instr_Out<14> , \Instr_Out<13> , \Instr_Out<12> ,
         \Instr_Out<11> , \Instr_Out<10> , \Instr_Out<9> , \Instr_Out<8> ,
         \Instr_Out<7> , \Instr_Out<6> , \Instr_Out<5> , \Instr_Out<4> ,
         \Instr_Out<3> , \Instr_Out<2> , \Instr_Out<1> , \Instr_Out<0> ,
         \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> , \IncPC_Out<12> ,
         \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> , \IncPC_Out<8> ,
         \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> , \IncPC_Out<4> ,
         \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> , \IncPC_Out<0> ,
         CPUActive;
  wire   \Instr_Muxed<11> , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n70, n71, n72, n73, n74, n75, n76;

  AOI22X1 U37 ( .A(\Instr_Out<9> ), .B(n4), .C(\Instr<9> ), .D(n6), .Y(n36) );
  AOI22X1 U38 ( .A(\Instr_Out<8> ), .B(n4), .C(\Instr<8> ), .D(n6), .Y(n39) );
  AOI22X1 U39 ( .A(\Instr_Out<7> ), .B(n4), .C(\Instr<7> ), .D(n6), .Y(n40) );
  AOI22X1 U40 ( .A(\Instr_Out<6> ), .B(n4), .C(\Instr<6> ), .D(n6), .Y(n41) );
  AOI22X1 U41 ( .A(\Instr_Out<5> ), .B(n4), .C(\Instr<5> ), .D(n6), .Y(n42) );
  AOI22X1 U42 ( .A(\Instr_Out<4> ), .B(n4), .C(\Instr<4> ), .D(n6), .Y(n43) );
  AOI22X1 U43 ( .A(\Instr_Out<3> ), .B(n4), .C(\Instr<3> ), .D(n6), .Y(n44) );
  AOI22X1 U44 ( .A(\Instr_Out<2> ), .B(n4), .C(\Instr<2> ), .D(n6), .Y(n45) );
  AOI22X1 U45 ( .A(\Instr_Out<1> ), .B(n4), .C(\Instr<1> ), .D(n5), .Y(n46) );
  AOI22X1 U46 ( .A(\Instr_Out<15> ), .B(n4), .C(\Instr<15> ), .D(n5), .Y(n47)
         );
  AOI22X1 U47 ( .A(\Instr_Out<14> ), .B(n4), .C(\Instr<14> ), .D(n5), .Y(n48)
         );
  AOI22X1 U48 ( .A(\Instr_Out<13> ), .B(n4), .C(\Instr<13> ), .D(n5), .Y(n49)
         );
  AOI22X1 U49 ( .A(\Instr_Out<12> ), .B(n4), .C(\Instr<12> ), .D(n5), .Y(n50)
         );
  NAND3X1 U50 ( .A(n10), .B(n9), .C(n51), .Y(\Instr_Muxed<11> ) );
  AOI22X1 U51 ( .A(\Instr_Out<11> ), .B(n4), .C(\Instr<11> ), .D(n5), .Y(n51)
         );
  AOI22X1 U52 ( .A(\Instr_Out<10> ), .B(n4), .C(\Instr<10> ), .D(n5), .Y(n52)
         );
  AOI22X1 U53 ( .A(\Instr_Out<0> ), .B(n4), .C(\Instr<0> ), .D(n5), .Y(n53) );
  NOR3X1 U54 ( .A(n2), .B(n7), .C(Flush), .Y(n38) );
  NOR3X1 U55 ( .A(Flush), .B(n7), .C(n76), .Y(n37) );
  AOI22X1 U56 ( .A(\IncPC<9> ), .B(n76), .C(\IncPC_Out<9> ), .D(n2), .Y(n54)
         );
  AOI22X1 U57 ( .A(\IncPC<8> ), .B(n76), .C(\IncPC_Out<8> ), .D(n2), .Y(n55)
         );
  AOI22X1 U58 ( .A(\IncPC<7> ), .B(n76), .C(\IncPC_Out<7> ), .D(n2), .Y(n56)
         );
  AOI22X1 U59 ( .A(\IncPC<6> ), .B(n76), .C(\IncPC_Out<6> ), .D(n2), .Y(n57)
         );
  AOI22X1 U60 ( .A(\IncPC<5> ), .B(n76), .C(\IncPC_Out<5> ), .D(n2), .Y(n58)
         );
  AOI22X1 U61 ( .A(\IncPC<4> ), .B(n76), .C(\IncPC_Out<4> ), .D(n2), .Y(n59)
         );
  AOI22X1 U62 ( .A(\IncPC<3> ), .B(n76), .C(\IncPC_Out<3> ), .D(n2), .Y(n60)
         );
  AOI22X1 U63 ( .A(\IncPC<2> ), .B(n76), .C(\IncPC_Out<2> ), .D(n2), .Y(n61)
         );
  AOI22X1 U64 ( .A(\IncPC<1> ), .B(n76), .C(\IncPC_Out<1> ), .D(n3), .Y(n62)
         );
  AOI22X1 U65 ( .A(\IncPC<15> ), .B(n76), .C(\IncPC_Out<15> ), .D(n3), .Y(n63)
         );
  AOI22X1 U66 ( .A(\IncPC<14> ), .B(n76), .C(\IncPC_Out<14> ), .D(n3), .Y(n64)
         );
  AOI22X1 U67 ( .A(\IncPC<13> ), .B(n76), .C(\IncPC_Out<13> ), .D(n3), .Y(n65)
         );
  AOI22X1 U68 ( .A(\IncPC<12> ), .B(n76), .C(\IncPC_Out<12> ), .D(n3), .Y(n66)
         );
  AOI22X1 U69 ( .A(\IncPC<11> ), .B(n76), .C(\IncPC_Out<11> ), .D(n3), .Y(n67)
         );
  AOI22X1 U70 ( .A(\IncPC<10> ), .B(n76), .C(\IncPC_Out<10> ), .D(n3), .Y(n68)
         );
  AOI22X1 U71 ( .A(\IncPC<0> ), .B(n76), .C(\IncPC_Out<0> ), .D(n3), .Y(n69)
         );
  dff_355 \instr_reg[0]  ( .q(\Instr_Out<0> ), .d(n33), .clk(clk), .rst(1'b0)
         );
  dff_356 \instr_reg[1]  ( .q(\Instr_Out<1> ), .d(n34), .clk(clk), .rst(1'b0)
         );
  dff_357 \instr_reg[2]  ( .q(\Instr_Out<2> ), .d(n35), .clk(clk), .rst(1'b0)
         );
  dff_358 \instr_reg[3]  ( .q(\Instr_Out<3> ), .d(n70), .clk(clk), .rst(1'b0)
         );
  dff_359 \instr_reg[4]  ( .q(\Instr_Out<4> ), .d(n71), .clk(clk), .rst(1'b0)
         );
  dff_360 \instr_reg[5]  ( .q(\Instr_Out<5> ), .d(n72), .clk(clk), .rst(1'b0)
         );
  dff_361 \instr_reg[6]  ( .q(\Instr_Out<6> ), .d(n73), .clk(clk), .rst(1'b0)
         );
  dff_362 \instr_reg[7]  ( .q(\Instr_Out<7> ), .d(n74), .clk(clk), .rst(1'b0)
         );
  dff_363 \instr_reg[8]  ( .q(\Instr_Out<8> ), .d(n32), .clk(clk), .rst(1'b0)
         );
  dff_364 \instr_reg[9]  ( .q(\Instr_Out<9> ), .d(n31), .clk(clk), .rst(1'b0)
         );
  dff_365 \instr_reg[10]  ( .q(\Instr_Out<10> ), .d(n30), .clk(clk), .rst(1'b0) );
  dff_366 \instr_reg[11]  ( .q(\Instr_Out<11> ), .d(n1), .clk(clk), .rst(1'b0)
         );
  dff_367 \instr_reg[12]  ( .q(\Instr_Out<12> ), .d(n29), .clk(clk), .rst(1'b0) );
  dff_368 \instr_reg[13]  ( .q(\Instr_Out<13> ), .d(n28), .clk(clk), .rst(1'b0) );
  dff_369 \instr_reg[14]  ( .q(\Instr_Out<14> ), .d(n27), .clk(clk), .rst(1'b0) );
  dff_370 \instr_reg[15]  ( .q(\Instr_Out<15> ), .d(n26), .clk(clk), .rst(1'b0) );
  dff_339 \incpc_reg[0]  ( .q(\IncPC_Out<0> ), .d(n75), .clk(clk), .rst(n8) );
  dff_340 \incpc_reg[1]  ( .q(\IncPC_Out<1> ), .d(n25), .clk(clk), .rst(n8) );
  dff_341 \incpc_reg[2]  ( .q(\IncPC_Out<2> ), .d(n23), .clk(clk), .rst(n8) );
  dff_342 \incpc_reg[3]  ( .q(\IncPC_Out<3> ), .d(n24), .clk(clk), .rst(n7) );
  dff_343 \incpc_reg[4]  ( .q(\IncPC_Out<4> ), .d(n11), .clk(clk), .rst(n7) );
  dff_344 \incpc_reg[5]  ( .q(\IncPC_Out<5> ), .d(n12), .clk(clk), .rst(n7) );
  dff_345 \incpc_reg[6]  ( .q(\IncPC_Out<6> ), .d(n13), .clk(clk), .rst(n7) );
  dff_346 \incpc_reg[7]  ( .q(\IncPC_Out<7> ), .d(n14), .clk(clk), .rst(n7) );
  dff_347 \incpc_reg[8]  ( .q(\IncPC_Out<8> ), .d(n15), .clk(clk), .rst(n7) );
  dff_348 \incpc_reg[9]  ( .q(\IncPC_Out<9> ), .d(n16), .clk(clk), .rst(n7) );
  dff_349 \incpc_reg[10]  ( .q(\IncPC_Out<10> ), .d(n17), .clk(clk), .rst(n7)
         );
  dff_350 \incpc_reg[11]  ( .q(\IncPC_Out<11> ), .d(n18), .clk(clk), .rst(n7)
         );
  dff_351 \incpc_reg[12]  ( .q(\IncPC_Out<12> ), .d(n19), .clk(clk), .rst(n7)
         );
  dff_352 \incpc_reg[13]  ( .q(\IncPC_Out<13> ), .d(n20), .clk(clk), .rst(n7)
         );
  dff_353 \incpc_reg[14]  ( .q(\IncPC_Out<14> ), .d(n21), .clk(clk), .rst(n7)
         );
  dff_354 \incpc_reg[15]  ( .q(\IncPC_Out<15> ), .d(n22), .clk(clk), .rst(n7)
         );
  dff_371 rst_ff ( .q(CPUActive), .d(n9), .clk(clk), .rst(n7) );
  BUFX2 U3 ( .A(n38), .Y(n6) );
  BUFX2 U4 ( .A(n38), .Y(n5) );
  INVX1 U5 ( .A(n9), .Y(n8) );
  BUFX2 U6 ( .A(Stall), .Y(n3) );
  INVX1 U7 ( .A(Flush), .Y(n10) );
  INVX1 U8 ( .A(rst), .Y(n9) );
  INVX2 U9 ( .A(n9), .Y(n7) );
  INVX1 U10 ( .A(n69), .Y(n75) );
  INVX1 U11 ( .A(n68), .Y(n17) );
  INVX1 U12 ( .A(n67), .Y(n18) );
  INVX1 U13 ( .A(n66), .Y(n19) );
  INVX1 U14 ( .A(n65), .Y(n20) );
  INVX1 U15 ( .A(n64), .Y(n21) );
  INVX1 U16 ( .A(n63), .Y(n22) );
  INVX1 U17 ( .A(n62), .Y(n25) );
  INVX1 U18 ( .A(n61), .Y(n23) );
  INVX1 U19 ( .A(n60), .Y(n24) );
  INVX1 U20 ( .A(n59), .Y(n11) );
  INVX1 U21 ( .A(n58), .Y(n12) );
  INVX1 U22 ( .A(n57), .Y(n13) );
  INVX1 U23 ( .A(n56), .Y(n14) );
  INVX1 U24 ( .A(n55), .Y(n15) );
  INVX1 U25 ( .A(n54), .Y(n16) );
  INVX1 U26 ( .A(n53), .Y(n33) );
  INVX1 U27 ( .A(n52), .Y(n30) );
  INVX1 U28 ( .A(n50), .Y(n29) );
  INVX1 U29 ( .A(n49), .Y(n28) );
  INVX1 U30 ( .A(n48), .Y(n27) );
  INVX1 U31 ( .A(n47), .Y(n26) );
  INVX1 U32 ( .A(n46), .Y(n34) );
  INVX1 U33 ( .A(n45), .Y(n35) );
  INVX1 U34 ( .A(n44), .Y(n70) );
  INVX1 U35 ( .A(n43), .Y(n71) );
  INVX1 U36 ( .A(n42), .Y(n72) );
  INVX1 U72 ( .A(n41), .Y(n73) );
  INVX1 U73 ( .A(n40), .Y(n74) );
  INVX1 U74 ( .A(n39), .Y(n32) );
  INVX1 U75 ( .A(n36), .Y(n31) );
  BUFX2 U76 ( .A(\Instr_Muxed<11> ), .Y(n1) );
  INVX8 U77 ( .A(n3), .Y(n76) );
  BUFX4 U78 ( .A(Stall), .Y(n2) );
  BUFX4 U79 ( .A(n37), .Y(n4) );
endmodule


module decode ( clk, rst, Stall, .Instr({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , 
        \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , 
        \Instr<1> , \Instr<0> }), .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .IncPC({\IncPC<15> , \IncPC<14> , 
        \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , 
        \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , 
        \IncPC<2> , \IncPC<1> , \IncPC<0> }), .ALUOp1({\ALUOp1<15> , 
        \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , 
        \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , 
        \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), 
    .ALUOp2({\ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , 
        \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , 
        \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , 
        \ALUOp2<1> , \ALUOp2<0> }), ALUSrc, .Immediate({\Immediate<15> , 
        \Immediate<14> , \Immediate<13> , \Immediate<12> , \Immediate<11> , 
        \Immediate<10> , \Immediate<9> , \Immediate<8> , \Immediate<7> , 
        \Immediate<6> , \Immediate<5> , \Immediate<4> , \Immediate<3> , 
        \Immediate<2> , \Immediate<1> , \Immediate<0> }), Branch, Jump, 
        JumpReg, Set, Btr, InvA, InvB, Cin, .ALUOpcode({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .Func({\Func<1> , \Func<0> }), 
        MemWrite, MemRead, MemToReg, Halt, Exception, Err, Rti, .Rs({\Rs<2> , 
        \Rs<1> , \Rs<0> }), .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({\Rd<2> , 
        \Rd<1> , \Rd<0> }), RegFileWrEn, RegFileWrEn_Out, .WriteReg({
        \WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), .WriteReg_Out({
        \WriteReg_Out<2> , \WriteReg_Out<1> , \WriteReg_Out<0> }), RtValid, 
        RsValid, RdValid, Link, Store );
  input clk, rst, Stall, \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> ,
         \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> ,
         \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> ,
         \Instr<1> , \Instr<0> , \WriteData<15> , \WriteData<14> ,
         \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> ,
         \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> ,
         \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> ,
         \WriteData<1> , \WriteData<0> , \IncPC<15> , \IncPC<14> , \IncPC<13> ,
         \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> ,
         \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> ,
         \IncPC<2> , \IncPC<1> , \IncPC<0> , RegFileWrEn, \WriteReg<2> ,
         \WriteReg<1> , \WriteReg<0> ;
  output \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> ,
         \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> ,
         \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> ,
         \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , ALUSrc, \Immediate<15> , \Immediate<14> ,
         \Immediate<13> , \Immediate<12> , \Immediate<11> , \Immediate<10> ,
         \Immediate<9> , \Immediate<8> , \Immediate<7> , \Immediate<6> ,
         \Immediate<5> , \Immediate<4> , \Immediate<3> , \Immediate<2> ,
         \Immediate<1> , \Immediate<0> , Branch, Jump, JumpReg, Set, Btr, InvA,
         InvB, Cin, \ALUOpcode<2> , \ALUOpcode<1> , \ALUOpcode<0> , \Func<1> ,
         \Func<0> , MemWrite, MemRead, MemToReg, Halt, Exception, Err, Rti,
         \Rs<2> , \Rs<1> , \Rs<0> , \Rt<2> , \Rt<1> , \Rt<0> , \Rd<2> ,
         \Rd<1> , \Rd<0> , RegFileWrEn_Out, \WriteReg_Out<2> ,
         \WriteReg_Out<1> , \WriteReg_Out<0> , RtValid, RsValid, RdValid, Link,
         Store;
  wire   Instr_15, Instr_14, Instr_13, n111, Rf, If1, If2, \rs_out<15> ,
         \rs_out<14> , \rs_out<13> , \rs_out<12> , \rs_out<11> , \rs_out<10> ,
         \rs_out<9> , \rs_out<8> , \rs_out<7> , \rs_out<6> , \rs_out<5> ,
         \rs_out<4> , \rs_out<3> , \rs_out<2> , \rs_out<1> , \rs_out<0> ,
         RfError, stu, slbi, lbi, ZeroExt, N73, N74, N75, N76, N77, N83, N84,
         n29, n30, n31, n38, n40, n42, n47, n48, n49, n55, n57, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n32, n33, n34, n35, n36, n37,
         n39, n41, n43, n44, n45, n46, n50, n51, n52, n53, n54, n56, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n78, n80, n82, n84, n89, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110;
  assign Instr_15 = \Instr<15> ;
  assign Instr_14 = \Instr<14> ;
  assign Instr_13 = \Instr<13> ;
  assign Err = 1'b0;

  LATCH \write_reg_reg<2>  ( .CLK(n22), .D(n19), .Q(\WriteReg_Out<2> ) );
  LATCH \write_reg_reg<1>  ( .CLK(n22), .D(n16), .Q(\WriteReg_Out<1> ) );
  LATCH \write_reg_reg<0>  ( .CLK(n22), .D(n13), .Q(\WriteReg_Out<0> ) );
  LATCH \ImmReg_reg<15>  ( .CLK(N83), .D(N84), .Q(\Immediate<15> ) );
  LATCH \ImmReg_reg<14>  ( .CLK(N83), .D(N84), .Q(\Immediate<14> ) );
  LATCH \ImmReg_reg<13>  ( .CLK(N83), .D(N84), .Q(\Immediate<13> ) );
  LATCH \ImmReg_reg<12>  ( .CLK(N83), .D(N84), .Q(\Immediate<12> ) );
  LATCH \ImmReg_reg<11>  ( .CLK(N83), .D(N84), .Q(\Immediate<11> ) );
  LATCH \ImmReg_reg<10>  ( .CLK(N83), .D(N84), .Q(\Immediate<10> ) );
  LATCH \ImmReg_reg<9>  ( .CLK(N83), .D(N77), .Q(\Immediate<9> ) );
  LATCH \ImmReg_reg<8>  ( .CLK(N83), .D(N76), .Q(\Immediate<8> ) );
  LATCH \ImmReg_reg<7>  ( .CLK(N83), .D(N75), .Q(\Immediate<7> ) );
  LATCH \ImmReg_reg<6>  ( .CLK(N83), .D(N74), .Q(\Immediate<6> ) );
  LATCH \ImmReg_reg<5>  ( .CLK(N83), .D(N73), .Q(\Immediate<5> ) );
  LATCH \ImmReg_reg<4>  ( .CLK(N83), .D(\Instr<4> ), .Q(\Immediate<4> ) );
  LATCH \ImmReg_reg<3>  ( .CLK(N83), .D(\Instr<3> ), .Q(\Immediate<3> ) );
  LATCH \ImmReg_reg<2>  ( .CLK(N83), .D(\Instr<2> ), .Q(\Immediate<2> ) );
  LATCH \ImmReg_reg<1>  ( .CLK(N83), .D(\Instr<1> ), .Q(\Immediate<1> ) );
  LATCH \ImmReg_reg<0>  ( .CLK(N83), .D(\Instr<0> ), .Q(\Immediate<0> ) );
  OR2X2 U3 ( .A(Instr_13), .B(Instr_14), .Y(n29) );
  OR2X2 U4 ( .A(RdValid), .B(If2), .Y(RsValid) );
  OR2X2 U5 ( .A(If1), .B(RtValid), .Y(RdValid) );
  AND2X2 U6 ( .A(Rf), .B(n31), .Y(RtValid) );
  NOR3X1 U42 ( .A(n29), .B(n110), .C(n30), .Y(Store) );
  XOR2X1 U43 ( .A(\Instr<12> ), .B(\Instr<11> ), .Y(n30) );
  NAND3X1 U44 ( .A(n107), .B(n109), .C(n11), .Y(n31) );
  OAI21X1 U46 ( .A(Rf), .B(n89), .C(n9), .Y(\Rd<2> ) );
  OAI21X1 U48 ( .A(Rf), .B(n78), .C(n7), .Y(\Rd<1> ) );
  OAI21X1 U50 ( .A(Rf), .B(n76), .C(n5), .Y(\Rd<0> ) );
  OAI21X1 U52 ( .A(Jump), .B(n65), .C(n102), .Y(N83) );
  OAI21X1 U53 ( .A(n24), .B(n91), .C(n92), .Y(N84) );
  OAI21X1 U54 ( .A(n24), .B(n82), .C(n92), .Y(N77) );
  OAI21X1 U55 ( .A(n24), .B(n80), .C(n92), .Y(N76) );
  OAI21X1 U56 ( .A(n89), .B(n73), .C(n40), .Y(n38) );
  OAI21X1 U57 ( .A(n102), .B(n89), .C(n40), .Y(N75) );
  OAI21X1 U58 ( .A(n102), .B(n78), .C(n40), .Y(N74) );
  OAI21X1 U59 ( .A(n102), .B(n76), .C(n40), .Y(N73) );
  NAND3X1 U60 ( .A(n64), .B(\Instr<4> ), .C(n59), .Y(n40) );
  NAND3X1 U62 ( .A(n73), .B(n24), .C(n56), .Y(n42) );
  AOI22X1 U68 ( .A(\Rs<2> ), .B(n48), .C(n49), .D(\Instr<4> ), .Y(n47) );
  AOI22X1 U73 ( .A(\Instr<9> ), .B(n48), .C(n49), .D(\Instr<3> ), .Y(n55) );
  AOI22X1 U76 ( .A(\Instr<8> ), .B(n48), .C(n49), .D(\Instr<2> ), .Y(n57) );
  NOR3X1 U77 ( .A(If1), .B(If2), .C(n106), .Y(n49) );
  OAI21X1 U78 ( .A(n70), .B(n104), .C(n63), .Y(n48) );
  OAI21X1 U85 ( .A(n75), .B(n94), .C(n52), .Y(\ALUOp1<9> ) );
  OAI21X1 U87 ( .A(n75), .B(n93), .C(n50), .Y(\ALUOp1<8> ) );
  OAI21X1 U89 ( .A(n75), .B(n100), .C(n45), .Y(\ALUOp1<15> ) );
  OAI21X1 U91 ( .A(n75), .B(n99), .C(n43), .Y(\ALUOp1<14> ) );
  OAI21X1 U93 ( .A(n75), .B(n98), .C(n39), .Y(\ALUOp1<13> ) );
  OAI21X1 U95 ( .A(n75), .B(n97), .C(n36), .Y(\ALUOp1<12> ) );
  OAI21X1 U97 ( .A(n75), .B(n96), .C(n34), .Y(\ALUOp1<11> ) );
  OAI21X1 U99 ( .A(n75), .B(n95), .C(n32), .Y(\ALUOp1<10> ) );
  rf_bypass regfile ( .read1data({\rs_out<15> , \rs_out<14> , \rs_out<13> , 
        \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> , \rs_out<8> , 
        \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> , \rs_out<3> , 
        \rs_out<2> , \rs_out<1> , \rs_out<0> }), .read2data({\ALUOp2<15> , 
        \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , 
        \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , 
        \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), 
        .err(RfError), .clk(clk), .rst(rst), .read1regsel({\Rs<2> , \Instr<9> , 
        \Instr<8> }), .read2regsel({\Rt<2> , \Instr<6> , \Instr<5> }), 
        .writeregsel({\WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), 
        .writedata({\WriteData<15> , \WriteData<14> , \WriteData<13> , 
        \WriteData<12> , \WriteData<11> , \WriteData<10> , \WriteData<9> , 
        \WriteData<8> , \WriteData<7> , \WriteData<6> , \WriteData<5> , 
        \WriteData<4> , \WriteData<3> , \WriteData<2> , \WriteData<1> , 
        \WriteData<0> }), .write(RegFileWrEn) );
  control_unit cu ( .opcode({Instr_15, Instr_14, Instr_13, \Instr<12> , 
        \Instr<11> }), .func({\Instr<1> , \Instr<0> }), .aluop({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .alusrc(ALUSrc), .branch(n111), 
        .jump(Jump), .i1(If1), .i2(If2), .r(Rf), .jumpreg(JumpReg), .set(Set), 
        .btr(Btr), .regwrite(RegFileWrEn_Out), .memwrite(MemWrite), .memread(
        MemRead), .memtoreg(MemToReg), .invA(InvA), .invB(InvB), .cin(Cin), 
        .excp(Exception), .zeroext(ZeroExt), .halt(Halt), .slbi(slbi), .link(
        Link), .lbi(lbi), .stu(stu), .rti(Rti) );
  INVX1 U7 ( .A(lbi), .Y(n101) );
  INVX1 U8 ( .A(Instr_13), .Y(n109) );
  INVX1 U9 ( .A(\Instr<12> ), .Y(n107) );
  AND2X1 U10 ( .A(\rs_out<2> ), .B(n61), .Y(\ALUOp1<2> ) );
  AND2X1 U11 ( .A(\rs_out<3> ), .B(n61), .Y(\ALUOp1<3> ) );
  AND2X1 U12 ( .A(\rs_out<4> ), .B(n61), .Y(\ALUOp1<4> ) );
  AND2X1 U13 ( .A(\rs_out<5> ), .B(n61), .Y(\ALUOp1<5> ) );
  AND2X1 U14 ( .A(\rs_out<6> ), .B(n61), .Y(\ALUOp1<6> ) );
  AND2X1 U15 ( .A(\rs_out<7> ), .B(n61), .Y(\ALUOp1<7> ) );
  INVX1 U16 ( .A(\rs_out<0> ), .Y(n93) );
  INVX1 U17 ( .A(\rs_out<1> ), .Y(n94) );
  INVX1 U18 ( .A(\rs_out<3> ), .Y(n96) );
  INVX1 U19 ( .A(\rs_out<4> ), .Y(n97) );
  INVX1 U20 ( .A(\rs_out<5> ), .Y(n98) );
  INVX1 U21 ( .A(\rs_out<6> ), .Y(n99) );
  INVX1 U22 ( .A(\Instr<7> ), .Y(n89) );
  INVX1 U23 ( .A(\Instr<10> ), .Y(n91) );
  INVX1 U24 ( .A(Instr_15), .Y(n110) );
  INVX1 U25 ( .A(ZeroExt), .Y(n105) );
  INVX1 U26 ( .A(If2), .Y(n103) );
  INVX1 U27 ( .A(stu), .Y(n104) );
  INVX1 U28 ( .A(Rf), .Y(n106) );
  AND2X1 U29 ( .A(\rs_out<0> ), .B(n61), .Y(\ALUOp1<0> ) );
  AND2X1 U30 ( .A(n61), .B(\rs_out<1> ), .Y(\ALUOp1<1> ) );
  INVX1 U31 ( .A(\rs_out<2> ), .Y(n95) );
  INVX1 U32 ( .A(\rs_out<7> ), .Y(n100) );
  INVX1 U33 ( .A(n38), .Y(n92) );
  INVX1 U34 ( .A(n91), .Y(\Rs<2> ) );
  INVX1 U35 ( .A(n89), .Y(\Rt<2> ) );
  AND2X1 U36 ( .A(n67), .B(n105), .Y(n72) );
  AND2X1 U37 ( .A(n69), .B(\Instr<6> ), .Y(n1) );
  AND2X1 U38 ( .A(n69), .B(\Instr<5> ), .Y(n2) );
  AND2X1 U39 ( .A(n69), .B(\Rt<2> ), .Y(n3) );
  INVX1 U40 ( .A(Jump), .Y(n108) );
  AND2X2 U41 ( .A(\Instr<2> ), .B(Rf), .Y(n4) );
  INVX1 U45 ( .A(n4), .Y(n5) );
  AND2X2 U47 ( .A(\Instr<3> ), .B(Rf), .Y(n6) );
  INVX1 U49 ( .A(n6), .Y(n7) );
  AND2X2 U51 ( .A(\Instr<4> ), .B(Rf), .Y(n8) );
  INVX1 U61 ( .A(n8), .Y(n9) );
  OR2X2 U63 ( .A(Instr_15), .B(Instr_14), .Y(n10) );
  INVX1 U64 ( .A(n10), .Y(n11) );
  BUFX2 U65 ( .A(n111), .Y(Branch) );
  OR2X1 U66 ( .A(n2), .B(n14), .Y(n13) );
  OR2X1 U67 ( .A(n15), .B(Link), .Y(n14) );
  INVX1 U69 ( .A(n57), .Y(n15) );
  OR2X1 U70 ( .A(n1), .B(n17), .Y(n16) );
  OR2X1 U71 ( .A(n18), .B(Link), .Y(n17) );
  INVX1 U72 ( .A(n55), .Y(n18) );
  OR2X1 U74 ( .A(n3), .B(n20), .Y(n19) );
  OR2X1 U75 ( .A(n21), .B(Link), .Y(n20) );
  INVX1 U79 ( .A(n47), .Y(n21) );
  OR2X1 U80 ( .A(n71), .B(n23), .Y(n22) );
  OR2X1 U81 ( .A(n26), .B(n62), .Y(n23) );
  OR2X1 U82 ( .A(n72), .B(n25), .Y(n24) );
  OR2X1 U83 ( .A(n27), .B(n108), .Y(n25) );
  OR2X1 U84 ( .A(n49), .B(Link), .Y(n26) );
  OR2X1 U86 ( .A(ZeroExt), .B(If1), .Y(n27) );
  AND2X1 U88 ( .A(\rs_out<10> ), .B(n61), .Y(n28) );
  INVX1 U90 ( .A(n28), .Y(n32) );
  AND2X1 U92 ( .A(\rs_out<11> ), .B(n61), .Y(n33) );
  INVX1 U94 ( .A(n33), .Y(n34) );
  AND2X1 U96 ( .A(\rs_out<12> ), .B(n61), .Y(n35) );
  INVX1 U98 ( .A(n35), .Y(n36) );
  AND2X1 U100 ( .A(\rs_out<13> ), .B(n61), .Y(n37) );
  INVX1 U101 ( .A(n37), .Y(n39) );
  AND2X1 U102 ( .A(\rs_out<14> ), .B(n61), .Y(n41) );
  INVX1 U103 ( .A(n41), .Y(n43) );
  AND2X1 U104 ( .A(\rs_out<15> ), .B(n61), .Y(n44) );
  INVX1 U105 ( .A(n44), .Y(n45) );
  AND2X1 U106 ( .A(\rs_out<8> ), .B(n61), .Y(n46) );
  INVX1 U107 ( .A(n46), .Y(n50) );
  AND2X1 U108 ( .A(\rs_out<9> ), .B(n61), .Y(n51) );
  INVX1 U109 ( .A(n51), .Y(n52) );
  BUFX2 U110 ( .A(n42), .Y(n53) );
  INVX1 U111 ( .A(n53), .Y(n102) );
  AND2X1 U112 ( .A(n67), .B(n108), .Y(n54) );
  INVX1 U113 ( .A(n54), .Y(n56) );
  OR2X1 U114 ( .A(ZeroExt), .B(Jump), .Y(n58) );
  INVX1 U115 ( .A(n58), .Y(n59) );
  OR2X1 U116 ( .A(lbi), .B(slbi), .Y(n60) );
  INVX1 U117 ( .A(n60), .Y(n61) );
  AND2X1 U118 ( .A(n67), .B(n106), .Y(n62) );
  INVX1 U119 ( .A(n62), .Y(n63) );
  AND2X1 U120 ( .A(If1), .B(n103), .Y(n64) );
  INVX1 U121 ( .A(n64), .Y(n65) );
  OR2X1 U122 ( .A(n103), .B(If1), .Y(n66) );
  INVX1 U123 ( .A(n66), .Y(n67) );
  OR2X1 U124 ( .A(n70), .B(stu), .Y(n68) );
  INVX1 U125 ( .A(n68), .Y(n69) );
  INVX1 U126 ( .A(n71), .Y(n70) );
  AND2X1 U127 ( .A(n64), .B(n106), .Y(n71) );
  INVX1 U128 ( .A(n72), .Y(n73) );
  AND2X1 U129 ( .A(slbi), .B(n101), .Y(n74) );
  INVX1 U130 ( .A(n74), .Y(n75) );
  INVX1 U131 ( .A(n107), .Y(\Func<1> ) );
  INVX1 U132 ( .A(n84), .Y(\Func<0> ) );
  INVX1 U133 ( .A(\Instr<11> ), .Y(n84) );
  INVX1 U134 ( .A(n82), .Y(\Rs<1> ) );
  INVX1 U135 ( .A(\Instr<9> ), .Y(n82) );
  INVX1 U136 ( .A(n80), .Y(\Rs<0> ) );
  INVX1 U137 ( .A(\Instr<8> ), .Y(n80) );
  INVX1 U138 ( .A(n78), .Y(\Rt<1> ) );
  INVX1 U139 ( .A(\Instr<6> ), .Y(n78) );
  INVX1 U140 ( .A(n76), .Y(\Rt<0> ) );
  INVX1 U141 ( .A(\Instr<5> ), .Y(n76) );
endmodule


module pipe_de ( clk, rst, Stall, Flush, .ALUOp1({\ALUOp1<15> , \ALUOp1<14> , 
        \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , 
        \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , 
        \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), .ALUOp2({
        \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , 
        \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , 
        \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , 
        \ALUOp2<0> }), .Immediate({\Immediate<15> , \Immediate<14> , 
        \Immediate<13> , \Immediate<12> , \Immediate<11> , \Immediate<10> , 
        \Immediate<9> , \Immediate<8> , \Immediate<7> , \Immediate<6> , 
        \Immediate<5> , \Immediate<4> , \Immediate<3> , \Immediate<2> , 
        \Immediate<1> , \Immediate<0> }), .ALUOpcode({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .Func({\Func<1> , \Func<0> }), 
        ALUSrc, Branch, Jump, JumpReg, Set, Btr, MemWrite, MemRead, MemToReg, 
        Halt, InvA, InvB, Cin, .IncPC({\IncPC<15> , \IncPC<14> , \IncPC<13> , 
        \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , 
        \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , 
        \IncPC<1> , \IncPC<0> }), CPUActive, .ALUOp1_Out({\ALUOp1_Out<15> , 
        \ALUOp1_Out<14> , \ALUOp1_Out<13> , \ALUOp1_Out<12> , \ALUOp1_Out<11> , 
        \ALUOp1_Out<10> , \ALUOp1_Out<9> , \ALUOp1_Out<8> , \ALUOp1_Out<7> , 
        \ALUOp1_Out<6> , \ALUOp1_Out<5> , \ALUOp1_Out<4> , \ALUOp1_Out<3> , 
        \ALUOp1_Out<2> , \ALUOp1_Out<1> , \ALUOp1_Out<0> }), .ALUOp2_Out({
        \ALUOp2_Out<15> , \ALUOp2_Out<14> , \ALUOp2_Out<13> , \ALUOp2_Out<12> , 
        \ALUOp2_Out<11> , \ALUOp2_Out<10> , \ALUOp2_Out<9> , \ALUOp2_Out<8> , 
        \ALUOp2_Out<7> , \ALUOp2_Out<6> , \ALUOp2_Out<5> , \ALUOp2_Out<4> , 
        \ALUOp2_Out<3> , \ALUOp2_Out<2> , \ALUOp2_Out<1> , \ALUOp2_Out<0> }), 
    .Immediate_Out({\Immediate_Out<15> , \Immediate_Out<14> , 
        \Immediate_Out<13> , \Immediate_Out<12> , \Immediate_Out<11> , 
        \Immediate_Out<10> , \Immediate_Out<9> , \Immediate_Out<8> , 
        \Immediate_Out<7> , \Immediate_Out<6> , \Immediate_Out<5> , 
        \Immediate_Out<4> , \Immediate_Out<3> , \Immediate_Out<2> , 
        \Immediate_Out<1> , \Immediate_Out<0> }), .ALUOpcode_Out({
        \ALUOpcode_Out<2> , \ALUOpcode_Out<1> , \ALUOpcode_Out<0> }), 
    .Func_Out({\Func_Out<1> , \Func_Out<0> }), ALUSrc_Out, Branch_Out, 
        Jump_Out, JumpReg_Out, Set_Out, Btr_Out, MemWrite_Out, MemRead_Out, 
        MemToReg_Out, Halt_Out, InvA_Out, InvB_Out, Cin_Out, .Rs({\Rs<2> , 
        \Rs<1> , \Rs<0> }), .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({\Rd<2> , 
        \Rd<1> , \Rd<0> }), .Rs_Out({\Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> }), 
    .Rt_Out({\Rt_Out<2> , \Rt_Out<1> , \Rt_Out<0> }), .Rd_Out({\Rd_Out<2> , 
        \Rd_Out<1> , \Rd_Out<0> }), RegFileWrEn, RegFileWrEn_Out, .IncPC_Out({
        \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> , \IncPC_Out<12> , 
        \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> , \IncPC_Out<8> , 
        \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> , \IncPC_Out<4> , 
        \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> , \IncPC_Out<0> }), 
    .WriteReg({\WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), .WriteReg_Out({
        \WriteReg_Out<2> , \WriteReg_Out<1> , \WriteReg_Out<0> }), RtValid, 
        RtValid_Out, CPUActive_Out, RsValid, RdValid, RsValid_Out, RdValid_Out, 
    .DecodeIncPC({\DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> , 
        \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> , 
        \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> , \DecodeIncPC<6> , 
        \DecodeIncPC<5> , \DecodeIncPC<4> , \DecodeIncPC<3> , \DecodeIncPC<2> , 
        \DecodeIncPC<1> , \DecodeIncPC<0> }), .DecodeIncPC_Out({
        \DecodeIncPC_Out<15> , \DecodeIncPC_Out<14> , \DecodeIncPC_Out<13> , 
        \DecodeIncPC_Out<12> , \DecodeIncPC_Out<11> , \DecodeIncPC_Out<10> , 
        \DecodeIncPC_Out<9> , \DecodeIncPC_Out<8> , \DecodeIncPC_Out<7> , 
        \DecodeIncPC_Out<6> , \DecodeIncPC_Out<5> , \DecodeIncPC_Out<4> , 
        \DecodeIncPC_Out<3> , \DecodeIncPC_Out<2> , \DecodeIncPC_Out<1> , 
        \DecodeIncPC_Out<0> }), Link, Link_Out );
  input clk, rst, Stall, Flush, \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> ,
         \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> ,
         \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> ,
         \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> ,
         \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> ,
         \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> ,
         \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> , \Immediate<15> ,
         \Immediate<14> , \Immediate<13> , \Immediate<12> , \Immediate<11> ,
         \Immediate<10> , \Immediate<9> , \Immediate<8> , \Immediate<7> ,
         \Immediate<6> , \Immediate<5> , \Immediate<4> , \Immediate<3> ,
         \Immediate<2> , \Immediate<1> , \Immediate<0> , \ALUOpcode<2> ,
         \ALUOpcode<1> , \ALUOpcode<0> , \Func<1> , \Func<0> , ALUSrc, Branch,
         Jump, JumpReg, Set, Btr, MemWrite, MemRead, MemToReg, Halt, InvA,
         InvB, Cin, \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> ,
         \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> ,
         \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> ,
         \IncPC<1> , \IncPC<0> , CPUActive, \Rs<2> , \Rs<1> , \Rs<0> , \Rt<2> ,
         \Rt<1> , \Rt<0> , \Rd<2> , \Rd<1> , \Rd<0> , RegFileWrEn,
         \WriteReg<2> , \WriteReg<1> , \WriteReg<0> , RtValid, RsValid,
         RdValid, \DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> ,
         \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> ,
         \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> ,
         \DecodeIncPC<6> , \DecodeIncPC<5> , \DecodeIncPC<4> ,
         \DecodeIncPC<3> , \DecodeIncPC<2> , \DecodeIncPC<1> ,
         \DecodeIncPC<0> , Link;
  output \ALUOp1_Out<15> , \ALUOp1_Out<14> , \ALUOp1_Out<13> ,
         \ALUOp1_Out<12> , \ALUOp1_Out<11> , \ALUOp1_Out<10> , \ALUOp1_Out<9> ,
         \ALUOp1_Out<8> , \ALUOp1_Out<7> , \ALUOp1_Out<6> , \ALUOp1_Out<5> ,
         \ALUOp1_Out<4> , \ALUOp1_Out<3> , \ALUOp1_Out<2> , \ALUOp1_Out<1> ,
         \ALUOp1_Out<0> , \ALUOp2_Out<15> , \ALUOp2_Out<14> , \ALUOp2_Out<13> ,
         \ALUOp2_Out<12> , \ALUOp2_Out<11> , \ALUOp2_Out<10> , \ALUOp2_Out<9> ,
         \ALUOp2_Out<8> , \ALUOp2_Out<7> , \ALUOp2_Out<6> , \ALUOp2_Out<5> ,
         \ALUOp2_Out<4> , \ALUOp2_Out<3> , \ALUOp2_Out<2> , \ALUOp2_Out<1> ,
         \ALUOp2_Out<0> , \Immediate_Out<15> , \Immediate_Out<14> ,
         \Immediate_Out<13> , \Immediate_Out<12> , \Immediate_Out<11> ,
         \Immediate_Out<10> , \Immediate_Out<9> , \Immediate_Out<8> ,
         \Immediate_Out<7> , \Immediate_Out<6> , \Immediate_Out<5> ,
         \Immediate_Out<4> , \Immediate_Out<3> , \Immediate_Out<2> ,
         \Immediate_Out<1> , \Immediate_Out<0> , \ALUOpcode_Out<2> ,
         \ALUOpcode_Out<1> , \ALUOpcode_Out<0> , \Func_Out<1> , \Func_Out<0> ,
         ALUSrc_Out, Branch_Out, Jump_Out, JumpReg_Out, Set_Out, Btr_Out,
         MemWrite_Out, MemRead_Out, MemToReg_Out, Halt_Out, InvA_Out, InvB_Out,
         Cin_Out, \Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> , \Rt_Out<2> ,
         \Rt_Out<1> , \Rt_Out<0> , \Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> ,
         RegFileWrEn_Out, \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> ,
         \IncPC_Out<12> , \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> ,
         \IncPC_Out<8> , \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> ,
         \IncPC_Out<4> , \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> ,
         \IncPC_Out<0> , \WriteReg_Out<2> , \WriteReg_Out<1> ,
         \WriteReg_Out<0> , RtValid_Out, CPUActive_Out, RsValid_Out,
         RdValid_Out, \DecodeIncPC_Out<15> , \DecodeIncPC_Out<14> ,
         \DecodeIncPC_Out<13> , \DecodeIncPC_Out<12> , \DecodeIncPC_Out<11> ,
         \DecodeIncPC_Out<10> , \DecodeIncPC_Out<9> , \DecodeIncPC_Out<8> ,
         \DecodeIncPC_Out<7> , \DecodeIncPC_Out<6> , \DecodeIncPC_Out<5> ,
         \DecodeIncPC_Out<4> , \DecodeIncPC_Out<3> , \DecodeIncPC_Out<2> ,
         \DecodeIncPC_Out<1> , \DecodeIncPC_Out<0> , Link_Out;
  wire   n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266;

  AOI22X1 U117 ( .A(\WriteReg<2> ), .B(n16), .C(\WriteReg_Out<2> ), .D(n6), 
        .Y(n118) );
  AOI22X1 U118 ( .A(\WriteReg<1> ), .B(n26), .C(\WriteReg_Out<1> ), .D(n6), 
        .Y(n119) );
  AOI22X1 U119 ( .A(\WriteReg<0> ), .B(n24), .C(\WriteReg_Out<0> ), .D(n6), 
        .Y(n120) );
  AOI22X1 U120 ( .A(Set), .B(n18), .C(Set_Out), .D(n6), .Y(n121) );
  AOI22X1 U121 ( .A(\Rt<2> ), .B(n18), .C(\Rt_Out<2> ), .D(n6), .Y(n122) );
  AOI22X1 U122 ( .A(\Rt<1> ), .B(n18), .C(\Rt_Out<1> ), .D(n6), .Y(n123) );
  AOI22X1 U123 ( .A(\Rt<0> ), .B(n18), .C(\Rt_Out<0> ), .D(n6), .Y(n124) );
  AOI22X1 U124 ( .A(RtValid), .B(n18), .C(RtValid_Out), .D(n6), .Y(n125) );
  AOI22X1 U125 ( .A(\Rs<2> ), .B(n18), .C(\Rs_Out<2> ), .D(n6), .Y(n126) );
  AOI22X1 U126 ( .A(\Rs<1> ), .B(n18), .C(\Rs_Out<1> ), .D(n6), .Y(n127) );
  AOI22X1 U127 ( .A(\Rs<0> ), .B(n18), .C(\Rs_Out<0> ), .D(n6), .Y(n128) );
  AOI22X1 U128 ( .A(RsValid), .B(n17), .C(RsValid_Out), .D(n6), .Y(n129) );
  AOI22X1 U129 ( .A(RegFileWrEn), .B(n17), .C(RegFileWrEn_Out), .D(n7), .Y(
        n130) );
  AOI22X1 U130 ( .A(\Rd<2> ), .B(n17), .C(\Rd_Out<2> ), .D(n7), .Y(n131) );
  AOI22X1 U131 ( .A(\Rd<1> ), .B(n17), .C(\Rd_Out<1> ), .D(n7), .Y(n132) );
  AOI22X1 U132 ( .A(\Rd<0> ), .B(n17), .C(\Rd_Out<0> ), .D(n7), .Y(n133) );
  AOI22X1 U133 ( .A(RdValid), .B(n17), .C(RdValid_Out), .D(n7), .Y(n134) );
  AOI22X1 U134 ( .A(MemWrite), .B(n17), .C(MemWrite_Out), .D(n7), .Y(n135) );
  AOI22X1 U135 ( .A(MemToReg), .B(n17), .C(MemToReg_Out), .D(n7), .Y(n136) );
  AOI22X1 U136 ( .A(MemRead), .B(n17), .C(MemRead_Out), .D(n7), .Y(n137) );
  AOI22X1 U137 ( .A(Link), .B(n17), .C(n3), .D(n7), .Y(n138) );
  AOI22X1 U138 ( .A(Jump), .B(n17), .C(Jump_Out), .D(n7), .Y(n139) );
  AOI22X1 U139 ( .A(JumpReg), .B(n18), .C(n4), .D(n7), .Y(n140) );
  AOI22X1 U140 ( .A(InvB), .B(n18), .C(InvB_Out), .D(n7), .Y(n141) );
  AOI22X1 U141 ( .A(InvA), .B(n18), .C(InvA_Out), .D(n8), .Y(n142) );
  AOI22X1 U142 ( .A(\IncPC<9> ), .B(n18), .C(\IncPC_Out<9> ), .D(n8), .Y(n143)
         );
  AOI22X1 U143 ( .A(\IncPC<8> ), .B(n18), .C(\IncPC_Out<8> ), .D(n8), .Y(n144)
         );
  AOI22X1 U144 ( .A(\IncPC<7> ), .B(n18), .C(\IncPC_Out<7> ), .D(n8), .Y(n145)
         );
  AOI22X1 U145 ( .A(\IncPC<6> ), .B(n18), .C(\IncPC_Out<6> ), .D(n8), .Y(n146)
         );
  AOI22X1 U146 ( .A(\IncPC<5> ), .B(n18), .C(\IncPC_Out<5> ), .D(n8), .Y(n147)
         );
  AOI22X1 U147 ( .A(\IncPC<4> ), .B(n18), .C(\IncPC_Out<4> ), .D(n8), .Y(n148)
         );
  AOI22X1 U148 ( .A(\IncPC<3> ), .B(n18), .C(\IncPC_Out<3> ), .D(n8), .Y(n149)
         );
  AOI22X1 U149 ( .A(\IncPC<2> ), .B(n18), .C(\IncPC_Out<2> ), .D(n8), .Y(n150)
         );
  AOI22X1 U150 ( .A(\IncPC<1> ), .B(n19), .C(\IncPC_Out<1> ), .D(n8), .Y(n151)
         );
  AOI22X1 U151 ( .A(\IncPC<15> ), .B(n19), .C(\IncPC_Out<15> ), .D(n8), .Y(
        n152) );
  AOI22X1 U152 ( .A(\IncPC<14> ), .B(n19), .C(\IncPC_Out<14> ), .D(n8), .Y(
        n153) );
  AOI22X1 U153 ( .A(\IncPC<13> ), .B(n19), .C(\IncPC_Out<13> ), .D(n9), .Y(
        n154) );
  AOI22X1 U154 ( .A(\IncPC<12> ), .B(n19), .C(\IncPC_Out<12> ), .D(n9), .Y(
        n155) );
  AOI22X1 U155 ( .A(\IncPC<11> ), .B(n19), .C(\IncPC_Out<11> ), .D(n9), .Y(
        n156) );
  AOI22X1 U156 ( .A(\IncPC<10> ), .B(n19), .C(\IncPC_Out<10> ), .D(n9), .Y(
        n157) );
  AOI22X1 U157 ( .A(\IncPC<0> ), .B(n19), .C(\IncPC_Out<0> ), .D(n9), .Y(n158)
         );
  AOI22X1 U158 ( .A(\Immediate<9> ), .B(n19), .C(\Immediate_Out<9> ), .D(n9), 
        .Y(n159) );
  AOI22X1 U159 ( .A(\Immediate<8> ), .B(n19), .C(\Immediate_Out<8> ), .D(n9), 
        .Y(n160) );
  AOI22X1 U160 ( .A(\Immediate<7> ), .B(n19), .C(\Immediate_Out<7> ), .D(n9), 
        .Y(n161) );
  AOI22X1 U161 ( .A(\Immediate<6> ), .B(n20), .C(\Immediate_Out<6> ), .D(n9), 
        .Y(n162) );
  AOI22X1 U162 ( .A(\Immediate<5> ), .B(n20), .C(\Immediate_Out<5> ), .D(n9), 
        .Y(n163) );
  AOI22X1 U163 ( .A(\Immediate<4> ), .B(n20), .C(\Immediate_Out<4> ), .D(n9), 
        .Y(n164) );
  AOI22X1 U164 ( .A(\Immediate<3> ), .B(n20), .C(\Immediate_Out<3> ), .D(n9), 
        .Y(n165) );
  AOI22X1 U165 ( .A(\Immediate<2> ), .B(n20), .C(\Immediate_Out<2> ), .D(n10), 
        .Y(n166) );
  AOI22X1 U166 ( .A(\Immediate<1> ), .B(n20), .C(\Immediate_Out<1> ), .D(n10), 
        .Y(n167) );
  AOI22X1 U167 ( .A(\Immediate<15> ), .B(n20), .C(\Immediate_Out<15> ), .D(n10), .Y(n168) );
  AOI22X1 U168 ( .A(\Immediate<14> ), .B(n20), .C(\Immediate_Out<14> ), .D(n10), .Y(n169) );
  AOI22X1 U169 ( .A(\Immediate<13> ), .B(n20), .C(\Immediate_Out<13> ), .D(n10), .Y(n170) );
  AOI22X1 U170 ( .A(\Immediate<12> ), .B(n20), .C(\Immediate_Out<12> ), .D(n10), .Y(n171) );
  AOI22X1 U171 ( .A(\Immediate<11> ), .B(n20), .C(\Immediate_Out<11> ), .D(n10), .Y(n172) );
  AOI22X1 U172 ( .A(\Immediate<10> ), .B(n21), .C(\Immediate_Out<10> ), .D(n10), .Y(n173) );
  AOI22X1 U173 ( .A(\Immediate<0> ), .B(n21), .C(\Immediate_Out<0> ), .D(n10), 
        .Y(n174) );
  AOI22X1 U174 ( .A(Halt), .B(n21), .C(Halt_Out), .D(n10), .Y(n175) );
  AOI22X1 U175 ( .A(\Func<1> ), .B(n21), .C(\Func_Out<1> ), .D(n10), .Y(n176)
         );
  AOI22X1 U176 ( .A(\Func<0> ), .B(n21), .C(\Func_Out<0> ), .D(n10), .Y(n177)
         );
  AOI22X1 U177 ( .A(\DecodeIncPC<9> ), .B(n21), .C(\DecodeIncPC_Out<9> ), .D(
        n11), .Y(n178) );
  AOI22X1 U178 ( .A(\DecodeIncPC<8> ), .B(n21), .C(\DecodeIncPC_Out<8> ), .D(
        n11), .Y(n179) );
  AOI22X1 U179 ( .A(\DecodeIncPC<7> ), .B(n21), .C(\DecodeIncPC_Out<7> ), .D(
        n11), .Y(n180) );
  AOI22X1 U180 ( .A(\DecodeIncPC<6> ), .B(n21), .C(\DecodeIncPC_Out<6> ), .D(
        n11), .Y(n181) );
  AOI22X1 U181 ( .A(\DecodeIncPC<5> ), .B(n21), .C(\DecodeIncPC_Out<5> ), .D(
        n11), .Y(n182) );
  AOI22X1 U182 ( .A(\DecodeIncPC<4> ), .B(n21), .C(\DecodeIncPC_Out<4> ), .D(
        n11), .Y(n183) );
  AOI22X1 U183 ( .A(\DecodeIncPC<3> ), .B(n22), .C(\DecodeIncPC_Out<3> ), .D(
        n11), .Y(n184) );
  AOI22X1 U184 ( .A(\DecodeIncPC<2> ), .B(n22), .C(\DecodeIncPC_Out<2> ), .D(
        n11), .Y(n185) );
  AOI22X1 U185 ( .A(\DecodeIncPC<1> ), .B(n22), .C(\DecodeIncPC_Out<1> ), .D(
        n11), .Y(n186) );
  AOI22X1 U186 ( .A(\DecodeIncPC<15> ), .B(n22), .C(\DecodeIncPC_Out<15> ), 
        .D(n11), .Y(n187) );
  AOI22X1 U187 ( .A(\DecodeIncPC<14> ), .B(n22), .C(\DecodeIncPC_Out<14> ), 
        .D(n11), .Y(n188) );
  AOI22X1 U188 ( .A(\DecodeIncPC<13> ), .B(n22), .C(\DecodeIncPC_Out<13> ), 
        .D(n11), .Y(n189) );
  AOI22X1 U189 ( .A(\DecodeIncPC<12> ), .B(n22), .C(\DecodeIncPC_Out<12> ), 
        .D(n12), .Y(n190) );
  AOI22X1 U190 ( .A(\DecodeIncPC<11> ), .B(n22), .C(\DecodeIncPC_Out<11> ), 
        .D(n12), .Y(n191) );
  AOI22X1 U191 ( .A(\DecodeIncPC<10> ), .B(n22), .C(\DecodeIncPC_Out<10> ), 
        .D(n12), .Y(n192) );
  AOI22X1 U192 ( .A(\DecodeIncPC<0> ), .B(n22), .C(n1), .D(n12), .Y(n193) );
  AOI22X1 U193 ( .A(Cin), .B(n22), .C(Cin_Out), .D(n12), .Y(n194) );
  AOI22X1 U194 ( .A(Btr), .B(n23), .C(Btr_Out), .D(n12), .Y(n195) );
  AOI22X1 U195 ( .A(Branch), .B(n23), .C(Branch_Out), .D(n12), .Y(n196) );
  AOI22X1 U196 ( .A(ALUSrc), .B(n23), .C(ALUSrc_Out), .D(n12), .Y(n197) );
  AOI22X1 U197 ( .A(\ALUOpcode<2> ), .B(n23), .C(\ALUOpcode_Out<2> ), .D(n12), 
        .Y(n198) );
  AOI22X1 U198 ( .A(\ALUOpcode<1> ), .B(n23), .C(\ALUOpcode_Out<1> ), .D(n12), 
        .Y(n199) );
  AOI22X1 U199 ( .A(\ALUOpcode<0> ), .B(n23), .C(n2), .D(n12), .Y(n200) );
  AOI22X1 U200 ( .A(\ALUOp2<9> ), .B(n23), .C(\ALUOp2_Out<9> ), .D(n12), .Y(
        n201) );
  AOI22X1 U201 ( .A(\ALUOp2<8> ), .B(n23), .C(\ALUOp2_Out<8> ), .D(n13), .Y(
        n202) );
  AOI22X1 U202 ( .A(\ALUOp2<7> ), .B(n23), .C(\ALUOp2_Out<7> ), .D(n13), .Y(
        n203) );
  AOI22X1 U203 ( .A(\ALUOp2<6> ), .B(n23), .C(\ALUOp2_Out<6> ), .D(n13), .Y(
        n204) );
  AOI22X1 U204 ( .A(\ALUOp2<5> ), .B(n23), .C(\ALUOp2_Out<5> ), .D(n13), .Y(
        n205) );
  AOI22X1 U205 ( .A(\ALUOp2<4> ), .B(n24), .C(\ALUOp2_Out<4> ), .D(n13), .Y(
        n206) );
  AOI22X1 U206 ( .A(\ALUOp2<3> ), .B(n24), .C(\ALUOp2_Out<3> ), .D(n13), .Y(
        n207) );
  AOI22X1 U207 ( .A(\ALUOp2<2> ), .B(n24), .C(\ALUOp2_Out<2> ), .D(n13), .Y(
        n208) );
  AOI22X1 U208 ( .A(\ALUOp2<1> ), .B(n24), .C(\ALUOp2_Out<1> ), .D(n13), .Y(
        n209) );
  AOI22X1 U209 ( .A(\ALUOp2<15> ), .B(n24), .C(\ALUOp2_Out<15> ), .D(n13), .Y(
        n210) );
  AOI22X1 U210 ( .A(\ALUOp2<14> ), .B(n24), .C(\ALUOp2_Out<14> ), .D(n13), .Y(
        n211) );
  AOI22X1 U211 ( .A(\ALUOp2<13> ), .B(n24), .C(\ALUOp2_Out<13> ), .D(n13), .Y(
        n212) );
  AOI22X1 U212 ( .A(\ALUOp2<12> ), .B(n24), .C(\ALUOp2_Out<12> ), .D(n13), .Y(
        n213) );
  AOI22X1 U213 ( .A(\ALUOp2<11> ), .B(n24), .C(\ALUOp2_Out<11> ), .D(n14), .Y(
        n214) );
  AOI22X1 U214 ( .A(\ALUOp2<10> ), .B(n24), .C(\ALUOp2_Out<10> ), .D(n14), .Y(
        n215) );
  AOI22X1 U215 ( .A(\ALUOp2<0> ), .B(n24), .C(\ALUOp2_Out<0> ), .D(n14), .Y(
        n216) );
  AOI22X1 U216 ( .A(\ALUOp1<9> ), .B(n25), .C(\ALUOp1_Out<9> ), .D(n14), .Y(
        n217) );
  AOI22X1 U217 ( .A(\ALUOp1<8> ), .B(n25), .C(\ALUOp1_Out<8> ), .D(n14), .Y(
        n218) );
  AOI22X1 U218 ( .A(\ALUOp1<7> ), .B(n25), .C(\ALUOp1_Out<7> ), .D(n14), .Y(
        n219) );
  AOI22X1 U219 ( .A(\ALUOp1<6> ), .B(n25), .C(\ALUOp1_Out<6> ), .D(n14), .Y(
        n220) );
  AOI22X1 U220 ( .A(\ALUOp1<5> ), .B(n25), .C(\ALUOp1_Out<5> ), .D(n14), .Y(
        n221) );
  AOI22X1 U221 ( .A(\ALUOp1<4> ), .B(n25), .C(\ALUOp1_Out<4> ), .D(n14), .Y(
        n222) );
  AOI22X1 U222 ( .A(\ALUOp1<3> ), .B(n25), .C(\ALUOp1_Out<3> ), .D(n14), .Y(
        n223) );
  AOI22X1 U223 ( .A(\ALUOp1<2> ), .B(n25), .C(\ALUOp1_Out<2> ), .D(n14), .Y(
        n224) );
  AOI22X1 U224 ( .A(\ALUOp1<1> ), .B(n25), .C(\ALUOp1_Out<1> ), .D(n14), .Y(
        n225) );
  AOI22X1 U225 ( .A(\ALUOp1<15> ), .B(n25), .C(\ALUOp1_Out<15> ), .D(n15), .Y(
        n226) );
  AOI22X1 U226 ( .A(\ALUOp1<14> ), .B(n25), .C(\ALUOp1_Out<14> ), .D(n15), .Y(
        n227) );
  AOI22X1 U227 ( .A(\ALUOp1<13> ), .B(n26), .C(\ALUOp1_Out<13> ), .D(n15), .Y(
        n228) );
  AOI22X1 U228 ( .A(\ALUOp1<12> ), .B(n26), .C(\ALUOp1_Out<12> ), .D(n15), .Y(
        n229) );
  AOI22X1 U229 ( .A(\ALUOp1<11> ), .B(n26), .C(\ALUOp1_Out<11> ), .D(n15), .Y(
        n230) );
  AOI22X1 U230 ( .A(\ALUOp1<10> ), .B(n26), .C(\ALUOp1_Out<10> ), .D(n15), .Y(
        n231) );
  AOI22X1 U231 ( .A(\ALUOp1<0> ), .B(n26), .C(\ALUOp1_Out<0> ), .D(n15), .Y(
        n232) );
  dff_338 LinkReg ( .q(Link_Out), .d(n114), .clk(clk), .rst(n35) );
  dff_304 \DecodeIncPC_Reg[0]  ( .q(\DecodeIncPC_Out<0> ), .d(n116), .clk(clk), 
        .rst(n35) );
  dff_305 \DecodeIncPC_Reg[1]  ( .q(\DecodeIncPC_Out<1> ), .d(n117), .clk(clk), 
        .rst(n35) );
  dff_306 \DecodeIncPC_Reg[2]  ( .q(\DecodeIncPC_Out<2> ), .d(n233), .clk(clk), 
        .rst(n35) );
  dff_307 \DecodeIncPC_Reg[3]  ( .q(\DecodeIncPC_Out<3> ), .d(n234), .clk(clk), 
        .rst(n35) );
  dff_308 \DecodeIncPC_Reg[4]  ( .q(\DecodeIncPC_Out<4> ), .d(n235), .clk(clk), 
        .rst(n35) );
  dff_309 \DecodeIncPC_Reg[5]  ( .q(\DecodeIncPC_Out<5> ), .d(n236), .clk(clk), 
        .rst(n35) );
  dff_310 \DecodeIncPC_Reg[6]  ( .q(\DecodeIncPC_Out<6> ), .d(n237), .clk(clk), 
        .rst(n35) );
  dff_311 \DecodeIncPC_Reg[7]  ( .q(\DecodeIncPC_Out<7> ), .d(n238), .clk(clk), 
        .rst(n35) );
  dff_312 \DecodeIncPC_Reg[8]  ( .q(\DecodeIncPC_Out<8> ), .d(n239), .clk(clk), 
        .rst(n35) );
  dff_313 \DecodeIncPC_Reg[9]  ( .q(\DecodeIncPC_Out<9> ), .d(n240), .clk(clk), 
        .rst(n35) );
  dff_314 \DecodeIncPC_Reg[10]  ( .q(\DecodeIncPC_Out<10> ), .d(n241), .clk(
        clk), .rst(n35) );
  dff_315 \DecodeIncPC_Reg[11]  ( .q(\DecodeIncPC_Out<11> ), .d(n242), .clk(
        clk), .rst(n34) );
  dff_316 \DecodeIncPC_Reg[12]  ( .q(\DecodeIncPC_Out<12> ), .d(n243), .clk(
        clk), .rst(n34) );
  dff_317 \DecodeIncPC_Reg[13]  ( .q(\DecodeIncPC_Out<13> ), .d(n244), .clk(
        clk), .rst(n34) );
  dff_318 \DecodeIncPC_Reg[14]  ( .q(\DecodeIncPC_Out<14> ), .d(n245), .clk(
        clk), .rst(n34) );
  dff_319 \DecodeIncPC_Reg[15]  ( .q(\DecodeIncPC_Out<15> ), .d(n246), .clk(
        clk), .rst(n34) );
  dff_337 RtValid_reg ( .q(RtValid_Out), .d(n64), .clk(clk), .rst(n34) );
  dff_336 RsValid_reg ( .q(RsValid_Out), .d(n111), .clk(clk), .rst(n34) );
  dff_335 RdValid_reg ( .q(RdValid_Out), .d(n112), .clk(clk), .rst(n34) );
  dff_301 \WriteReg_reg[0]  ( .q(\WriteReg_Out<0> ), .d(n247), .clk(clk), 
        .rst(n34) );
  dff_302 \WriteReg_reg[1]  ( .q(\WriteReg_Out<1> ), .d(n248), .clk(clk), 
        .rst(n34) );
  dff_303 \WriteReg_reg[2]  ( .q(\WriteReg_Out<2> ), .d(n249), .clk(clk), 
        .rst(n34) );
  dff_285 \incpc_reg[0]  ( .q(\IncPC_Out<0> ), .d(n250), .clk(clk), .rst(n34)
         );
  dff_286 \incpc_reg[1]  ( .q(\IncPC_Out<1> ), .d(n51), .clk(clk), .rst(n34)
         );
  dff_287 \incpc_reg[2]  ( .q(\IncPC_Out<2> ), .d(n49), .clk(clk), .rst(n33)
         );
  dff_288 \incpc_reg[3]  ( .q(\IncPC_Out<3> ), .d(n50), .clk(clk), .rst(n33)
         );
  dff_289 \incpc_reg[4]  ( .q(\IncPC_Out<4> ), .d(n37), .clk(clk), .rst(n33)
         );
  dff_290 \incpc_reg[5]  ( .q(\IncPC_Out<5> ), .d(n38), .clk(clk), .rst(n33)
         );
  dff_291 \incpc_reg[6]  ( .q(\IncPC_Out<6> ), .d(n39), .clk(clk), .rst(n33)
         );
  dff_292 \incpc_reg[7]  ( .q(\IncPC_Out<7> ), .d(n40), .clk(clk), .rst(n33)
         );
  dff_293 \incpc_reg[8]  ( .q(\IncPC_Out<8> ), .d(n41), .clk(clk), .rst(n33)
         );
  dff_294 \incpc_reg[9]  ( .q(\IncPC_Out<9> ), .d(n42), .clk(clk), .rst(n33)
         );
  dff_295 \incpc_reg[10]  ( .q(\IncPC_Out<10> ), .d(n43), .clk(clk), .rst(n33)
         );
  dff_296 \incpc_reg[11]  ( .q(\IncPC_Out<11> ), .d(n44), .clk(clk), .rst(n33)
         );
  dff_297 \incpc_reg[12]  ( .q(\IncPC_Out<12> ), .d(n45), .clk(clk), .rst(n33)
         );
  dff_298 \incpc_reg[13]  ( .q(\IncPC_Out<13> ), .d(n46), .clk(clk), .rst(n33)
         );
  dff_299 \incpc_reg[14]  ( .q(\IncPC_Out<14> ), .d(n47), .clk(clk), .rst(n33)
         );
  dff_300 \incpc_reg[15]  ( .q(\IncPC_Out<15> ), .d(n48), .clk(clk), .rst(n32)
         );
  dff_334 rf_wr_en_reg ( .q(RegFileWrEn_Out), .d(n63), .clk(clk), .rst(n32) );
  dff_282 \rs_reg[0]  ( .q(\Rs_Out<0> ), .d(n108), .clk(clk), .rst(n32) );
  dff_283 \rs_reg[1]  ( .q(\Rs_Out<1> ), .d(n109), .clk(clk), .rst(n32) );
  dff_284 \rs_reg[2]  ( .q(\Rs_Out<2> ), .d(n110), .clk(clk), .rst(n32) );
  dff_279 \rt_reg[0]  ( .q(\Rt_Out<0> ), .d(n89), .clk(clk), .rst(n32) );
  dff_280 \rt_reg[1]  ( .q(\Rt_Out<1> ), .d(n90), .clk(clk), .rst(n32) );
  dff_281 \rt_reg[2]  ( .q(\Rt_Out<2> ), .d(n91), .clk(clk), .rst(n32) );
  dff_276 \rd_reg[0]  ( .q(\Rd_Out<0> ), .d(n57), .clk(clk), .rst(n32) );
  dff_277 \rd_reg[1]  ( .q(\Rd_Out<1> ), .d(n71), .clk(clk), .rst(n32) );
  dff_278 \rd_reg[2]  ( .q(\Rd_Out<2> ), .d(n72), .clk(clk), .rst(n32) );
  dff_260 \ALUOp1_reg[0]  ( .q(\ALUOp1_Out<0> ), .d(n93), .clk(clk), .rst(n32)
         );
  dff_261 \ALUOp1_reg[1]  ( .q(\ALUOp1_Out<1> ), .d(n101), .clk(clk), .rst(n32) );
  dff_262 \ALUOp1_reg[2]  ( .q(\ALUOp1_Out<2> ), .d(n102), .clk(clk), .rst(n31) );
  dff_263 \ALUOp1_reg[3]  ( .q(\ALUOp1_Out<3> ), .d(n103), .clk(clk), .rst(n31) );
  dff_264 \ALUOp1_reg[4]  ( .q(\ALUOp1_Out<4> ), .d(n104), .clk(clk), .rst(n31) );
  dff_265 \ALUOp1_reg[5]  ( .q(\ALUOp1_Out<5> ), .d(n105), .clk(clk), .rst(n31) );
  dff_266 \ALUOp1_reg[6]  ( .q(\ALUOp1_Out<6> ), .d(n106), .clk(clk), .rst(n31) );
  dff_267 \ALUOp1_reg[7]  ( .q(\ALUOp1_Out<7> ), .d(n107), .clk(clk), .rst(n31) );
  dff_268 \ALUOp1_reg[8]  ( .q(\ALUOp1_Out<8> ), .d(n92), .clk(clk), .rst(n31)
         );
  dff_269 \ALUOp1_reg[9]  ( .q(\ALUOp1_Out<9> ), .d(n100), .clk(clk), .rst(n31) );
  dff_270 \ALUOp1_reg[10]  ( .q(\ALUOp1_Out<10> ), .d(n94), .clk(clk), .rst(
        n31) );
  dff_271 \ALUOp1_reg[11]  ( .q(\ALUOp1_Out<11> ), .d(n95), .clk(clk), .rst(
        n31) );
  dff_272 \ALUOp1_reg[12]  ( .q(\ALUOp1_Out<12> ), .d(n96), .clk(clk), .rst(
        n31) );
  dff_273 \ALUOp1_reg[13]  ( .q(\ALUOp1_Out<13> ), .d(n97), .clk(clk), .rst(
        n31) );
  dff_274 \ALUOp1_reg[14]  ( .q(\ALUOp1_Out<14> ), .d(n98), .clk(clk), .rst(
        n31) );
  dff_275 \ALUOp1_reg[15]  ( .q(\ALUOp1_Out<15> ), .d(n99), .clk(clk), .rst(
        n30) );
  dff_244 \ALUOp2_reg[0]  ( .q(\ALUOp2_Out<0> ), .d(n73), .clk(clk), .rst(n30)
         );
  dff_245 \ALUOp2_reg[1]  ( .q(\ALUOp2_Out<1> ), .d(n80), .clk(clk), .rst(n30)
         );
  dff_246 \ALUOp2_reg[2]  ( .q(\ALUOp2_Out<2> ), .d(n81), .clk(clk), .rst(n30)
         );
  dff_247 \ALUOp2_reg[3]  ( .q(\ALUOp2_Out<3> ), .d(n82), .clk(clk), .rst(n30)
         );
  dff_248 \ALUOp2_reg[4]  ( .q(\ALUOp2_Out<4> ), .d(n83), .clk(clk), .rst(n30)
         );
  dff_249 \ALUOp2_reg[5]  ( .q(\ALUOp2_Out<5> ), .d(n84), .clk(clk), .rst(n30)
         );
  dff_250 \ALUOp2_reg[6]  ( .q(\ALUOp2_Out<6> ), .d(n85), .clk(clk), .rst(n30)
         );
  dff_251 \ALUOp2_reg[7]  ( .q(\ALUOp2_Out<7> ), .d(n86), .clk(clk), .rst(n30)
         );
  dff_252 \ALUOp2_reg[8]  ( .q(\ALUOp2_Out<8> ), .d(n87), .clk(clk), .rst(n30)
         );
  dff_253 \ALUOp2_reg[9]  ( .q(\ALUOp2_Out<9> ), .d(n88), .clk(clk), .rst(n30)
         );
  dff_254 \ALUOp2_reg[10]  ( .q(\ALUOp2_Out<10> ), .d(n74), .clk(clk), .rst(
        n30) );
  dff_255 \ALUOp2_reg[11]  ( .q(\ALUOp2_Out<11> ), .d(n75), .clk(clk), .rst(
        n30) );
  dff_256 \ALUOp2_reg[12]  ( .q(\ALUOp2_Out<12> ), .d(n76), .clk(clk), .rst(
        n29) );
  dff_257 \ALUOp2_reg[13]  ( .q(\ALUOp2_Out<13> ), .d(n77), .clk(clk), .rst(
        n29) );
  dff_258 \ALUOp2_reg[14]  ( .q(\ALUOp2_Out<14> ), .d(n78), .clk(clk), .rst(
        n29) );
  dff_259 \ALUOp2_reg[15]  ( .q(\ALUOp2_Out<15> ), .d(n79), .clk(clk), .rst(
        n29) );
  dff_228 \Immediate_reg[0]  ( .q(\Immediate_Out<0> ), .d(n251), .clk(clk), 
        .rst(n29) );
  dff_229 \Immediate_reg[1]  ( .q(\Immediate_Out<1> ), .d(n252), .clk(clk), 
        .rst(n29) );
  dff_230 \Immediate_reg[2]  ( .q(\Immediate_Out<2> ), .d(n253), .clk(clk), 
        .rst(n29) );
  dff_231 \Immediate_reg[3]  ( .q(\Immediate_Out<3> ), .d(n254), .clk(clk), 
        .rst(n29) );
  dff_232 \Immediate_reg[4]  ( .q(\Immediate_Out<4> ), .d(n255), .clk(clk), 
        .rst(n29) );
  dff_233 \Immediate_reg[5]  ( .q(\Immediate_Out<5> ), .d(n256), .clk(clk), 
        .rst(n29) );
  dff_234 \Immediate_reg[6]  ( .q(\Immediate_Out<6> ), .d(n257), .clk(clk), 
        .rst(n29) );
  dff_235 \Immediate_reg[7]  ( .q(\Immediate_Out<7> ), .d(n258), .clk(clk), 
        .rst(n29) );
  dff_236 \Immediate_reg[8]  ( .q(\Immediate_Out<8> ), .d(n259), .clk(clk), 
        .rst(n29) );
  dff_237 \Immediate_reg[9]  ( .q(\Immediate_Out<9> ), .d(n260), .clk(clk), 
        .rst(n28) );
  dff_238 \Immediate_reg[10]  ( .q(\Immediate_Out<10> ), .d(n261), .clk(clk), 
        .rst(n28) );
  dff_239 \Immediate_reg[11]  ( .q(\Immediate_Out<11> ), .d(n262), .clk(clk), 
        .rst(n28) );
  dff_240 \Immediate_reg[12]  ( .q(\Immediate_Out<12> ), .d(n263), .clk(clk), 
        .rst(n28) );
  dff_241 \Immediate_reg[13]  ( .q(\Immediate_Out<13> ), .d(n264), .clk(clk), 
        .rst(n28) );
  dff_242 \Immediate_reg[14]  ( .q(\Immediate_Out<14> ), .d(n265), .clk(clk), 
        .rst(n28) );
  dff_243 \Immediate_reg[15]  ( .q(\Immediate_Out<15> ), .d(n266), .clk(clk), 
        .rst(n28) );
  dff_225 \ALUOpcode_reg[0]  ( .q(\ALUOpcode_Out<0> ), .d(n52), .clk(clk), 
        .rst(n28) );
  dff_226 \ALUOpcode_reg[1]  ( .q(\ALUOpcode_Out<1> ), .d(n56), .clk(clk), 
        .rst(n28) );
  dff_227 \ALUOpcode_reg[2]  ( .q(\ALUOpcode_Out<2> ), .d(n113), .clk(clk), 
        .rst(n28) );
  dff_223 \Func_reg[0]  ( .q(\Func_Out<0> ), .d(n62), .clk(clk), .rst(n28) );
  dff_224 \Func_reg[1]  ( .q(\Func_Out<1> ), .d(n115), .clk(clk), .rst(n28) );
  dff_333 ALUSrc_reg ( .q(ALUSrc_Out), .d(n61), .clk(clk), .rst(n28) );
  dff_332 Branch_reg ( .q(Branch_Out), .d(n60), .clk(clk), .rst(n27) );
  dff_331 Jump_reg ( .q(Jump_Out), .d(n59), .clk(clk), .rst(n27) );
  dff_330 JumpReg_reg ( .q(JumpReg_Out), .d(n58), .clk(clk), .rst(n27) );
  dff_329 Set_reg ( .q(Set_Out), .d(n69), .clk(clk), .rst(n27) );
  dff_328 Btr_reg ( .q(Btr_Out), .d(n68), .clk(clk), .rst(n27) );
  dff_327 MemWrite_reg ( .q(MemWrite_Out), .d(n67), .clk(clk), .rst(n27) );
  dff_326 MemRead_reg ( .q(MemRead_Out), .d(n66), .clk(clk), .rst(n27) );
  dff_325 MemToReg_reg ( .q(MemToReg_Out), .d(n65), .clk(clk), .rst(n27) );
  dff_324 Halt_reg ( .q(Halt_Out), .d(n70), .clk(clk), .rst(n27) );
  dff_323 InvA_reg ( .q(InvA_Out), .d(n54), .clk(clk), .rst(n27) );
  dff_322 InvB_reg ( .q(InvB_Out), .d(n53), .clk(clk), .rst(n27) );
  dff_321 Cin_reg ( .q(Cin_Out), .d(n55), .clk(clk), .rst(n27) );
  dff_320 CPUActive_reg ( .q(CPUActive_Out), .d(CPUActive), .clk(clk), .rst(
        n27) );
  INVX1 U1 ( .A(n16), .Y(n15) );
  INVX1 U2 ( .A(n16), .Y(n14) );
  INVX1 U3 ( .A(n5), .Y(n23) );
  INVX1 U4 ( .A(n232), .Y(n93) );
  INVX1 U5 ( .A(n225), .Y(n101) );
  INVX1 U6 ( .A(n137), .Y(n66) );
  INVX1 U7 ( .A(n16), .Y(n13) );
  INVX1 U8 ( .A(n130), .Y(n63) );
  INVX1 U9 ( .A(n224), .Y(n102) );
  INVX1 U10 ( .A(n223), .Y(n103) );
  INVX1 U11 ( .A(n222), .Y(n104) );
  INVX1 U12 ( .A(n221), .Y(n105) );
  INVX1 U13 ( .A(n220), .Y(n106) );
  INVX1 U14 ( .A(n219), .Y(n107) );
  INVX1 U15 ( .A(n177), .Y(n62) );
  INVX1 U16 ( .A(n139), .Y(n59) );
  INVX1 U17 ( .A(n140), .Y(n58) );
  INVX1 U18 ( .A(n121), .Y(n69) );
  INVX1 U19 ( .A(n195), .Y(n68) );
  INVX1 U20 ( .A(n136), .Y(n65) );
  INVX1 U21 ( .A(n142), .Y(n54) );
  INVX1 U22 ( .A(n141), .Y(n53) );
  INVX1 U23 ( .A(n194), .Y(n55) );
  INVX1 U24 ( .A(n5), .Y(n24) );
  INVX1 U25 ( .A(n17), .Y(n5) );
  INVX1 U26 ( .A(n10), .Y(n25) );
  INVX1 U27 ( .A(rst), .Y(n36) );
  INVX1 U28 ( .A(Stall), .Y(n17) );
  INVX1 U29 ( .A(n5), .Y(n18) );
  INVX1 U30 ( .A(n5), .Y(n26) );
  BUFX2 U31 ( .A(\DecodeIncPC_Out<0> ), .Y(n1) );
  INVX1 U32 ( .A(n125), .Y(n64) );
  INVX1 U33 ( .A(n36), .Y(n27) );
  INVX1 U34 ( .A(n36), .Y(n28) );
  INVX1 U35 ( .A(n36), .Y(n29) );
  INVX1 U36 ( .A(n36), .Y(n30) );
  INVX1 U37 ( .A(n36), .Y(n31) );
  INVX1 U38 ( .A(n36), .Y(n32) );
  INVX1 U39 ( .A(n36), .Y(n33) );
  INVX1 U40 ( .A(n36), .Y(n34) );
  INVX1 U41 ( .A(n36), .Y(n35) );
  INVX1 U42 ( .A(n231), .Y(n94) );
  INVX1 U43 ( .A(n230), .Y(n95) );
  INVX1 U44 ( .A(n229), .Y(n96) );
  INVX1 U45 ( .A(n228), .Y(n97) );
  INVX1 U46 ( .A(n227), .Y(n98) );
  INVX1 U47 ( .A(n226), .Y(n99) );
  INVX1 U48 ( .A(n218), .Y(n92) );
  INVX1 U49 ( .A(n217), .Y(n100) );
  INVX1 U50 ( .A(n216), .Y(n73) );
  INVX1 U51 ( .A(n215), .Y(n74) );
  INVX1 U52 ( .A(n214), .Y(n75) );
  INVX1 U53 ( .A(n213), .Y(n76) );
  INVX1 U54 ( .A(n212), .Y(n77) );
  INVX1 U55 ( .A(n211), .Y(n78) );
  INVX1 U56 ( .A(n210), .Y(n79) );
  INVX1 U57 ( .A(n209), .Y(n80) );
  INVX1 U58 ( .A(n208), .Y(n81) );
  INVX1 U59 ( .A(n207), .Y(n82) );
  INVX1 U60 ( .A(n206), .Y(n83) );
  INVX1 U61 ( .A(n205), .Y(n84) );
  INVX1 U62 ( .A(n204), .Y(n85) );
  INVX1 U63 ( .A(n203), .Y(n86) );
  INVX1 U64 ( .A(n202), .Y(n87) );
  INVX1 U65 ( .A(n201), .Y(n88) );
  INVX1 U66 ( .A(n200), .Y(n52) );
  INVX1 U67 ( .A(n199), .Y(n56) );
  INVX1 U68 ( .A(n198), .Y(n113) );
  INVX1 U69 ( .A(n197), .Y(n61) );
  INVX1 U70 ( .A(n196), .Y(n60) );
  INVX1 U71 ( .A(n193), .Y(n116) );
  INVX1 U72 ( .A(n192), .Y(n241) );
  INVX1 U73 ( .A(n191), .Y(n242) );
  INVX1 U74 ( .A(n190), .Y(n243) );
  INVX1 U75 ( .A(n5), .Y(n22) );
  INVX1 U76 ( .A(n17), .Y(n12) );
  INVX1 U77 ( .A(n189), .Y(n244) );
  INVX1 U78 ( .A(n188), .Y(n245) );
  INVX1 U79 ( .A(n187), .Y(n246) );
  INVX1 U80 ( .A(n186), .Y(n117) );
  INVX1 U81 ( .A(n185), .Y(n233) );
  INVX1 U82 ( .A(n184), .Y(n234) );
  INVX1 U83 ( .A(n183), .Y(n235) );
  INVX1 U84 ( .A(n182), .Y(n236) );
  INVX1 U85 ( .A(n181), .Y(n237) );
  INVX1 U86 ( .A(n180), .Y(n238) );
  INVX1 U87 ( .A(n179), .Y(n239) );
  INVX1 U88 ( .A(n178), .Y(n240) );
  INVX1 U89 ( .A(n11), .Y(n21) );
  INVX1 U90 ( .A(n17), .Y(n11) );
  INVX1 U91 ( .A(n176), .Y(n115) );
  INVX1 U92 ( .A(n175), .Y(n70) );
  INVX1 U93 ( .A(n174), .Y(n251) );
  INVX1 U94 ( .A(n173), .Y(n261) );
  INVX1 U95 ( .A(n172), .Y(n262) );
  INVX1 U96 ( .A(n171), .Y(n263) );
  INVX1 U97 ( .A(n170), .Y(n264) );
  INVX1 U98 ( .A(n169), .Y(n265) );
  INVX1 U99 ( .A(n168), .Y(n266) );
  INVX1 U100 ( .A(n167), .Y(n252) );
  INVX1 U101 ( .A(n166), .Y(n253) );
  INVX1 U102 ( .A(n11), .Y(n20) );
  INVX1 U103 ( .A(n17), .Y(n10) );
  INVX1 U104 ( .A(n165), .Y(n254) );
  INVX1 U105 ( .A(n164), .Y(n255) );
  INVX1 U106 ( .A(n163), .Y(n256) );
  INVX1 U107 ( .A(n162), .Y(n257) );
  INVX1 U108 ( .A(n161), .Y(n258) );
  INVX1 U109 ( .A(n160), .Y(n259) );
  INVX1 U110 ( .A(n159), .Y(n260) );
  INVX1 U111 ( .A(n158), .Y(n250) );
  INVX1 U112 ( .A(n11), .Y(n19) );
  INVX1 U113 ( .A(n26), .Y(n9) );
  INVX1 U114 ( .A(n157), .Y(n43) );
  INVX1 U115 ( .A(n156), .Y(n44) );
  INVX1 U116 ( .A(n155), .Y(n45) );
  INVX1 U232 ( .A(n154), .Y(n46) );
  INVX1 U233 ( .A(n153), .Y(n47) );
  INVX1 U234 ( .A(n152), .Y(n48) );
  INVX1 U235 ( .A(n151), .Y(n51) );
  INVX1 U236 ( .A(n26), .Y(n8) );
  INVX1 U237 ( .A(n150), .Y(n49) );
  INVX1 U238 ( .A(n149), .Y(n50) );
  INVX1 U239 ( .A(n148), .Y(n37) );
  INVX1 U240 ( .A(n147), .Y(n38) );
  INVX1 U241 ( .A(n146), .Y(n39) );
  INVX1 U242 ( .A(n145), .Y(n40) );
  INVX1 U243 ( .A(n144), .Y(n41) );
  INVX1 U244 ( .A(n143), .Y(n42) );
  INVX1 U245 ( .A(n138), .Y(n114) );
  INVX1 U246 ( .A(n135), .Y(n67) );
  INVX1 U247 ( .A(n134), .Y(n112) );
  INVX1 U248 ( .A(n133), .Y(n57) );
  INVX1 U249 ( .A(n132), .Y(n71) );
  INVX1 U250 ( .A(n131), .Y(n72) );
  INVX1 U251 ( .A(n26), .Y(n7) );
  INVX1 U252 ( .A(n129), .Y(n111) );
  INVX1 U253 ( .A(n128), .Y(n108) );
  INVX1 U254 ( .A(n127), .Y(n109) );
  INVX1 U255 ( .A(n126), .Y(n110) );
  INVX1 U256 ( .A(n124), .Y(n89) );
  INVX1 U257 ( .A(n123), .Y(n90) );
  INVX1 U258 ( .A(n122), .Y(n91) );
  INVX1 U259 ( .A(n120), .Y(n247) );
  INVX1 U260 ( .A(n119), .Y(n248) );
  INVX1 U261 ( .A(n118), .Y(n249) );
  INVX1 U262 ( .A(n12), .Y(n16) );
  INVX1 U263 ( .A(n17), .Y(n6) );
  BUFX2 U264 ( .A(\ALUOpcode_Out<0> ), .Y(n2) );
  BUFX2 U265 ( .A(Link_Out), .Y(n3) );
  BUFX2 U266 ( .A(JumpReg_Out), .Y(n4) );
endmodule


module execute ( .ALUOp1({\ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , 
        \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , 
        \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , 
        \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), .ALUOp2({\ALUOp2<15> , 
        \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , 
        \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , 
        \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), 
    .Opcode({\Opcode<2> , \Opcode<1> , \Opcode<0> }), .IncPC({\IncPC<15> , 
        \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , 
        \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , 
        \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> }), Jump, Branch, 
        JumpReg, Set, InvA, InvB, Cin, Btr, .Func({\Func<1> , \Func<0> }), 
    .Imm({\Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> , \Imm<11> , \Imm<10> , 
        \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> , \Imm<5> , \Imm<4> , \Imm<3> , 
        \Imm<2> , \Imm<1> , \Imm<0> }), ALUSrc, .Result({\Result<15> , 
        \Result<14> , \Result<13> , \Result<12> , \Result<11> , \Result<10> , 
        \Result<9> , \Result<8> , \Result<7> , \Result<6> , \Result<5> , 
        \Result<4> , \Result<3> , \Result<2> , \Result<1> , \Result<0> }), 
    .NextPC({\NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> , 
        \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> , 
        \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> , 
        \NextPC<1> , \NextPC<0> }), Err, BranchJumpTaken, rst, .DecodeIncPC({
        \DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> , 
        \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> , 
        \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> , \DecodeIncPC<6> , 
        \DecodeIncPC<5> , \DecodeIncPC<4> , \DecodeIncPC<3> , \DecodeIncPC<2> , 
        \DecodeIncPC<1> , \DecodeIncPC<0> }), Link, .ForwardALUOp1({
        \ForwardALUOp1<1> , \ForwardALUOp1<0> }), .ForwardALUOp2({
        \ForwardALUOp2<1> , \ForwardALUOp2<0> }), .PipeMW_Result({
        \PipeMW_Result<15> , \PipeMW_Result<14> , \PipeMW_Result<13> , 
        \PipeMW_Result<12> , \PipeMW_Result<11> , \PipeMW_Result<10> , 
        \PipeMW_Result<9> , \PipeMW_Result<8> , \PipeMW_Result<7> , 
        \PipeMW_Result<6> , \PipeMW_Result<5> , \PipeMW_Result<4> , 
        \PipeMW_Result<3> , \PipeMW_Result<2> , \PipeMW_Result<1> , 
        \PipeMW_Result<0> }), .PipeEM_Result({\PipeEM_Result<15> , 
        \PipeEM_Result<14> , \PipeEM_Result<13> , \PipeEM_Result<12> , 
        \PipeEM_Result<11> , \PipeEM_Result<10> , \PipeEM_Result<9> , 
        \PipeEM_Result<8> , \PipeEM_Result<7> , \PipeEM_Result<6> , 
        \PipeEM_Result<5> , \PipeEM_Result<4> , \PipeEM_Result<3> , 
        \PipeEM_Result<2> , \PipeEM_Result<1> , \PipeEM_Result<0> }) );
  input \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> ,
         \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> ,
         \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> ,
         \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , \Opcode<2> , \Opcode<1> , \Opcode<0> ,
         \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> ,
         \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> ,
         \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> ,
         \IncPC<0> , Jump, Branch, JumpReg, Set, InvA, InvB, Cin, Btr,
         \Func<1> , \Func<0> , \Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> ,
         \Imm<11> , \Imm<10> , \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> ,
         \Imm<5> , \Imm<4> , \Imm<3> , \Imm<2> , \Imm<1> , \Imm<0> , ALUSrc,
         rst, \DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> ,
         \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> ,
         \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> ,
         \DecodeIncPC<6> , \DecodeIncPC<5> , \DecodeIncPC<4> ,
         \DecodeIncPC<3> , \DecodeIncPC<2> , \DecodeIncPC<1> ,
         \DecodeIncPC<0> , Link, \ForwardALUOp1<1> , \ForwardALUOp1<0> ,
         \ForwardALUOp2<1> , \ForwardALUOp2<0> , \PipeMW_Result<15> ,
         \PipeMW_Result<14> , \PipeMW_Result<13> , \PipeMW_Result<12> ,
         \PipeMW_Result<11> , \PipeMW_Result<10> , \PipeMW_Result<9> ,
         \PipeMW_Result<8> , \PipeMW_Result<7> , \PipeMW_Result<6> ,
         \PipeMW_Result<5> , \PipeMW_Result<4> , \PipeMW_Result<3> ,
         \PipeMW_Result<2> , \PipeMW_Result<1> , \PipeMW_Result<0> ,
         \PipeEM_Result<15> , \PipeEM_Result<14> , \PipeEM_Result<13> ,
         \PipeEM_Result<12> , \PipeEM_Result<11> , \PipeEM_Result<10> ,
         \PipeEM_Result<9> , \PipeEM_Result<8> , \PipeEM_Result<7> ,
         \PipeEM_Result<6> , \PipeEM_Result<5> , \PipeEM_Result<4> ,
         \PipeEM_Result<3> , \PipeEM_Result<2> , \PipeEM_Result<1> ,
         \PipeEM_Result<0> ;
  output \Result<15> , \Result<14> , \Result<13> , \Result<12> , \Result<11> ,
         \Result<10> , \Result<9> , \Result<8> , \Result<7> , \Result<6> ,
         \Result<5> , \Result<4> , \Result<3> , \Result<2> , \Result<1> ,
         \Result<0> , \NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> ,
         \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> ,
         \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> ,
         \NextPC<1> , \NextPC<0> , Err, BranchJumpTaken;
  wire   n514, n515, n516, n517, n518, n519, \alu_operand_a<10> ,
         \alu_operand_a<0> , \alu_operand_b<15> , \alu_operand_b<14> ,
         \alu_operand_b<11> , \aluResult<15> , \aluResult<14> ,
         \aluResult<13> , \aluResult<12> , \aluResult<11> , \aluResult<10> ,
         \aluResult<9> , \aluResult<8> , \aluResult<7> , \aluResult<6> ,
         \aluResult<5> , \aluResult<4> , \aluResult<3> , \aluResult<2> ,
         \aluResult<1> , \aluResult<0> , Zero, cout, \OpAReg<15> ,
         \OpAReg<14> , \OpAReg<13> , \OpAReg<12> , \OpAReg<11> , \OpAReg<10> ,
         \OpAReg<9> , \OpAReg<8> , \OpAReg<7> , \OpAReg<6> , \OpAReg<5> ,
         \OpAReg<4> , \OpAReg<3> , \OpAReg<2> , \OpAReg<1> , \OpAReg<0> ,
         \OpBReg<15> , \OpBReg<14> , \OpBReg<13> , \OpBReg<12> , \OpBReg<11> ,
         \OpBReg<10> , \OpBReg<9> , \OpBReg<8> , \OpBReg<7> , \OpBReg<6> ,
         \OpBReg<5> , \OpBReg<4> , \OpBReg<3> , \OpBReg<2> , \OpBReg<1> ,
         \OpBReg<0> , N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N54, \_2_net_<0> , \setResult<15> ,
         \setResult<14> , \setResult<13> , \setResult<12> , \setResult<11> ,
         \setResult<10> , \setResult<9> , \setResult<8> , \setResult<7> ,
         \setResult<6> , \setResult<5> , \setResult<4> , \setResult<3> ,
         \setResult<2> , \setResult<1> , \setResult<0> , \offsetAddr<15> ,
         \offsetAddr<14> , \offsetAddr<13> , \offsetAddr<12> ,
         \offsetAddr<11> , \offsetAddr<10> , \offsetAddr<9> , \offsetAddr<8> ,
         \offsetAddr<7> , \offsetAddr<6> , \offsetAddr<5> , \offsetAddr<4> ,
         \offsetAddr<3> , \offsetAddr<2> , \offsetAddr<1> , \offsetAddr<0> ,
         branch_en, _7_net_, n83, n84, n85, n86, n87, n88, n89, n90, n91, n113,
         n114, n146, n147, n148, n149, n150, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n185, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n137, n139, n141, n143, n145, n152, n184, n187, n204, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n217, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n306, n307, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513;
  assign Err = 1'b0;

  LATCH \OpAReg_reg<15>  ( .CLK(n300), .D(N54), .Q(\OpAReg<15> ) );
  LATCH \OpAReg_reg<14>  ( .CLK(n300), .D(N52), .Q(\OpAReg<14> ) );
  LATCH \OpAReg_reg<13>  ( .CLK(n300), .D(N51), .Q(\OpAReg<13> ) );
  LATCH \OpAReg_reg<12>  ( .CLK(n300), .D(N50), .Q(\OpAReg<12> ) );
  LATCH \OpAReg_reg<11>  ( .CLK(n300), .D(N49), .Q(\OpAReg<11> ) );
  LATCH \OpAReg_reg<10>  ( .CLK(n300), .D(N48), .Q(\OpAReg<10> ) );
  LATCH \OpAReg_reg<9>  ( .CLK(n300), .D(N47), .Q(\OpAReg<9> ) );
  LATCH \OpAReg_reg<8>  ( .CLK(n300), .D(N46), .Q(\OpAReg<8> ) );
  LATCH \OpAReg_reg<7>  ( .CLK(n300), .D(N45), .Q(\OpAReg<7> ) );
  LATCH \OpAReg_reg<6>  ( .CLK(n300), .D(N44), .Q(\OpAReg<6> ) );
  LATCH \OpAReg_reg<5>  ( .CLK(n300), .D(N43), .Q(\OpAReg<5> ) );
  LATCH \OpAReg_reg<4>  ( .CLK(n300), .D(N42), .Q(\OpAReg<4> ) );
  LATCH \OpAReg_reg<3>  ( .CLK(n300), .D(N41), .Q(\OpAReg<3> ) );
  LATCH \OpAReg_reg<2>  ( .CLK(n300), .D(N40), .Q(\OpAReg<2> ) );
  LATCH \OpAReg_reg<1>  ( .CLK(n300), .D(N39), .Q(\OpAReg<1> ) );
  LATCH \OpAReg_reg<0>  ( .CLK(n300), .D(N38), .Q(\OpAReg<0> ) );
  LATCH \OpBReg_reg<15>  ( .CLK(n302), .D(n299), .Q(\OpBReg<15> ) );
  LATCH \OpBReg_reg<14>  ( .CLK(n302), .D(n297), .Q(\OpBReg<14> ) );
  LATCH \OpBReg_reg<13>  ( .CLK(n302), .D(n295), .Q(\OpBReg<13> ) );
  LATCH \OpBReg_reg<12>  ( .CLK(n302), .D(n293), .Q(\OpBReg<12> ) );
  LATCH \OpBReg_reg<11>  ( .CLK(n302), .D(n291), .Q(\OpBReg<11> ) );
  LATCH \OpBReg_reg<10>  ( .CLK(n302), .D(n289), .Q(\OpBReg<10> ) );
  LATCH \OpBReg_reg<9>  ( .CLK(n302), .D(n287), .Q(\OpBReg<9> ) );
  LATCH \OpBReg_reg<8>  ( .CLK(n302), .D(n285), .Q(\OpBReg<8> ) );
  LATCH \OpBReg_reg<7>  ( .CLK(n302), .D(n283), .Q(\OpBReg<7> ) );
  LATCH \OpBReg_reg<6>  ( .CLK(n302), .D(n281), .Q(\OpBReg<6> ) );
  LATCH \OpBReg_reg<5>  ( .CLK(n302), .D(n279), .Q(\OpBReg<5> ) );
  LATCH \OpBReg_reg<4>  ( .CLK(n302), .D(n277), .Q(\OpBReg<4> ) );
  LATCH \OpBReg_reg<3>  ( .CLK(n302), .D(n275), .Q(\OpBReg<3> ) );
  LATCH \OpBReg_reg<2>  ( .CLK(n302), .D(n273), .Q(\OpBReg<2> ) );
  LATCH \OpBReg_reg<1>  ( .CLK(n302), .D(n271), .Q(\OpBReg<1> ) );
  LATCH \OpBReg_reg<0>  ( .CLK(n302), .D(n269), .Q(\OpBReg<0> ) );
  AND2X2 U20 ( .A(n503), .B(n502), .Y(n89) );
  NAND3X1 U120 ( .A(n83), .B(n84), .C(n85), .Y(_7_net_) );
  NOR3X1 U121 ( .A(n86), .B(n87), .C(n88), .Y(n85) );
  NAND2X1 U122 ( .A(n496), .B(n497), .Y(n88) );
  NAND2X1 U123 ( .A(n498), .B(n499), .Y(n87) );
  NAND3X1 U124 ( .A(n500), .B(n501), .C(n89), .Y(n86) );
  NOR3X1 U125 ( .A(n90), .B(\ALUOp1<1> ), .C(\ALUOp1<15> ), .Y(n84) );
  NAND2X1 U126 ( .A(n507), .B(n508), .Y(n90) );
  NOR3X1 U127 ( .A(n91), .B(\ALUOp1<10> ), .C(\ALUOp1<0> ), .Y(n83) );
  NAND2X1 U128 ( .A(n505), .B(n506), .Y(n91) );
  AOI22X1 U158 ( .A(\setResult<1> ), .B(n490), .C(\ALUOp1<14> ), .D(Btr), .Y(
        n113) );
  AOI22X1 U216 ( .A(n400), .B(\ALUOp2<15> ), .C(n150), .D(\Imm<15> ), .Y(n148)
         );
  AOI22X1 U217 ( .A(\PipeEM_Result<15> ), .B(n350), .C(\PipeMW_Result<15> ), 
        .D(n351), .Y(n147) );
  AOI22X1 U220 ( .A(\ALUOp2<14> ), .B(n400), .C(n150), .D(\Imm<14> ), .Y(n155)
         );
  AOI22X1 U221 ( .A(\PipeEM_Result<14> ), .B(n350), .C(\PipeMW_Result<14> ), 
        .D(n351), .Y(n154) );
  AOI22X1 U223 ( .A(\ALUOp2<13> ), .B(n400), .C(n150), .D(\Imm<13> ), .Y(n157)
         );
  AOI22X1 U224 ( .A(\PipeEM_Result<13> ), .B(n350), .C(\PipeMW_Result<13> ), 
        .D(n351), .Y(n156) );
  AOI22X1 U226 ( .A(\ALUOp2<12> ), .B(n400), .C(n150), .D(\Imm<12> ), .Y(n159)
         );
  AOI22X1 U227 ( .A(\PipeEM_Result<12> ), .B(n350), .C(\PipeMW_Result<12> ), 
        .D(n351), .Y(n158) );
  AOI22X1 U229 ( .A(\ALUOp2<11> ), .B(n400), .C(n150), .D(\Imm<11> ), .Y(n161)
         );
  AOI22X1 U230 ( .A(\PipeEM_Result<11> ), .B(n350), .C(\PipeMW_Result<11> ), 
        .D(n351), .Y(n160) );
  AOI22X1 U232 ( .A(\ALUOp2<10> ), .B(n400), .C(n150), .D(\Imm<10> ), .Y(n163)
         );
  AOI22X1 U233 ( .A(\PipeEM_Result<10> ), .B(n350), .C(\PipeMW_Result<10> ), 
        .D(n351), .Y(n162) );
  AOI22X1 U235 ( .A(\ALUOp2<9> ), .B(n400), .C(n150), .D(\Imm<9> ), .Y(n165)
         );
  AOI22X1 U236 ( .A(\PipeEM_Result<9> ), .B(n350), .C(\PipeMW_Result<9> ), .D(
        n351), .Y(n164) );
  AOI22X1 U238 ( .A(\ALUOp2<8> ), .B(n400), .C(n150), .D(\Imm<8> ), .Y(n167)
         );
  AOI22X1 U239 ( .A(\PipeEM_Result<8> ), .B(n350), .C(\PipeMW_Result<8> ), .D(
        n351), .Y(n166) );
  AOI22X1 U241 ( .A(\ALUOp2<7> ), .B(n400), .C(n150), .D(\Imm<7> ), .Y(n169)
         );
  AOI22X1 U242 ( .A(\PipeEM_Result<7> ), .B(n350), .C(\PipeMW_Result<7> ), .D(
        n351), .Y(n168) );
  AOI22X1 U244 ( .A(\ALUOp2<6> ), .B(n400), .C(n150), .D(\Imm<6> ), .Y(n171)
         );
  AOI22X1 U245 ( .A(\PipeEM_Result<6> ), .B(n350), .C(\PipeMW_Result<6> ), .D(
        n351), .Y(n170) );
  AOI22X1 U247 ( .A(\ALUOp2<5> ), .B(n400), .C(n150), .D(\Imm<5> ), .Y(n173)
         );
  AOI22X1 U248 ( .A(\PipeEM_Result<5> ), .B(n350), .C(\PipeMW_Result<5> ), .D(
        n351), .Y(n172) );
  AOI22X1 U250 ( .A(\ALUOp2<4> ), .B(n400), .C(n150), .D(\Imm<4> ), .Y(n175)
         );
  AOI22X1 U251 ( .A(\PipeEM_Result<4> ), .B(n350), .C(\PipeMW_Result<4> ), .D(
        n351), .Y(n174) );
  AOI22X1 U253 ( .A(\ALUOp2<3> ), .B(n400), .C(n150), .D(\Imm<3> ), .Y(n177)
         );
  AOI22X1 U254 ( .A(\PipeEM_Result<3> ), .B(n350), .C(\PipeMW_Result<3> ), .D(
        n351), .Y(n176) );
  AOI22X1 U256 ( .A(\ALUOp2<2> ), .B(n400), .C(n150), .D(\Imm<2> ), .Y(n179)
         );
  AOI22X1 U257 ( .A(\PipeEM_Result<2> ), .B(n350), .C(\PipeMW_Result<2> ), .D(
        n351), .Y(n178) );
  AOI22X1 U259 ( .A(\ALUOp2<1> ), .B(n400), .C(n150), .D(\Imm<1> ), .Y(n181)
         );
  AOI22X1 U260 ( .A(\PipeEM_Result<1> ), .B(n350), .C(\PipeMW_Result<1> ), .D(
        n351), .Y(n180) );
  AOI22X1 U262 ( .A(\ALUOp2<0> ), .B(n400), .C(n150), .D(\Imm<0> ), .Y(n183)
         );
  NOR2X1 U263 ( .A(n353), .B(ALUSrc), .Y(n149) );
  AOI22X1 U265 ( .A(\PipeEM_Result<0> ), .B(n350), .C(\PipeMW_Result<0> ), .D(
        n351), .Y(n182) );
  OAI21X1 U268 ( .A(n509), .B(n399), .C(n185), .Y(N54) );
  AOI22X1 U269 ( .A(n348), .B(\PipeEM_Result<15> ), .C(n349), .D(
        \PipeMW_Result<15> ), .Y(n185) );
  OAI21X1 U271 ( .A(n508), .B(n399), .C(n188), .Y(N52) );
  AOI22X1 U272 ( .A(n348), .B(\PipeEM_Result<14> ), .C(n349), .D(
        \PipeMW_Result<14> ), .Y(n188) );
  OAI21X1 U273 ( .A(n507), .B(n399), .C(n189), .Y(N51) );
  AOI22X1 U274 ( .A(n348), .B(\PipeEM_Result<13> ), .C(n349), .D(
        \PipeMW_Result<13> ), .Y(n189) );
  OAI21X1 U275 ( .A(n506), .B(n399), .C(n190), .Y(N50) );
  AOI22X1 U276 ( .A(n348), .B(\PipeEM_Result<12> ), .C(n349), .D(
        \PipeMW_Result<12> ), .Y(n190) );
  OAI21X1 U277 ( .A(n505), .B(n399), .C(n191), .Y(N49) );
  AOI22X1 U278 ( .A(n348), .B(\PipeEM_Result<11> ), .C(n349), .D(
        \PipeMW_Result<11> ), .Y(n191) );
  OAI21X1 U279 ( .A(n504), .B(n399), .C(n192), .Y(N48) );
  AOI22X1 U280 ( .A(n348), .B(\PipeEM_Result<10> ), .C(n349), .D(
        \PipeMW_Result<10> ), .Y(n192) );
  OAI21X1 U281 ( .A(n503), .B(n399), .C(n193), .Y(N47) );
  AOI22X1 U282 ( .A(n348), .B(\PipeEM_Result<9> ), .C(n349), .D(
        \PipeMW_Result<9> ), .Y(n193) );
  OAI21X1 U283 ( .A(n502), .B(n398), .C(n194), .Y(N46) );
  AOI22X1 U284 ( .A(n348), .B(\PipeEM_Result<8> ), .C(n349), .D(
        \PipeMW_Result<8> ), .Y(n194) );
  OAI21X1 U285 ( .A(n501), .B(n398), .C(n195), .Y(N45) );
  AOI22X1 U286 ( .A(n348), .B(\PipeEM_Result<7> ), .C(n349), .D(
        \PipeMW_Result<7> ), .Y(n195) );
  OAI21X1 U287 ( .A(n500), .B(n398), .C(n196), .Y(N44) );
  AOI22X1 U288 ( .A(n348), .B(\PipeEM_Result<6> ), .C(n349), .D(
        \PipeMW_Result<6> ), .Y(n196) );
  OAI21X1 U289 ( .A(n499), .B(n398), .C(n197), .Y(N43) );
  AOI22X1 U290 ( .A(n348), .B(\PipeEM_Result<5> ), .C(n349), .D(
        \PipeMW_Result<5> ), .Y(n197) );
  OAI21X1 U291 ( .A(n498), .B(n398), .C(n198), .Y(N42) );
  AOI22X1 U292 ( .A(n348), .B(\PipeEM_Result<4> ), .C(n349), .D(
        \PipeMW_Result<4> ), .Y(n198) );
  OAI21X1 U293 ( .A(n497), .B(n398), .C(n199), .Y(N41) );
  AOI22X1 U294 ( .A(n348), .B(\PipeEM_Result<3> ), .C(n349), .D(
        \PipeMW_Result<3> ), .Y(n199) );
  OAI21X1 U295 ( .A(n496), .B(n398), .C(n200), .Y(N40) );
  AOI22X1 U296 ( .A(n348), .B(\PipeEM_Result<2> ), .C(n349), .D(
        \PipeMW_Result<2> ), .Y(n200) );
  OAI21X1 U297 ( .A(n495), .B(n398), .C(n201), .Y(N39) );
  AOI22X1 U298 ( .A(n348), .B(\PipeEM_Result<1> ), .C(n349), .D(
        \PipeMW_Result<1> ), .Y(n201) );
  OAI21X1 U299 ( .A(n494), .B(n398), .C(n202), .Y(N38) );
  AOI22X1 U300 ( .A(n348), .B(\PipeEM_Result<0> ), .C(n349), .D(
        \PipeMW_Result<0> ), .Y(n202) );
  AOI21X1 U305 ( .A(branch_en), .B(Branch), .C(Jump), .Y(n146) );
  alu primary_alu ( .A({n214, n134, n132, n130, n342, \alu_operand_a<10> , 
        n128, n126, n124, n212, n122, n120, n118, n112, n110, 
        \alu_operand_a<0> }), .B({\alu_operand_b<15> , \alu_operand_b<14> , 
        n106, n209, \alu_operand_b<11> , n98, n94, n108, n82, n79, n75, n72, 
        n70, n67, n64, n61}), .Cin(Cin), .Op({\Opcode<2> , \Opcode<1> , 
        \Opcode<0> }), .invA(InvA), .invB(InvB), .sign(1'b1), .Out({
        \aluResult<15> , \aluResult<14> , \aluResult<13> , \aluResult<12> , 
        \aluResult<11> , \aluResult<10> , \aluResult<9> , \aluResult<8> , 
        \aluResult<7> , \aluResult<6> , \aluResult<5> , \aluResult<4> , 
        \aluResult<3> , \aluResult<2> , \aluResult<1> , \aluResult<0> }), 
        .Ofl(), .Z(Zero), .Cout(cout) );
  mux4to1_16_5 set_mux ( .InA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n59}), .InB({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \_2_net_<0> }), .InC({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n116}), .InD({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout}), .S({\Func<1> , \Func<0> }), .Out({\setResult<15> , 
        \setResult<14> , \setResult<13> , \setResult<12> , \setResult<11> , 
        \setResult<10> , \setResult<9> , \setResult<8> , \setResult<7> , 
        \setResult<6> , \setResult<5> , \setResult<4> , \setResult<3> , 
        \setResult<2> , \setResult<1> , \setResult<0> }) );
  cla16_1 addr_adder ( .A({\DecodeIncPC<15> , \DecodeIncPC<14> , 
        \DecodeIncPC<13> , \DecodeIncPC<12> , \DecodeIncPC<11> , 
        \DecodeIncPC<10> , \DecodeIncPC<9> , \DecodeIncPC<8> , 
        \DecodeIncPC<7> , \DecodeIncPC<6> , \DecodeIncPC<5> , \DecodeIncPC<4> , 
        \DecodeIncPC<3> , \DecodeIncPC<2> , \DecodeIncPC<1> , n23}), .B({
        \Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> , \Imm<11> , \Imm<10> , 
        \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> , \Imm<5> , \Imm<4> , \Imm<3> , 
        \Imm<2> , \Imm<1> , \Imm<0> }), .Cin(1'b0), .S({\offsetAddr<15> , 
        \offsetAddr<14> , \offsetAddr<13> , \offsetAddr<12> , \offsetAddr<11> , 
        \offsetAddr<10> , \offsetAddr<9> , \offsetAddr<8> , \offsetAddr<7> , 
        \offsetAddr<6> , \offsetAddr<5> , \offsetAddr<4> , \offsetAddr<3> , 
        \offsetAddr<2> , \offsetAddr<1> , \offsetAddr<0> }), .Cout() );
  mux4to1 branchMux ( .InA(n345), .InB(n346), .InC(\ALUOp1<15> ), .InD(n509), 
        .S({\Func<1> , \Func<0> }), .Out(branch_en) );
  INVX1 U3 ( .A(n354), .Y(n1) );
  AND2X2 U4 ( .A(n365), .B(\OpBReg<6> ), .Y(n2) );
  INVX2 U5 ( .A(n210), .Y(n371) );
  INVX2 U6 ( .A(n402), .Y(n377) );
  INVX1 U7 ( .A(\Imm<1> ), .Y(n35) );
  INVX1 U8 ( .A(\Imm<0> ), .Y(n56) );
  INVX1 U9 ( .A(\Imm<3> ), .Y(n38) );
  INVX1 U10 ( .A(Btr), .Y(n469) );
  INVX1 U11 ( .A(\DecodeIncPC<4> ), .Y(n44) );
  INVX1 U12 ( .A(\Imm<5> ), .Y(n19) );
  INVX1 U13 ( .A(\Imm<6> ), .Y(n58) );
  INVX1 U14 ( .A(\DecodeIncPC<7> ), .Y(n26) );
  INVX1 U15 ( .A(\OpBReg<14> ), .Y(n426) );
  INVX1 U16 ( .A(\OpBReg<15> ), .Y(n428) );
  INVX1 U17 ( .A(\ALUOp1<8> ), .Y(n502) );
  INVX1 U18 ( .A(\ALUOp1<9> ), .Y(n503) );
  INVX1 U19 ( .A(\OpAReg<4> ), .Y(n432) );
  INVX1 U21 ( .A(\OpAReg<13> ), .Y(n440) );
  INVX1 U22 ( .A(\OpAReg<12> ), .Y(n439) );
  INVX1 U23 ( .A(\OpBReg<2> ), .Y(n382) );
  INVX1 U24 ( .A(\OpAReg<9> ), .Y(n437) );
  INVX1 U25 ( .A(\OpAReg<14> ), .Y(n441) );
  INVX1 U26 ( .A(\OpAReg<3> ), .Y(n431) );
  INVX1 U27 ( .A(\OpAReg<7> ), .Y(n435) );
  INVX1 U28 ( .A(\OpAReg<11> ), .Y(n438) );
  INVX1 U29 ( .A(Set), .Y(n466) );
  INVX1 U30 ( .A(n443), .Y(n462) );
  OR2X1 U31 ( .A(n384), .B(n47), .Y(n443) );
  INVX1 U32 ( .A(\OpAReg<15> ), .Y(n442) );
  BUFX2 U33 ( .A(n488), .Y(n397) );
  INVX1 U34 ( .A(n355), .Y(n389) );
  INVX1 U35 ( .A(\aluResult<0> ), .Y(n492) );
  INVX1 U36 ( .A(\ForwardALUOp2<1> ), .Y(n511) );
  INVX1 U37 ( .A(\ForwardALUOp2<0> ), .Y(n510) );
  INVX1 U38 ( .A(\ForwardALUOp1<1> ), .Y(n513) );
  INVX1 U39 ( .A(\ForwardALUOp1<0> ), .Y(n512) );
  INVX1 U40 ( .A(\ALUOp1<6> ), .Y(n500) );
  INVX1 U41 ( .A(\ALUOp1<7> ), .Y(n501) );
  BUFX2 U42 ( .A(n344), .Y(n398) );
  INVX1 U43 ( .A(\ALUOp1<15> ), .Y(n509) );
  INVX1 U44 ( .A(\ALUOp1<0> ), .Y(n494) );
  INVX1 U45 ( .A(\ALUOp1<1> ), .Y(n495) );
  INVX1 U46 ( .A(\ALUOp1<10> ), .Y(n504) );
  AND2X2 U47 ( .A(n403), .B(n17), .Y(n3) );
  AND2X2 U48 ( .A(n366), .B(\OpBReg<1> ), .Y(n4) );
  AND2X2 U49 ( .A(n365), .B(\OpBReg<10> ), .Y(n5) );
  AND2X2 U50 ( .A(n358), .B(\OpBReg<0> ), .Y(n6) );
  AND2X2 U51 ( .A(n387), .B(\OpBReg<3> ), .Y(n7) );
  AND2X2 U52 ( .A(n365), .B(\OpBReg<4> ), .Y(n8) );
  AND2X2 U53 ( .A(n27), .B(\OpBReg<7> ), .Y(n9) );
  AND2X2 U54 ( .A(\aluResult<11> ), .B(n397), .Y(n332) );
  INVX1 U55 ( .A(n368), .Y(n10) );
  INVX1 U56 ( .A(Link), .Y(n11) );
  INVX1 U57 ( .A(Link), .Y(n12) );
  INVX1 U58 ( .A(n402), .Y(n13) );
  INVX1 U59 ( .A(n12), .Y(n376) );
  INVX4 U60 ( .A(n24), .Y(n358) );
  INVX1 U61 ( .A(n17), .Y(n14) );
  INVX1 U62 ( .A(\Imm<2> ), .Y(n21) );
  INVX1 U63 ( .A(n33), .Y(n15) );
  INVX1 U64 ( .A(n378), .Y(n16) );
  INVX1 U65 ( .A(\DecodeIncPC<2> ), .Y(n29) );
  INVX1 U66 ( .A(\DecodeIncPC<3> ), .Y(n40) );
  INVX1 U67 ( .A(n51), .Y(n17) );
  NOR3X1 U68 ( .A(n10), .B(n19), .C(n31), .Y(n18) );
  NOR3X1 U69 ( .A(n21), .B(n15), .C(n358), .Y(n20) );
  INVX1 U70 ( .A(\DecodeIncPC<0> ), .Y(n22) );
  INVX2 U71 ( .A(n22), .Y(n23) );
  INVX1 U72 ( .A(n369), .Y(n24) );
  AND2X2 U73 ( .A(\aluResult<13> ), .B(n397), .Y(n336) );
  NOR3X1 U74 ( .A(n364), .B(n26), .C(n14), .Y(n25) );
  INVX1 U75 ( .A(n381), .Y(n27) );
  INVX1 U76 ( .A(n13), .Y(n30) );
  NOR3X1 U77 ( .A(n29), .B(n388), .C(n30), .Y(n28) );
  INVX1 U78 ( .A(n386), .Y(n31) );
  INVX1 U79 ( .A(n31), .Y(n32) );
  INVX1 U80 ( .A(n12), .Y(n386) );
  INVX1 U81 ( .A(n367), .Y(n33) );
  NOR3X1 U82 ( .A(n27), .B(n35), .C(n375), .Y(n34) );
  INVX1 U83 ( .A(\Imm<9> ), .Y(n50) );
  INVX1 U84 ( .A(JumpReg), .Y(n36) );
  INVX1 U85 ( .A(n381), .Y(n365) );
  NOR3X1 U86 ( .A(n1), .B(n38), .C(n387), .Y(n37) );
  NOR3X1 U87 ( .A(n40), .B(n395), .C(n354), .Y(n39) );
  INVX1 U88 ( .A(n54), .Y(n41) );
  INVX2 U89 ( .A(n41), .Y(n42) );
  INVX1 U90 ( .A(JumpReg), .Y(n404) );
  NOR3X1 U91 ( .A(n387), .B(n355), .C(n44), .Y(n43) );
  INVX1 U92 ( .A(n395), .Y(n380) );
  INVX1 U93 ( .A(n386), .Y(n51) );
  AND2X2 U94 ( .A(n48), .B(n32), .Y(n45) );
  AND2X2 U95 ( .A(\DecodeIncPC<15> ), .B(n489), .Y(n46) );
  BUFX2 U96 ( .A(n146), .Y(n47) );
  INVX1 U97 ( .A(n368), .Y(n48) );
  INVX1 U98 ( .A(n367), .Y(n368) );
  NOR3X1 U99 ( .A(n385), .B(n50), .C(n51), .Y(n49) );
  INVX1 U100 ( .A(n376), .Y(n52) );
  INVX1 U101 ( .A(n30), .Y(n53) );
  OR2X2 U102 ( .A(n53), .B(n382), .Y(n409) );
  AND2X2 U103 ( .A(n368), .B(n376), .Y(n54) );
  INVX1 U104 ( .A(n381), .Y(n366) );
  INVX1 U105 ( .A(n23), .Y(n467) );
  NOR3X1 U106 ( .A(n403), .B(n56), .C(n358), .Y(n55) );
  NOR3X1 U107 ( .A(n404), .B(n58), .C(n358), .Y(n57) );
  BUFX2 U108 ( .A(Zero), .Y(n59) );
  INVX1 U109 ( .A(n54), .Y(n60) );
  OR2X2 U110 ( .A(n6), .B(n62), .Y(n61) );
  OR2X2 U111 ( .A(n55), .B(n63), .Y(n62) );
  INVX1 U112 ( .A(n407), .Y(n63) );
  OR2X2 U113 ( .A(n66), .B(n65), .Y(n64) );
  OR2X2 U114 ( .A(n34), .B(n4), .Y(n65) );
  INVX1 U115 ( .A(n408), .Y(n66) );
  OR2X2 U116 ( .A(n69), .B(n68), .Y(n67) );
  OR2X2 U117 ( .A(n20), .B(n28), .Y(n68) );
  INVX1 U118 ( .A(n409), .Y(n69) );
  OR2X2 U119 ( .A(n7), .B(n71), .Y(n70) );
  OR2X2 U129 ( .A(n37), .B(n39), .Y(n71) );
  OR2X2 U130 ( .A(n8), .B(n73), .Y(n72) );
  OR2X2 U131 ( .A(n43), .B(n74), .Y(n73) );
  INVX1 U132 ( .A(n410), .Y(n74) );
  OR2X2 U133 ( .A(n78), .B(n76), .Y(n75) );
  OR2X2 U134 ( .A(n18), .B(n77), .Y(n76) );
  INVX1 U135 ( .A(n412), .Y(n77) );
  INVX1 U136 ( .A(n411), .Y(n78) );
  OR2X2 U137 ( .A(n81), .B(n80), .Y(n79) );
  OR2X2 U138 ( .A(n57), .B(n2), .Y(n80) );
  INVX1 U139 ( .A(n413), .Y(n81) );
  OR2X2 U140 ( .A(n9), .B(n92), .Y(n82) );
  OR2X2 U141 ( .A(n93), .B(n25), .Y(n92) );
  INVX1 U142 ( .A(n414), .Y(n93) );
  OR2X2 U143 ( .A(n97), .B(n95), .Y(n94) );
  OR2X2 U144 ( .A(n49), .B(n96), .Y(n95) );
  INVX1 U145 ( .A(n417), .Y(n96) );
  INVX1 U146 ( .A(n418), .Y(n97) );
  OR2X2 U147 ( .A(n101), .B(n99), .Y(n98) );
  OR2X2 U148 ( .A(n100), .B(n5), .Y(n99) );
  INVX1 U149 ( .A(n419), .Y(n100) );
  INVX1 U150 ( .A(n420), .Y(n101) );
  OR2X2 U151 ( .A(n46), .B(n103), .Y(\Result<15> ) );
  OR2X2 U152 ( .A(n340), .B(n104), .Y(n103) );
  INVX1 U153 ( .A(n487), .Y(n104) );
  AND2X2 U154 ( .A(n362), .B(n424), .Y(n105) );
  INVX1 U155 ( .A(n105), .Y(n106) );
  AND2X2 U156 ( .A(n374), .B(n415), .Y(n107) );
  INVX1 U157 ( .A(n107), .Y(n108) );
  AND2X2 U159 ( .A(n390), .B(n429), .Y(n109) );
  INVX1 U160 ( .A(n109), .Y(n110) );
  AND2X2 U161 ( .A(n430), .B(n396), .Y(n111) );
  INVX1 U162 ( .A(n111), .Y(n112) );
  AND2X2 U163 ( .A(n405), .B(n406), .Y(n115) );
  INVX1 U164 ( .A(n115), .Y(n116) );
  OR2X2 U165 ( .A(n393), .B(n431), .Y(n117) );
  INVX1 U166 ( .A(n117), .Y(n118) );
  OR2X2 U167 ( .A(n391), .B(n432), .Y(n119) );
  INVX1 U168 ( .A(n119), .Y(n120) );
  OR2X2 U169 ( .A(n391), .B(n433), .Y(n121) );
  INVX1 U170 ( .A(n121), .Y(n122) );
  OR2X2 U171 ( .A(n393), .B(n435), .Y(n123) );
  INVX1 U172 ( .A(n123), .Y(n124) );
  OR2X2 U173 ( .A(n391), .B(n436), .Y(n125) );
  INVX1 U174 ( .A(n125), .Y(n126) );
  OR2X2 U175 ( .A(n393), .B(n437), .Y(n127) );
  INVX1 U176 ( .A(n127), .Y(n128) );
  OR2X2 U177 ( .A(n372), .B(n439), .Y(n129) );
  INVX1 U178 ( .A(n129), .Y(n130) );
  OR2X2 U179 ( .A(n372), .B(n440), .Y(n131) );
  INVX1 U180 ( .A(n131), .Y(n132) );
  OR2X2 U181 ( .A(n371), .B(n441), .Y(n133) );
  INVX1 U182 ( .A(n133), .Y(n134) );
  AND2X2 U183 ( .A(n452), .B(n224), .Y(n135) );
  INVX1 U184 ( .A(n135), .Y(\NextPC<6> ) );
  AND2X2 U185 ( .A(n453), .B(n226), .Y(n137) );
  INVX1 U186 ( .A(n137), .Y(\NextPC<7> ) );
  AND2X2 U187 ( .A(n454), .B(n228), .Y(n139) );
  INVX1 U188 ( .A(n139), .Y(\NextPC<8> ) );
  AND2X2 U189 ( .A(n455), .B(n230), .Y(n141) );
  INVX1 U190 ( .A(n141), .Y(\NextPC<9> ) );
  AND2X2 U191 ( .A(n456), .B(n232), .Y(n143) );
  INVX1 U192 ( .A(n143), .Y(\NextPC<10> ) );
  AND2X2 U193 ( .A(n457), .B(n458), .Y(n145) );
  INVX1 U194 ( .A(n145), .Y(\NextPC<11> ) );
  AND2X2 U195 ( .A(n459), .B(n234), .Y(n152) );
  INVX1 U196 ( .A(n152), .Y(\NextPC<12> ) );
  AND2X2 U197 ( .A(n460), .B(n236), .Y(n184) );
  INVX1 U198 ( .A(n184), .Y(\NextPC<13> ) );
  AND2X2 U199 ( .A(n461), .B(n238), .Y(n187) );
  INVX1 U200 ( .A(n187), .Y(\NextPC<14> ) );
  AND2X2 U201 ( .A(n464), .B(n465), .Y(n204) );
  INVX1 U202 ( .A(n204), .Y(\NextPC<15> ) );
  AND2X2 U203 ( .A(n113), .B(n114), .Y(n206) );
  INVX1 U204 ( .A(n206), .Y(\Result<1> ) );
  AND2X2 U205 ( .A(n360), .B(n423), .Y(n208) );
  INVX1 U206 ( .A(n208), .Y(n209) );
  OR2X2 U207 ( .A(n33), .B(n52), .Y(n210) );
  OR2X2 U208 ( .A(n391), .B(n434), .Y(n211) );
  INVX1 U209 ( .A(n211), .Y(n212) );
  OR2X2 U210 ( .A(n371), .B(n442), .Y(n213) );
  INVX1 U211 ( .A(n213), .Y(n214) );
  AND2X2 U212 ( .A(n448), .B(n220), .Y(n215) );
  INVX1 U213 ( .A(n215), .Y(\NextPC<3> ) );
  AND2X2 U214 ( .A(n451), .B(n222), .Y(n217) );
  INVX1 U215 ( .A(n217), .Y(\NextPC<5> ) );
  AND2X1 U218 ( .A(\aluResult<3> ), .B(n384), .Y(n219) );
  INVX1 U219 ( .A(n219), .Y(n220) );
  AND2X1 U222 ( .A(\aluResult<5> ), .B(n384), .Y(n221) );
  INVX1 U225 ( .A(n221), .Y(n222) );
  AND2X1 U228 ( .A(\aluResult<6> ), .B(n384), .Y(n223) );
  INVX1 U231 ( .A(n223), .Y(n224) );
  AND2X1 U234 ( .A(\aluResult<7> ), .B(n384), .Y(n225) );
  INVX1 U237 ( .A(n225), .Y(n226) );
  AND2X1 U240 ( .A(\aluResult<8> ), .B(n384), .Y(n227) );
  INVX1 U243 ( .A(n227), .Y(n228) );
  AND2X1 U246 ( .A(\aluResult<9> ), .B(n384), .Y(n229) );
  INVX1 U249 ( .A(n229), .Y(n230) );
  AND2X1 U252 ( .A(\aluResult<10> ), .B(n384), .Y(n231) );
  INVX1 U255 ( .A(n231), .Y(n232) );
  AND2X1 U258 ( .A(\aluResult<12> ), .B(n384), .Y(n233) );
  INVX1 U261 ( .A(n233), .Y(n234) );
  AND2X1 U264 ( .A(\aluResult<13> ), .B(n384), .Y(n235) );
  INVX1 U266 ( .A(n235), .Y(n236) );
  AND2X1 U267 ( .A(\aluResult<14> ), .B(n384), .Y(n237) );
  INVX1 U270 ( .A(n237), .Y(n238) );
  AND2X2 U301 ( .A(\DecodeIncPC<2> ), .B(n489), .Y(n239) );
  INVX1 U302 ( .A(n239), .Y(n240) );
  AND2X2 U303 ( .A(\DecodeIncPC<3> ), .B(n489), .Y(n241) );
  INVX1 U304 ( .A(n241), .Y(n242) );
  AND2X2 U307 ( .A(\DecodeIncPC<4> ), .B(n489), .Y(n243) );
  INVX1 U308 ( .A(n243), .Y(n244) );
  AND2X2 U309 ( .A(\DecodeIncPC<5> ), .B(n489), .Y(n245) );
  INVX1 U310 ( .A(n245), .Y(n246) );
  AND2X2 U311 ( .A(\DecodeIncPC<6> ), .B(n489), .Y(n247) );
  INVX1 U312 ( .A(n247), .Y(n248) );
  AND2X2 U313 ( .A(\DecodeIncPC<7> ), .B(n489), .Y(n249) );
  INVX1 U314 ( .A(n249), .Y(n250) );
  AND2X2 U315 ( .A(\DecodeIncPC<8> ), .B(n489), .Y(n251) );
  INVX1 U316 ( .A(n251), .Y(n252) );
  AND2X2 U317 ( .A(\DecodeIncPC<9> ), .B(n489), .Y(n253) );
  INVX1 U318 ( .A(n253), .Y(n254) );
  AND2X2 U319 ( .A(\DecodeIncPC<10> ), .B(n489), .Y(n255) );
  INVX1 U320 ( .A(n255), .Y(n256) );
  AND2X2 U321 ( .A(\DecodeIncPC<11> ), .B(n489), .Y(n257) );
  INVX1 U322 ( .A(n257), .Y(n258) );
  AND2X2 U323 ( .A(\DecodeIncPC<12> ), .B(n489), .Y(n259) );
  INVX1 U324 ( .A(n259), .Y(n260) );
  AND2X2 U325 ( .A(\DecodeIncPC<13> ), .B(n489), .Y(n261) );
  INVX1 U326 ( .A(n261), .Y(n262) );
  AND2X2 U327 ( .A(\DecodeIncPC<14> ), .B(n489), .Y(n263) );
  INVX1 U328 ( .A(n263), .Y(n264) );
  BUFX2 U329 ( .A(\aluResult<15> ), .Y(n265) );
  AND2X2 U330 ( .A(n449), .B(n450), .Y(n266) );
  INVX1 U331 ( .A(n266), .Y(\NextPC<4> ) );
  AND2X2 U332 ( .A(n182), .B(n183), .Y(n268) );
  INVX1 U333 ( .A(n268), .Y(n269) );
  AND2X2 U334 ( .A(n180), .B(n181), .Y(n270) );
  INVX1 U335 ( .A(n270), .Y(n271) );
  AND2X2 U336 ( .A(n178), .B(n179), .Y(n272) );
  INVX1 U337 ( .A(n272), .Y(n273) );
  AND2X2 U338 ( .A(n176), .B(n177), .Y(n274) );
  INVX1 U339 ( .A(n274), .Y(n275) );
  AND2X2 U340 ( .A(n174), .B(n175), .Y(n276) );
  INVX1 U341 ( .A(n276), .Y(n277) );
  AND2X2 U342 ( .A(n172), .B(n173), .Y(n278) );
  INVX1 U343 ( .A(n278), .Y(n279) );
  AND2X2 U344 ( .A(n170), .B(n171), .Y(n280) );
  INVX1 U345 ( .A(n280), .Y(n281) );
  AND2X2 U346 ( .A(n168), .B(n169), .Y(n282) );
  INVX1 U347 ( .A(n282), .Y(n283) );
  AND2X2 U348 ( .A(n166), .B(n167), .Y(n284) );
  INVX1 U349 ( .A(n284), .Y(n285) );
  AND2X2 U350 ( .A(n164), .B(n165), .Y(n286) );
  INVX1 U351 ( .A(n286), .Y(n287) );
  AND2X2 U352 ( .A(n162), .B(n163), .Y(n288) );
  INVX1 U353 ( .A(n288), .Y(n289) );
  AND2X2 U354 ( .A(n160), .B(n161), .Y(n290) );
  INVX1 U355 ( .A(n290), .Y(n291) );
  AND2X2 U356 ( .A(n158), .B(n159), .Y(n292) );
  INVX1 U357 ( .A(n292), .Y(n293) );
  AND2X2 U358 ( .A(n156), .B(n157), .Y(n294) );
  INVX1 U359 ( .A(n294), .Y(n295) );
  AND2X2 U360 ( .A(n154), .B(n155), .Y(n296) );
  INVX1 U361 ( .A(n296), .Y(n297) );
  AND2X2 U362 ( .A(n147), .B(n148), .Y(n298) );
  INVX1 U363 ( .A(n298), .Y(n299) );
  OR2X1 U364 ( .A(n349), .B(n301), .Y(n300) );
  OR2X1 U365 ( .A(n348), .B(n343), .Y(n301) );
  OR2X1 U366 ( .A(n351), .B(n303), .Y(n302) );
  OR2X1 U367 ( .A(n350), .B(n352), .Y(n303) );
  AND2X2 U368 ( .A(n446), .B(n447), .Y(n304) );
  INVX1 U369 ( .A(n304), .Y(\NextPC<2> ) );
  AND2X1 U370 ( .A(\aluResult<0> ), .B(n397), .Y(n306) );
  INVX1 U371 ( .A(n306), .Y(n307) );
  BUFX2 U372 ( .A(n149), .Y(n400) );
  AND2X1 U373 ( .A(ALUSrc), .B(n352), .Y(n150) );
  BUFX2 U374 ( .A(n519), .Y(\Result<3> ) );
  BUFX2 U375 ( .A(n518), .Y(\Result<4> ) );
  BUFX2 U376 ( .A(n517), .Y(\Result<7> ) );
  BUFX2 U377 ( .A(n516), .Y(\Result<8> ) );
  BUFX2 U378 ( .A(n515), .Y(\Result<9> ) );
  BUFX2 U379 ( .A(n514), .Y(\Result<11> ) );
  AND2X1 U380 ( .A(\aluResult<2> ), .B(n397), .Y(n314) );
  INVX1 U381 ( .A(n314), .Y(n315) );
  AND2X1 U382 ( .A(\aluResult<3> ), .B(n397), .Y(n316) );
  INVX1 U383 ( .A(n316), .Y(n317) );
  AND2X1 U384 ( .A(\aluResult<4> ), .B(n397), .Y(n318) );
  INVX1 U385 ( .A(n318), .Y(n319) );
  AND2X1 U386 ( .A(\aluResult<5> ), .B(n397), .Y(n320) );
  INVX1 U387 ( .A(n320), .Y(n321) );
  AND2X1 U388 ( .A(\aluResult<6> ), .B(n397), .Y(n322) );
  INVX1 U389 ( .A(n322), .Y(n323) );
  AND2X1 U390 ( .A(\aluResult<7> ), .B(n397), .Y(n324) );
  INVX1 U391 ( .A(n324), .Y(n325) );
  AND2X1 U392 ( .A(\aluResult<8> ), .B(n397), .Y(n326) );
  INVX1 U393 ( .A(n326), .Y(n327) );
  AND2X1 U394 ( .A(\aluResult<9> ), .B(n397), .Y(n328) );
  INVX1 U395 ( .A(n328), .Y(n329) );
  AND2X1 U396 ( .A(\aluResult<10> ), .B(n397), .Y(n330) );
  INVX1 U397 ( .A(n330), .Y(n331) );
  INVX1 U398 ( .A(n332), .Y(n333) );
  AND2X1 U399 ( .A(\aluResult<12> ), .B(n397), .Y(n334) );
  INVX1 U400 ( .A(n334), .Y(n335) );
  INVX1 U401 ( .A(n336), .Y(n337) );
  AND2X1 U402 ( .A(\aluResult<14> ), .B(n397), .Y(n338) );
  INVX1 U403 ( .A(n338), .Y(n339) );
  AND2X2 U404 ( .A(n265), .B(n397), .Y(n340) );
  INVX1 U405 ( .A(\ALUOp1<12> ), .Y(n506) );
  INVX1 U406 ( .A(\ALUOp1<11> ), .Y(n505) );
  INVX1 U407 ( .A(\ALUOp1<14> ), .Y(n508) );
  INVX1 U408 ( .A(\ALUOp1<13> ), .Y(n507) );
  INVX1 U409 ( .A(\ALUOp1<5> ), .Y(n499) );
  INVX1 U410 ( .A(\ALUOp1<4> ), .Y(n498) );
  INVX1 U411 ( .A(\ALUOp1<3> ), .Y(n497) );
  INVX1 U412 ( .A(\ALUOp1<2> ), .Y(n496) );
  OR2X2 U413 ( .A(n45), .B(n438), .Y(n341) );
  INVX1 U414 ( .A(n341), .Y(n342) );
  AND2X1 U415 ( .A(n512), .B(n513), .Y(n343) );
  INVX1 U416 ( .A(n343), .Y(n344) );
  INVX1 U417 ( .A(\aluResult<1> ), .Y(n493) );
  INVX1 U418 ( .A(n347), .Y(n345) );
  INVX1 U419 ( .A(n345), .Y(n346) );
  BUFX2 U420 ( .A(_7_net_), .Y(n347) );
  AND2X1 U421 ( .A(\ForwardALUOp1<1> ), .B(n512), .Y(n348) );
  AND2X1 U422 ( .A(\ForwardALUOp1<0> ), .B(n513), .Y(n349) );
  AND2X1 U423 ( .A(\ForwardALUOp2<1> ), .B(n510), .Y(n350) );
  AND2X1 U424 ( .A(\ForwardALUOp2<0> ), .B(n511), .Y(n351) );
  INVX1 U425 ( .A(n472), .Y(n489) );
  INVX1 U426 ( .A(n473), .Y(n490) );
  AND2X1 U427 ( .A(n510), .B(n511), .Y(n352) );
  INVX1 U428 ( .A(n352), .Y(n353) );
  INVX1 U429 ( .A(BranchJumpTaken), .Y(n463) );
  BUFX2 U430 ( .A(n344), .Y(n399) );
  OAI21X1 U431 ( .A(n470), .B(n473), .C(n471), .Y(\Result<0> ) );
  INVX1 U432 ( .A(n385), .Y(n354) );
  INVX1 U433 ( .A(n404), .Y(n355) );
  INVX1 U434 ( .A(n36), .Y(n388) );
  INVX1 U435 ( .A(n11), .Y(n356) );
  INVX1 U436 ( .A(n370), .Y(n357) );
  NAND2X1 U437 ( .A(n403), .B(n377), .Y(n359) );
  NAND2X1 U438 ( .A(\OpBReg<12> ), .B(n378), .Y(n360) );
  INVX1 U439 ( .A(n354), .Y(n361) );
  OR2X2 U440 ( .A(n60), .B(n416), .Y(n374) );
  NAND2X1 U441 ( .A(\OpBReg<13> ), .B(n14), .Y(n362) );
  INVX1 U442 ( .A(n54), .Y(n363) );
  INVX1 U443 ( .A(n404), .Y(n364) );
  INVX1 U444 ( .A(n401), .Y(n387) );
  INVX1 U445 ( .A(JumpReg), .Y(n367) );
  INVX1 U446 ( .A(Link), .Y(n369) );
  INVX1 U447 ( .A(n369), .Y(n370) );
  INVX1 U448 ( .A(n210), .Y(n372) );
  INVX1 U449 ( .A(n10), .Y(n373) );
  INVX1 U450 ( .A(\Imm<8> ), .Y(n416) );
  INVX1 U451 ( .A(n355), .Y(n375) );
  AND2X2 U452 ( .A(n392), .B(\OpAReg<0> ), .Y(\alu_operand_a<0> ) );
  INVX1 U453 ( .A(n357), .Y(n401) );
  INVX1 U454 ( .A(n401), .Y(n378) );
  INVX1 U455 ( .A(n378), .Y(n379) );
  INVX1 U456 ( .A(n12), .Y(n381) );
  INVX1 U457 ( .A(JumpReg), .Y(n403) );
  INVX1 U458 ( .A(n384), .Y(n383) );
  INVX1 U459 ( .A(n389), .Y(n384) );
  INVX1 U460 ( .A(Link), .Y(n402) );
  INVX1 U461 ( .A(JumpReg), .Y(n385) );
  NAND2X1 U462 ( .A(n52), .B(\OpAReg<1> ), .Y(n390) );
  AND2X2 U463 ( .A(n36), .B(n13), .Y(n391) );
  INVX1 U464 ( .A(n45), .Y(n392) );
  AND2X2 U465 ( .A(n370), .B(n385), .Y(n393) );
  MUX2X1 U466 ( .B(\ALUOp1<15> ), .A(n265), .S(n394), .Y(n405) );
  XNOR2X1 U467 ( .A(\ALUOp1<15> ), .B(\ALUOp2<15> ), .Y(n394) );
  AND2X2 U468 ( .A(\OpAReg<10> ), .B(n359), .Y(\alu_operand_a<10> ) );
  NAND2X1 U469 ( .A(n395), .B(\OpAReg<2> ), .Y(n396) );
  INVX1 U470 ( .A(n370), .Y(n395) );
  INVX1 U471 ( .A(n405), .Y(\_2_net_<0> ) );
  INVX1 U472 ( .A(Zero), .Y(n406) );
  INVX1 U473 ( .A(\setResult<0> ), .Y(n470) );
  NAND3X1 U474 ( .A(n403), .B(\DecodeIncPC<0> ), .C(n356), .Y(n407) );
  NAND3X1 U475 ( .A(n48), .B(\DecodeIncPC<1> ), .C(n13), .Y(n408) );
  NAND3X1 U476 ( .A(n373), .B(\Imm<4> ), .C(n379), .Y(n410) );
  NAND2X1 U477 ( .A(n358), .B(\OpBReg<5> ), .Y(n412) );
  NAND3X1 U478 ( .A(n48), .B(\DecodeIncPC<5> ), .C(n376), .Y(n411) );
  NAND3X1 U479 ( .A(n361), .B(\DecodeIncPC<6> ), .C(n377), .Y(n413) );
  NAND3X1 U480 ( .A(n373), .B(\Imm<7> ), .C(n16), .Y(n414) );
  AOI22X1 U481 ( .A(\DecodeIncPC<8> ), .B(n393), .C(n14), .D(\OpBReg<8> ), .Y(
        n415) );
  NAND3X1 U482 ( .A(n361), .B(\DecodeIncPC<9> ), .C(n377), .Y(n418) );
  NAND2X1 U483 ( .A(\OpBReg<9> ), .B(n357), .Y(n417) );
  NAND3X1 U484 ( .A(n364), .B(\Imm<10> ), .C(n32), .Y(n420) );
  NAND3X1 U485 ( .A(n377), .B(n389), .C(\DecodeIncPC<10> ), .Y(n419) );
  INVX2 U486 ( .A(\Imm<11> ), .Y(n422) );
  AOI22X1 U487 ( .A(\DecodeIncPC<11> ), .B(n3), .C(n366), .D(\OpBReg<11> ), 
        .Y(n421) );
  OAI21X1 U488 ( .A(n363), .B(n422), .C(n421), .Y(\alu_operand_b<11> ) );
  AOI22X1 U489 ( .A(\DecodeIncPC<12> ), .B(n372), .C(\Imm<12> ), .D(n42), .Y(
        n423) );
  AOI22X1 U490 ( .A(\DecodeIncPC<13> ), .B(n371), .C(\Imm<13> ), .D(n42), .Y(
        n424) );
  AOI22X1 U491 ( .A(\DecodeIncPC<14> ), .B(n3), .C(\Imm<14> ), .D(n42), .Y(
        n425) );
  OAI21X1 U492 ( .A(n426), .B(n380), .C(n425), .Y(\alu_operand_b<14> ) );
  AOI22X1 U493 ( .A(\DecodeIncPC<15> ), .B(n371), .C(\Imm<15> ), .D(n42), .Y(
        n427) );
  OAI21X1 U494 ( .A(n428), .B(n380), .C(n427), .Y(\alu_operand_b<15> ) );
  NAND2X1 U495 ( .A(\OpAReg<1> ), .B(n364), .Y(n429) );
  NAND2X1 U496 ( .A(\OpAReg<2> ), .B(n33), .Y(n430) );
  INVX2 U497 ( .A(\OpAReg<5> ), .Y(n433) );
  INVX2 U498 ( .A(\OpAReg<6> ), .Y(n434) );
  INVX2 U499 ( .A(\OpAReg<8> ), .Y(n436) );
  NAND2X1 U500 ( .A(n146), .B(n383), .Y(BranchJumpTaken) );
  AOI22X1 U501 ( .A(\IncPC<0> ), .B(n463), .C(\offsetAddr<0> ), .D(n462), .Y(
        n444) );
  OAI21X1 U502 ( .A(n389), .B(n492), .C(n444), .Y(\NextPC<0> ) );
  AOI22X1 U503 ( .A(\IncPC<1> ), .B(n463), .C(\offsetAddr<1> ), .D(n462), .Y(
        n445) );
  OAI21X1 U504 ( .A(n389), .B(n493), .C(n445), .Y(\NextPC<1> ) );
  NAND2X1 U505 ( .A(\aluResult<2> ), .B(n384), .Y(n447) );
  AOI22X1 U506 ( .A(\IncPC<2> ), .B(n463), .C(\offsetAddr<2> ), .D(n462), .Y(
        n446) );
  AOI22X1 U507 ( .A(\IncPC<3> ), .B(n463), .C(\offsetAddr<3> ), .D(n462), .Y(
        n448) );
  NAND2X1 U508 ( .A(\aluResult<4> ), .B(n384), .Y(n450) );
  AOI22X1 U509 ( .A(\IncPC<4> ), .B(n463), .C(\offsetAddr<4> ), .D(n462), .Y(
        n449) );
  AOI22X1 U510 ( .A(\IncPC<5> ), .B(n463), .C(\offsetAddr<5> ), .D(n462), .Y(
        n451) );
  AOI22X1 U511 ( .A(\IncPC<6> ), .B(n463), .C(\offsetAddr<6> ), .D(n462), .Y(
        n452) );
  AOI22X1 U512 ( .A(\IncPC<7> ), .B(n463), .C(\offsetAddr<7> ), .D(n462), .Y(
        n453) );
  AOI22X1 U513 ( .A(\IncPC<8> ), .B(n463), .C(\offsetAddr<8> ), .D(n462), .Y(
        n454) );
  AOI22X1 U514 ( .A(\IncPC<9> ), .B(n463), .C(\offsetAddr<9> ), .D(n462), .Y(
        n455) );
  AOI22X1 U515 ( .A(\IncPC<10> ), .B(n463), .C(\offsetAddr<10> ), .D(n462), 
        .Y(n456) );
  NAND2X1 U516 ( .A(n384), .B(\aluResult<11> ), .Y(n458) );
  AOI22X1 U517 ( .A(\IncPC<11> ), .B(n463), .C(\offsetAddr<11> ), .D(n462), 
        .Y(n457) );
  AOI22X1 U518 ( .A(\IncPC<12> ), .B(n463), .C(\offsetAddr<12> ), .D(n462), 
        .Y(n459) );
  AOI22X1 U519 ( .A(\IncPC<13> ), .B(n463), .C(\offsetAddr<13> ), .D(n462), 
        .Y(n460) );
  AOI22X1 U520 ( .A(\IncPC<14> ), .B(n463), .C(\offsetAddr<14> ), .D(n462), 
        .Y(n461) );
  NAND2X1 U521 ( .A(n384), .B(n265), .Y(n465) );
  AOI22X1 U522 ( .A(\IncPC<15> ), .B(n463), .C(\offsetAddr<15> ), .D(n462), 
        .Y(n464) );
  NAND3X1 U523 ( .A(n466), .B(n384), .C(n469), .Y(n472) );
  NOR3X1 U524 ( .A(Btr), .B(n384), .C(Set), .Y(n488) );
  OAI21X1 U525 ( .A(n472), .B(n467), .C(n307), .Y(n468) );
  AOI21X1 U526 ( .A(\ALUOp1<15> ), .B(Btr), .C(n468), .Y(n471) );
  NAND2X1 U527 ( .A(n469), .B(Set), .Y(n473) );
  AOI22X1 U528 ( .A(\ALUOp1<13> ), .B(Btr), .C(\setResult<2> ), .D(n490), .Y(
        n474) );
  NAND3X1 U529 ( .A(n240), .B(n474), .C(n315), .Y(\Result<2> ) );
  AOI22X1 U530 ( .A(\ALUOp1<12> ), .B(Btr), .C(\setResult<3> ), .D(n490), .Y(
        n475) );
  NAND3X1 U531 ( .A(n242), .B(n475), .C(n317), .Y(n519) );
  AOI22X1 U532 ( .A(\ALUOp1<11> ), .B(Btr), .C(\setResult<4> ), .D(n490), .Y(
        n476) );
  NAND3X1 U533 ( .A(n244), .B(n476), .C(n319), .Y(n518) );
  AOI22X1 U534 ( .A(\ALUOp1<10> ), .B(Btr), .C(\setResult<5> ), .D(n490), .Y(
        n477) );
  NAND3X1 U535 ( .A(n246), .B(n477), .C(n321), .Y(\Result<5> ) );
  AOI22X1 U536 ( .A(\ALUOp1<9> ), .B(Btr), .C(\setResult<6> ), .D(n490), .Y(
        n478) );
  NAND3X1 U537 ( .A(n248), .B(n478), .C(n323), .Y(\Result<6> ) );
  AOI22X1 U538 ( .A(\ALUOp1<8> ), .B(Btr), .C(\setResult<7> ), .D(n490), .Y(
        n479) );
  NAND3X1 U539 ( .A(n250), .B(n479), .C(n325), .Y(n517) );
  AOI22X1 U540 ( .A(\ALUOp1<7> ), .B(Btr), .C(\setResult<8> ), .D(n490), .Y(
        n480) );
  NAND3X1 U541 ( .A(n252), .B(n480), .C(n327), .Y(n516) );
  AOI22X1 U542 ( .A(\ALUOp1<6> ), .B(Btr), .C(\setResult<9> ), .D(n490), .Y(
        n481) );
  NAND3X1 U543 ( .A(n254), .B(n481), .C(n329), .Y(n515) );
  AOI22X1 U544 ( .A(\ALUOp1<5> ), .B(Btr), .C(\setResult<10> ), .D(n490), .Y(
        n482) );
  NAND3X1 U545 ( .A(n256), .B(n482), .C(n331), .Y(\Result<10> ) );
  AOI22X1 U546 ( .A(\ALUOp1<4> ), .B(Btr), .C(\setResult<11> ), .D(n490), .Y(
        n483) );
  NAND3X1 U547 ( .A(n258), .B(n483), .C(n333), .Y(n514) );
  AOI22X1 U548 ( .A(\ALUOp1<3> ), .B(Btr), .C(\setResult<12> ), .D(n490), .Y(
        n484) );
  NAND3X1 U549 ( .A(n260), .B(n484), .C(n335), .Y(\Result<12> ) );
  AOI22X1 U550 ( .A(\ALUOp1<2> ), .B(Btr), .C(\setResult<13> ), .D(n490), .Y(
        n485) );
  NAND3X1 U551 ( .A(n262), .B(n485), .C(n337), .Y(\Result<13> ) );
  AOI22X1 U552 ( .A(\ALUOp1<1> ), .B(Btr), .C(\setResult<14> ), .D(n490), .Y(
        n486) );
  NAND3X1 U553 ( .A(n264), .B(n486), .C(n339), .Y(\Result<14> ) );
  AOI22X1 U554 ( .A(\ALUOp1<0> ), .B(Btr), .C(\setResult<15> ), .D(n490), .Y(
        n487) );
  AOI22X1 U555 ( .A(\DecodeIncPC<1> ), .B(n489), .C(\aluResult<1> ), .D(n397), 
        .Y(n114) );
endmodule


module pipe_em ( Stall, rst, clk, .Result({\Result<15> , \Result<14> , 
        \Result<13> , \Result<12> , \Result<11> , \Result<10> , \Result<9> , 
        \Result<8> , \Result<7> , \Result<6> , \Result<5> , \Result<4> , 
        \Result<3> , \Result<2> , \Result<1> , \Result<0> }), MemRead, 
        MemWrite, MemToReg, Halt, .ALUOp2({\ALUOp2<15> , \ALUOp2<14> , 
        \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , 
        \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , 
        \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), RegFileWrEn, 
    .Rs({\Rs<2> , \Rs<1> , \Rs<0> }), .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({
        \Rd<2> , \Rd<1> , \Rd<0> }), .WriteReg({\WriteReg<2> , \WriteReg<1> , 
        \WriteReg<0> }), .Address({\Address<15> , \Address<14> , \Address<13> , 
        \Address<12> , \Address<11> , \Address<10> , \Address<9> , 
        \Address<8> , \Address<7> , \Address<6> , \Address<5> , \Address<4> , 
        \Address<3> , \Address<2> , \Address<1> , \Address<0> }), MemRead_Out, 
        MemWrite_Out, MemToReg_Out, Halt_Out, .WriteData({\WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), RegFileWrEn_Out, 
    .Rs_Out({\Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> }), .Rt_Out({\Rt_Out<2> , 
        \Rt_Out<1> , \Rt_Out<0> }), .Rd_Out({\Rd_Out<2> , \Rd_Out<1> , 
        \Rd_Out<0> }), .WriteReg_Out({\WriteReg_Out<2> , \WriteReg_Out<1> , 
        \WriteReg_Out<0> }) );
  input Stall, rst, clk, \Result<15> , \Result<14> , \Result<13> ,
         \Result<12> , \Result<11> , \Result<10> , \Result<9> , \Result<8> ,
         \Result<7> , \Result<6> , \Result<5> , \Result<4> , \Result<3> ,
         \Result<2> , \Result<1> , \Result<0> , MemRead, MemWrite, MemToReg,
         Halt, \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , RegFileWrEn, \Rs<2> , \Rs<1> , \Rs<0> ,
         \Rt<2> , \Rt<1> , \Rt<0> , \Rd<2> , \Rd<1> , \Rd<0> , \WriteReg<2> ,
         \WriteReg<1> , \WriteReg<0> ;
  output \Address<15> , \Address<14> , \Address<13> , \Address<12> ,
         \Address<11> , \Address<10> , \Address<9> , \Address<8> ,
         \Address<7> , \Address<6> , \Address<5> , \Address<4> , \Address<3> ,
         \Address<2> , \Address<1> , \Address<0> , MemRead_Out, MemWrite_Out,
         MemToReg_Out, Halt_Out, \WriteData<15> , \WriteData<14> ,
         \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> ,
         \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> ,
         \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> ,
         \WriteData<1> , \WriteData<0> , RegFileWrEn_Out, \Rs_Out<2> ,
         \Rs_Out<1> , \Rs_Out<0> , \Rt_Out<2> , \Rt_Out<1> , \Rt_Out<0> ,
         \Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> , \WriteReg_Out<2> ,
         \WriteReg_Out<1> , \WriteReg_Out<0> ;
  wire   n125, n126, n127, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n77, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n2, n4, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n69, n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82,
         n83, n84, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124;

  AOI22X1 U51 ( .A(\WriteReg<2> ), .B(n10), .C(\WriteReg_Out<2> ), .D(n9), .Y(
        n52) );
  AOI22X1 U52 ( .A(\WriteReg<1> ), .B(n10), .C(\WriteReg_Out<1> ), .D(n9), .Y(
        n53) );
  AOI22X1 U53 ( .A(\WriteReg<0> ), .B(n10), .C(\WriteReg_Out<0> ), .D(n9), .Y(
        n54) );
  AOI22X1 U54 ( .A(\Rt<2> ), .B(n10), .C(\Rt_Out<2> ), .D(n9), .Y(n55) );
  AOI22X1 U55 ( .A(\Rt<1> ), .B(n10), .C(\Rt_Out<1> ), .D(n9), .Y(n56) );
  AOI22X1 U56 ( .A(\Rt<0> ), .B(n10), .C(\Rt_Out<0> ), .D(n9), .Y(n57) );
  AOI22X1 U57 ( .A(\Rs<2> ), .B(n10), .C(\Rs_Out<2> ), .D(n9), .Y(n58) );
  AOI22X1 U58 ( .A(\Rs<1> ), .B(n10), .C(\Rs_Out<1> ), .D(n9), .Y(n59) );
  AOI22X1 U59 ( .A(\Rs<0> ), .B(n10), .C(\Rs_Out<0> ), .D(n9), .Y(n60) );
  AOI22X1 U60 ( .A(RegFileWrEn), .B(n10), .C(RegFileWrEn_Out), .D(n9), .Y(n61)
         );
  AOI22X1 U61 ( .A(\Rd<2> ), .B(n10), .C(\Rd_Out<2> ), .D(n9), .Y(n62) );
  AOI22X1 U62 ( .A(\Rd<1> ), .B(n10), .C(\Rd_Out<1> ), .D(n9), .Y(n63) );
  AOI22X1 U63 ( .A(\Rd<0> ), .B(n10), .C(\Rd_Out<0> ), .D(n9), .Y(n64) );
  AOI22X1 U64 ( .A(MemWrite), .B(n10), .C(MemWrite_Out), .D(n9), .Y(n65) );
  AOI22X1 U65 ( .A(MemToReg), .B(n10), .C(MemToReg_Out), .D(n9), .Y(n66) );
  AOI22X1 U66 ( .A(MemRead), .B(n10), .C(MemRead_Out), .D(n9), .Y(n67) );
  AOI22X1 U67 ( .A(Halt), .B(n10), .C(Halt_Out), .D(n9), .Y(n68) );
  AOI22X1 U76 ( .A(\Address<1> ), .B(n7), .C(\Result<1> ), .D(n10), .Y(n77) );
  AOI22X1 U84 ( .A(\ALUOp2<9> ), .B(n10), .C(\WriteData<9> ), .D(n8), .Y(n85)
         );
  AOI22X1 U85 ( .A(\ALUOp2<8> ), .B(n10), .C(\WriteData<8> ), .D(n8), .Y(n86)
         );
  AOI22X1 U86 ( .A(\ALUOp2<7> ), .B(n10), .C(\WriteData<7> ), .D(n8), .Y(n87)
         );
  AOI22X1 U87 ( .A(\ALUOp2<6> ), .B(n10), .C(\WriteData<6> ), .D(n8), .Y(n88)
         );
  AOI22X1 U88 ( .A(\ALUOp2<5> ), .B(n10), .C(\WriteData<5> ), .D(n8), .Y(n89)
         );
  AOI22X1 U89 ( .A(\ALUOp2<4> ), .B(n10), .C(\WriteData<4> ), .D(n8), .Y(n90)
         );
  AOI22X1 U90 ( .A(\ALUOp2<3> ), .B(n10), .C(\WriteData<3> ), .D(n8), .Y(n91)
         );
  AOI22X1 U91 ( .A(\ALUOp2<2> ), .B(n10), .C(\WriteData<2> ), .D(n8), .Y(n92)
         );
  AOI22X1 U92 ( .A(\ALUOp2<1> ), .B(n10), .C(\WriteData<1> ), .D(n8), .Y(n93)
         );
  AOI22X1 U93 ( .A(\ALUOp2<15> ), .B(n10), .C(\WriteData<15> ), .D(n8), .Y(n94) );
  AOI22X1 U94 ( .A(\ALUOp2<14> ), .B(n10), .C(\WriteData<14> ), .D(n8), .Y(n95) );
  AOI22X1 U95 ( .A(\ALUOp2<13> ), .B(n10), .C(\WriteData<13> ), .D(n8), .Y(n96) );
  AOI22X1 U96 ( .A(\ALUOp2<12> ), .B(n10), .C(\WriteData<12> ), .D(n8), .Y(n97) );
  AOI22X1 U97 ( .A(\ALUOp2<11> ), .B(n10), .C(\WriteData<11> ), .D(n8), .Y(n98) );
  AOI22X1 U98 ( .A(\ALUOp2<10> ), .B(n10), .C(\WriteData<10> ), .D(n8), .Y(n99) );
  AOI22X1 U99 ( .A(\ALUOp2<0> ), .B(n10), .C(\WriteData<0> ), .D(n9), .Y(n100)
         );
  dff_215 \WriteReg_reg[0]  ( .q(\WriteReg_Out<0> ), .d(n75), .clk(clk), .rst(
        n12) );
  dff_216 \WriteReg_reg[1]  ( .q(\WriteReg_Out<1> ), .d(n76), .clk(clk), .rst(
        n12) );
  dff_217 \WriteReg_reg[2]  ( .q(\WriteReg_Out<2> ), .d(n78), .clk(clk), .rst(
        n12) );
  dff_212 \rs_reg[0]  ( .q(\Rs_Out<0> ), .d(n80), .clk(clk), .rst(n12) );
  dff_213 \rs_reg[1]  ( .q(\Rs_Out<1> ), .d(n81), .clk(clk), .rst(n12) );
  dff_214 \rs_reg[2]  ( .q(\Rs_Out<2> ), .d(n82), .clk(clk), .rst(n12) );
  dff_209 \rt_reg[0]  ( .q(\Rt_Out<0> ), .d(n83), .clk(clk), .rst(n12) );
  dff_210 \rt_reg[1]  ( .q(\Rt_Out<1> ), .d(n84), .clk(clk), .rst(n12) );
  dff_211 \rt_reg[2]  ( .q(\Rt_Out<2> ), .d(n101), .clk(clk), .rst(n12) );
  dff_206 \rd_reg[0]  ( .q(\Rd_Out<0> ), .d(n102), .clk(clk), .rst(n12) );
  dff_207 \rd_reg[1]  ( .q(\Rd_Out<1> ), .d(n103), .clk(clk), .rst(n12) );
  dff_208 \rd_reg[2]  ( .q(\Rd_Out<2> ), .d(n104), .clk(clk), .rst(n12) );
  dff_222 rf_wr_en_reg ( .q(RegFileWrEn_Out), .d(n79), .clk(clk), .rst(n12) );
  dff_190 \address_reg[0]  ( .q(\Address<0> ), .d(n42), .clk(clk), .rst(n11)
         );
  dff_191 \address_reg[1]  ( .q(\Address<1> ), .d(n74), .clk(clk), .rst(n12)
         );
  dff_192 \address_reg[2]  ( .q(n127), .d(n43), .clk(clk), .rst(n11) );
  dff_193 \address_reg[3]  ( .q(n126), .d(n44), .clk(clk), .rst(n11) );
  dff_194 \address_reg[4]  ( .q(n125), .d(n45), .clk(clk), .rst(n11) );
  dff_195 \address_reg[5]  ( .q(\Address<5> ), .d(n46), .clk(clk), .rst(n11)
         );
  dff_196 \address_reg[6]  ( .q(\Address<6> ), .d(n47), .clk(clk), .rst(n11)
         );
  dff_197 \address_reg[7]  ( .q(\Address<7> ), .d(n48), .clk(clk), .rst(n11)
         );
  dff_198 \address_reg[8]  ( .q(\Address<8> ), .d(n49), .clk(clk), .rst(n12)
         );
  dff_199 \address_reg[9]  ( .q(\Address<9> ), .d(n50), .clk(clk), .rst(n11)
         );
  dff_200 \address_reg[10]  ( .q(\Address<10> ), .d(n51), .clk(clk), .rst(n12)
         );
  dff_201 \address_reg[11]  ( .q(\Address<11> ), .d(n69), .clk(clk), .rst(n11)
         );
  dff_202 \address_reg[12]  ( .q(\Address<12> ), .d(n70), .clk(clk), .rst(n11)
         );
  dff_203 \address_reg[13]  ( .q(\Address<13> ), .d(n71), .clk(clk), .rst(n11)
         );
  dff_204 \address_reg[14]  ( .q(\Address<14> ), .d(n72), .clk(clk), .rst(n12)
         );
  dff_205 \address_reg[15]  ( .q(\Address<15> ), .d(n73), .clk(clk), .rst(n11)
         );
  dff_221 memread_reg ( .q(MemRead_Out), .d(n122), .clk(clk), .rst(n12) );
  dff_220 memwrite_reg ( .q(MemWrite_Out), .d(n121), .clk(clk), .rst(n12) );
  dff_219 memtoreg_reg ( .q(MemToReg_Out), .d(n123), .clk(clk), .rst(n12) );
  dff_174 \writedata_reg[0]  ( .q(\WriteData<0> ), .d(n105), .clk(clk), .rst(
        n12) );
  dff_175 \writedata_reg[1]  ( .q(\WriteData<1> ), .d(n106), .clk(clk), .rst(
        n12) );
  dff_176 \writedata_reg[2]  ( .q(\WriteData<2> ), .d(n107), .clk(clk), .rst(
        n12) );
  dff_177 \writedata_reg[3]  ( .q(\WriteData<3> ), .d(n108), .clk(clk), .rst(
        n12) );
  dff_178 \writedata_reg[4]  ( .q(\WriteData<4> ), .d(n109), .clk(clk), .rst(
        n12) );
  dff_179 \writedata_reg[5]  ( .q(\WriteData<5> ), .d(n110), .clk(clk), .rst(
        n12) );
  dff_180 \writedata_reg[6]  ( .q(\WriteData<6> ), .d(n111), .clk(clk), .rst(
        n12) );
  dff_181 \writedata_reg[7]  ( .q(\WriteData<7> ), .d(n112), .clk(clk), .rst(
        n12) );
  dff_182 \writedata_reg[8]  ( .q(\WriteData<8> ), .d(n113), .clk(clk), .rst(
        n12) );
  dff_183 \writedata_reg[9]  ( .q(\WriteData<9> ), .d(n114), .clk(clk), .rst(
        n12) );
  dff_184 \writedata_reg[10]  ( .q(\WriteData<10> ), .d(n115), .clk(clk), 
        .rst(n12) );
  dff_185 \writedata_reg[11]  ( .q(\WriteData<11> ), .d(n116), .clk(clk), 
        .rst(n12) );
  dff_186 \writedata_reg[12]  ( .q(\WriteData<12> ), .d(n117), .clk(clk), 
        .rst(n12) );
  dff_187 \writedata_reg[13]  ( .q(\WriteData<13> ), .d(n118), .clk(clk), 
        .rst(n12) );
  dff_188 \writedata_reg[14]  ( .q(\WriteData<14> ), .d(n119), .clk(clk), 
        .rst(n12) );
  dff_189 \writedata_reg[15]  ( .q(\WriteData<15> ), .d(n120), .clk(clk), 
        .rst(n12) );
  dff_218 halt_reg ( .q(Halt_Out), .d(n124), .clk(clk), .rst(n12) );
  INVX1 U1 ( .A(rst), .Y(n13) );
  INVX1 U2 ( .A(n13), .Y(n11) );
  INVX1 U3 ( .A(\Address<10> ), .Y(n24) );
  INVX1 U4 ( .A(n127), .Y(n2) );
  INVX1 U5 ( .A(n126), .Y(n4) );
  INVX1 U6 ( .A(n125), .Y(n6) );
  INVX1 U7 ( .A(\Address<5> ), .Y(n34) );
  INVX1 U8 ( .A(\Address<6> ), .Y(n32) );
  INVX1 U9 ( .A(\Address<7> ), .Y(n30) );
  INVX1 U10 ( .A(\Address<8> ), .Y(n28) );
  INVX1 U11 ( .A(\Address<9> ), .Y(n26) );
  INVX1 U12 ( .A(\Address<11> ), .Y(n22) );
  INVX1 U13 ( .A(\Address<12> ), .Y(n20) );
  INVX1 U14 ( .A(\Address<13> ), .Y(n18) );
  INVX1 U15 ( .A(\Address<14> ), .Y(n16) );
  INVX1 U16 ( .A(\Address<15> ), .Y(n14) );
  INVX1 U17 ( .A(n13), .Y(n12) );
  INVX1 U18 ( .A(n10), .Y(n7) );
  INVX1 U19 ( .A(Stall), .Y(n10) );
  INVX1 U20 ( .A(n77), .Y(n74) );
  INVX1 U21 ( .A(n100), .Y(n105) );
  INVX1 U22 ( .A(n99), .Y(n115) );
  INVX1 U23 ( .A(n98), .Y(n116) );
  INVX1 U24 ( .A(n97), .Y(n117) );
  INVX1 U25 ( .A(n96), .Y(n118) );
  INVX1 U26 ( .A(n95), .Y(n119) );
  INVX1 U27 ( .A(n94), .Y(n120) );
  INVX1 U28 ( .A(n93), .Y(n106) );
  INVX1 U29 ( .A(n92), .Y(n107) );
  INVX1 U30 ( .A(n91), .Y(n108) );
  INVX1 U31 ( .A(n90), .Y(n109) );
  INVX1 U32 ( .A(n89), .Y(n110) );
  INVX1 U33 ( .A(n88), .Y(n111) );
  INVX1 U34 ( .A(n87), .Y(n112) );
  INVX1 U35 ( .A(n86), .Y(n113) );
  INVX1 U36 ( .A(n85), .Y(n114) );
  INVX1 U37 ( .A(n10), .Y(n8) );
  INVX1 U38 ( .A(n68), .Y(n124) );
  INVX1 U39 ( .A(n67), .Y(n122) );
  INVX1 U40 ( .A(n66), .Y(n123) );
  INVX1 U41 ( .A(n65), .Y(n121) );
  INVX1 U42 ( .A(n64), .Y(n102) );
  INVX1 U43 ( .A(n63), .Y(n103) );
  INVX1 U44 ( .A(n62), .Y(n104) );
  INVX1 U45 ( .A(n61), .Y(n79) );
  INVX1 U46 ( .A(n60), .Y(n80) );
  INVX1 U47 ( .A(n59), .Y(n81) );
  INVX1 U48 ( .A(n58), .Y(n82) );
  INVX1 U49 ( .A(n57), .Y(n83) );
  INVX1 U50 ( .A(n56), .Y(n84) );
  INVX1 U68 ( .A(n55), .Y(n101) );
  INVX1 U69 ( .A(n54), .Y(n75) );
  INVX1 U70 ( .A(n53), .Y(n76) );
  INVX1 U71 ( .A(n52), .Y(n78) );
  INVX1 U72 ( .A(n10), .Y(n9) );
  INVX1 U73 ( .A(n2), .Y(\Address<2> ) );
  INVX1 U74 ( .A(n4), .Y(\Address<3> ) );
  INVX1 U75 ( .A(n6), .Y(\Address<4> ) );
  INVX1 U77 ( .A(\Result<2> ), .Y(n38) );
  INVX1 U78 ( .A(\Result<3> ), .Y(n37) );
  INVX1 U79 ( .A(\Result<4> ), .Y(n36) );
  INVX1 U80 ( .A(\Result<5> ), .Y(n35) );
  INVX1 U81 ( .A(\Result<6> ), .Y(n33) );
  INVX1 U82 ( .A(\Result<7> ), .Y(n31) );
  INVX1 U83 ( .A(\Result<8> ), .Y(n29) );
  INVX1 U100 ( .A(\Result<9> ), .Y(n27) );
  INVX1 U101 ( .A(\Result<10> ), .Y(n25) );
  INVX1 U102 ( .A(\Result<11> ), .Y(n23) );
  INVX1 U103 ( .A(\Result<12> ), .Y(n21) );
  INVX1 U104 ( .A(\Result<13> ), .Y(n19) );
  INVX1 U105 ( .A(\Result<14> ), .Y(n17) );
  INVX1 U106 ( .A(\Result<15> ), .Y(n15) );
  INVX1 U107 ( .A(\Result<0> ), .Y(n41) );
  MUX2X1 U108 ( .B(n15), .A(n14), .S(n7), .Y(n73) );
  MUX2X1 U109 ( .B(n17), .A(n16), .S(n7), .Y(n72) );
  MUX2X1 U110 ( .B(n19), .A(n18), .S(n7), .Y(n71) );
  MUX2X1 U111 ( .B(n21), .A(n20), .S(n7), .Y(n70) );
  MUX2X1 U112 ( .B(n23), .A(n22), .S(n7), .Y(n69) );
  MUX2X1 U113 ( .B(n25), .A(n24), .S(n7), .Y(n51) );
  MUX2X1 U114 ( .B(n27), .A(n26), .S(n7), .Y(n50) );
  MUX2X1 U115 ( .B(n29), .A(n28), .S(n7), .Y(n49) );
  MUX2X1 U116 ( .B(n31), .A(n30), .S(n7), .Y(n48) );
  MUX2X1 U117 ( .B(n33), .A(n32), .S(n7), .Y(n47) );
  MUX2X1 U118 ( .B(n35), .A(n34), .S(n7), .Y(n46) );
  MUX2X1 U119 ( .B(n36), .A(n6), .S(n7), .Y(n45) );
  MUX2X1 U120 ( .B(n37), .A(n4), .S(n8), .Y(n44) );
  MUX2X1 U121 ( .B(n38), .A(n2), .S(n8), .Y(n43) );
  NAND2X1 U122 ( .A(\Address<0> ), .B(n7), .Y(n40) );
  AND2X2 U123 ( .A(n7), .B(n40), .Y(n39) );
  AOI21X1 U124 ( .A(n41), .B(n40), .C(n39), .Y(n42) );
endmodule


module memory ( MemRead, MemWrite, halt, clk, rst, .Address({\Address<15> , 
        \Address<14> , \Address<13> , \Address<12> , \Address<11> , 
        \Address<10> , \Address<9> , \Address<8> , \Address<7> , \Address<6> , 
        \Address<5> , \Address<4> , \Address<3> , \Address<2> , \Address<1> , 
        \Address<0> }), .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .ReadData({\ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }), Err, DataMemStall, 
        CacheHit );
  input MemRead, MemWrite, halt, clk, rst, \Address<15> , \Address<14> ,
         \Address<13> , \Address<12> , \Address<11> , \Address<10> ,
         \Address<9> , \Address<8> , \Address<7> , \Address<6> , \Address<5> ,
         \Address<4> , \Address<3> , \Address<2> , \Address<1> , \Address<0> ,
         \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ;
  output \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> ,
         \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> ,
         \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> ,
         \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> , Err,
         DataMemStall, CacheHit;
  wire   n2;
  assign CacheHit = 1'b0;

  stallmem data_mem ( .DataOut({\ReadData<15> , \ReadData<14> , \ReadData<13> , 
        \ReadData<12> , \ReadData<11> , \ReadData<10> , \ReadData<9> , 
        \ReadData<8> , \ReadData<7> , \ReadData<6> , \ReadData<5> , 
        \ReadData<4> , \ReadData<3> , \ReadData<2> , \ReadData<1> , 
        \ReadData<0> }), .Done(), .Stall(DataMemStall), .CacheHit(), .err(n2), 
        .Addr({\Address<15> , \Address<14> , \Address<13> , \Address<12> , 
        \Address<11> , \Address<10> , \Address<9> , \Address<8> , \Address<7> , 
        \Address<6> , \Address<5> , \Address<4> , \Address<3> , \Address<2> , 
        \Address<1> , \Address<0> }), .DataIn({\WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .Rd(MemRead), .Wr(
        MemWrite), .createdump(halt), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(n2), .Y(Err) );
endmodule


module pipe_mw ( Stall, rst, clk, .ExecuteOut({\ExecuteOut<15> , 
        \ExecuteOut<14> , \ExecuteOut<13> , \ExecuteOut<12> , \ExecuteOut<11> , 
        \ExecuteOut<10> , \ExecuteOut<9> , \ExecuteOut<8> , \ExecuteOut<7> , 
        \ExecuteOut<6> , \ExecuteOut<5> , \ExecuteOut<4> , \ExecuteOut<3> , 
        \ExecuteOut<2> , \ExecuteOut<1> , \ExecuteOut<0> }), .MemOut({
        \MemOut<15> , \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> , 
        \MemOut<10> , \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> , 
        \MemOut<5> , \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> , 
        \MemOut<0> }), MemToReg, RegFileWrEn, .Rs({\Rs<2> , \Rs<1> , \Rs<0> }), 
    .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({\Rd<2> , \Rd<1> , \Rd<0> }), 
    .WriteReg({\WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), 
    .ExecuteOut_Out({\ExecuteOut_Out<15> , \ExecuteOut_Out<14> , 
        \ExecuteOut_Out<13> , \ExecuteOut_Out<12> , \ExecuteOut_Out<11> , 
        \ExecuteOut_Out<10> , \ExecuteOut_Out<9> , \ExecuteOut_Out<8> , 
        \ExecuteOut_Out<7> , \ExecuteOut_Out<6> , \ExecuteOut_Out<5> , 
        \ExecuteOut_Out<4> , \ExecuteOut_Out<3> , \ExecuteOut_Out<2> , 
        \ExecuteOut_Out<1> , \ExecuteOut_Out<0> }), .MemOut_Out({
        \MemOut_Out<15> , \MemOut_Out<14> , \MemOut_Out<13> , \MemOut_Out<12> , 
        \MemOut_Out<11> , \MemOut_Out<10> , \MemOut_Out<9> , \MemOut_Out<8> , 
        \MemOut_Out<7> , \MemOut_Out<6> , \MemOut_Out<5> , \MemOut_Out<4> , 
        \MemOut_Out<3> , \MemOut_Out<2> , \MemOut_Out<1> , \MemOut_Out<0> }), 
        MemToReg_Out, RegFileWrEn_Out, .WriteReg_Out({\WriteReg_Out<2> , 
        \WriteReg_Out<1> , \WriteReg_Out<0> }), .Rs_Out({\Rs_Out<2> , 
        \Rs_Out<1> , \Rs_Out<0> }), .Rt_Out({\Rt_Out<2> , \Rt_Out<1> , 
        \Rt_Out<0> }), .Rd_Out({\Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> }) );
  input Stall, rst, clk, \ExecuteOut<15> , \ExecuteOut<14> , \ExecuteOut<13> ,
         \ExecuteOut<12> , \ExecuteOut<11> , \ExecuteOut<10> , \ExecuteOut<9> ,
         \ExecuteOut<8> , \ExecuteOut<7> , \ExecuteOut<6> , \ExecuteOut<5> ,
         \ExecuteOut<4> , \ExecuteOut<3> , \ExecuteOut<2> , \ExecuteOut<1> ,
         \ExecuteOut<0> , \MemOut<15> , \MemOut<14> , \MemOut<13> ,
         \MemOut<12> , \MemOut<11> , \MemOut<10> , \MemOut<9> , \MemOut<8> ,
         \MemOut<7> , \MemOut<6> , \MemOut<5> , \MemOut<4> , \MemOut<3> ,
         \MemOut<2> , \MemOut<1> , \MemOut<0> , MemToReg, RegFileWrEn, \Rs<2> ,
         \Rs<1> , \Rs<0> , \Rt<2> , \Rt<1> , \Rt<0> , \Rd<2> , \Rd<1> ,
         \Rd<0> , \WriteReg<2> , \WriteReg<1> , \WriteReg<0> ;
  output \ExecuteOut_Out<15> , \ExecuteOut_Out<14> , \ExecuteOut_Out<13> ,
         \ExecuteOut_Out<12> , \ExecuteOut_Out<11> , \ExecuteOut_Out<10> ,
         \ExecuteOut_Out<9> , \ExecuteOut_Out<8> , \ExecuteOut_Out<7> ,
         \ExecuteOut_Out<6> , \ExecuteOut_Out<5> , \ExecuteOut_Out<4> ,
         \ExecuteOut_Out<3> , \ExecuteOut_Out<2> , \ExecuteOut_Out<1> ,
         \ExecuteOut_Out<0> , \MemOut_Out<15> , \MemOut_Out<14> ,
         \MemOut_Out<13> , \MemOut_Out<12> , \MemOut_Out<11> ,
         \MemOut_Out<10> , \MemOut_Out<9> , \MemOut_Out<8> , \MemOut_Out<7> ,
         \MemOut_Out<6> , \MemOut_Out<5> , \MemOut_Out<4> , \MemOut_Out<3> ,
         \MemOut_Out<2> , \MemOut_Out<1> , \MemOut_Out<0> , MemToReg_Out,
         RegFileWrEn_Out, \WriteReg_Out<2> , \WriteReg_Out<1> ,
         \WriteReg_Out<0> , \Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> , \Rt_Out<2> ,
         \Rt_Out<1> , \Rt_Out<0> , \Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> ;
  wire   n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n95, n96, n97;

  AOI22X1 U48 ( .A(\WriteReg<2> ), .B(n97), .C(\WriteReg_Out<2> ), .D(Stall), 
        .Y(n49) );
  AOI22X1 U49 ( .A(\WriteReg<1> ), .B(n97), .C(\WriteReg_Out<1> ), .D(Stall), 
        .Y(n50) );
  AOI22X1 U50 ( .A(\WriteReg<0> ), .B(n97), .C(\WriteReg_Out<0> ), .D(Stall), 
        .Y(n51) );
  AOI22X1 U51 ( .A(\Rt<2> ), .B(n97), .C(\Rt_Out<2> ), .D(Stall), .Y(n52) );
  AOI22X1 U52 ( .A(\Rt<1> ), .B(n97), .C(\Rt_Out<1> ), .D(Stall), .Y(n53) );
  AOI22X1 U53 ( .A(\Rt<0> ), .B(n97), .C(\Rt_Out<0> ), .D(Stall), .Y(n54) );
  AOI22X1 U54 ( .A(\Rs<2> ), .B(n97), .C(\Rs_Out<2> ), .D(Stall), .Y(n55) );
  AOI22X1 U55 ( .A(\Rs<1> ), .B(n97), .C(\Rs_Out<1> ), .D(Stall), .Y(n56) );
  AOI22X1 U56 ( .A(\Rs<0> ), .B(n97), .C(\Rs_Out<0> ), .D(Stall), .Y(n57) );
  AOI22X1 U57 ( .A(RegFileWrEn), .B(n97), .C(RegFileWrEn_Out), .D(Stall), .Y(
        n58) );
  AOI22X1 U58 ( .A(\Rd<2> ), .B(n97), .C(\Rd_Out<2> ), .D(Stall), .Y(n59) );
  AOI22X1 U59 ( .A(\Rd<1> ), .B(n97), .C(\Rd_Out<1> ), .D(Stall), .Y(n60) );
  AOI22X1 U60 ( .A(\Rd<0> ), .B(n97), .C(\Rd_Out<0> ), .D(Stall), .Y(n61) );
  AOI22X1 U61 ( .A(MemToReg), .B(n97), .C(MemToReg_Out), .D(Stall), .Y(n62) );
  AOI22X1 U62 ( .A(\MemOut<9> ), .B(n97), .C(\MemOut_Out<9> ), .D(Stall), .Y(
        n63) );
  AOI22X1 U63 ( .A(\MemOut<8> ), .B(n97), .C(\MemOut_Out<8> ), .D(Stall), .Y(
        n64) );
  AOI22X1 U64 ( .A(\MemOut<7> ), .B(n97), .C(\MemOut_Out<7> ), .D(Stall), .Y(
        n65) );
  AOI22X1 U65 ( .A(\MemOut<6> ), .B(n97), .C(\MemOut_Out<6> ), .D(Stall), .Y(
        n66) );
  AOI22X1 U66 ( .A(\MemOut<5> ), .B(n97), .C(\MemOut_Out<5> ), .D(Stall), .Y(
        n67) );
  AOI22X1 U67 ( .A(\MemOut<4> ), .B(n97), .C(\MemOut_Out<4> ), .D(Stall), .Y(
        n68) );
  AOI22X1 U68 ( .A(\MemOut<3> ), .B(n97), .C(\MemOut_Out<3> ), .D(Stall), .Y(
        n69) );
  AOI22X1 U69 ( .A(\MemOut<2> ), .B(n97), .C(\MemOut_Out<2> ), .D(Stall), .Y(
        n70) );
  AOI22X1 U70 ( .A(\MemOut<1> ), .B(n97), .C(\MemOut_Out<1> ), .D(Stall), .Y(
        n71) );
  AOI22X1 U71 ( .A(\MemOut<15> ), .B(n97), .C(\MemOut_Out<15> ), .D(Stall), 
        .Y(n72) );
  AOI22X1 U72 ( .A(\MemOut<14> ), .B(n97), .C(\MemOut_Out<14> ), .D(Stall), 
        .Y(n73) );
  AOI22X1 U73 ( .A(\MemOut<13> ), .B(n97), .C(\MemOut_Out<13> ), .D(Stall), 
        .Y(n74) );
  AOI22X1 U74 ( .A(\MemOut<12> ), .B(n97), .C(\MemOut_Out<12> ), .D(Stall), 
        .Y(n75) );
  AOI22X1 U75 ( .A(\MemOut<11> ), .B(n97), .C(\MemOut_Out<11> ), .D(Stall), 
        .Y(n76) );
  AOI22X1 U76 ( .A(\MemOut<10> ), .B(n97), .C(\MemOut_Out<10> ), .D(Stall), 
        .Y(n77) );
  AOI22X1 U77 ( .A(\MemOut<0> ), .B(n97), .C(\MemOut_Out<0> ), .D(Stall), .Y(
        n78) );
  AOI22X1 U78 ( .A(\ExecuteOut<9> ), .B(n97), .C(\ExecuteOut_Out<9> ), .D(
        Stall), .Y(n79) );
  AOI22X1 U79 ( .A(\ExecuteOut<8> ), .B(n97), .C(\ExecuteOut_Out<8> ), .D(
        Stall), .Y(n80) );
  AOI22X1 U80 ( .A(\ExecuteOut<7> ), .B(n97), .C(\ExecuteOut_Out<7> ), .D(
        Stall), .Y(n81) );
  AOI22X1 U81 ( .A(\ExecuteOut<6> ), .B(n97), .C(\ExecuteOut_Out<6> ), .D(
        Stall), .Y(n82) );
  AOI22X1 U82 ( .A(\ExecuteOut<5> ), .B(n97), .C(\ExecuteOut_Out<5> ), .D(
        Stall), .Y(n83) );
  AOI22X1 U83 ( .A(\ExecuteOut<4> ), .B(n97), .C(\ExecuteOut_Out<4> ), .D(
        Stall), .Y(n84) );
  AOI22X1 U84 ( .A(\ExecuteOut<3> ), .B(n97), .C(\ExecuteOut_Out<3> ), .D(
        Stall), .Y(n85) );
  AOI22X1 U85 ( .A(\ExecuteOut<2> ), .B(n97), .C(\ExecuteOut_Out<2> ), .D(
        Stall), .Y(n86) );
  AOI22X1 U86 ( .A(\ExecuteOut<1> ), .B(n97), .C(\ExecuteOut_Out<1> ), .D(
        Stall), .Y(n87) );
  AOI22X1 U87 ( .A(\ExecuteOut<15> ), .B(n97), .C(\ExecuteOut_Out<15> ), .D(
        Stall), .Y(n88) );
  AOI22X1 U88 ( .A(\ExecuteOut<14> ), .B(n97), .C(\ExecuteOut_Out<14> ), .D(
        Stall), .Y(n89) );
  AOI22X1 U89 ( .A(\ExecuteOut<13> ), .B(n97), .C(\ExecuteOut_Out<13> ), .D(
        Stall), .Y(n90) );
  AOI22X1 U90 ( .A(\ExecuteOut<12> ), .B(n97), .C(\ExecuteOut_Out<12> ), .D(
        Stall), .Y(n91) );
  AOI22X1 U91 ( .A(\ExecuteOut<11> ), .B(n97), .C(\ExecuteOut_Out<11> ), .D(
        Stall), .Y(n92) );
  AOI22X1 U92 ( .A(\ExecuteOut<10> ), .B(n97), .C(\ExecuteOut_Out<10> ), .D(
        Stall), .Y(n93) );
  AOI22X1 U93 ( .A(\ExecuteOut<0> ), .B(n97), .C(\ExecuteOut_Out<0> ), .D(
        Stall), .Y(n94) );
  dff_169 \WriteReg_reg[0]  ( .q(\WriteReg_Out<0> ), .d(n5), .clk(clk), .rst(
        n3) );
  dff_170 \WriteReg_reg[1]  ( .q(\WriteReg_Out<1> ), .d(n6), .clk(clk), .rst(
        n3) );
  dff_171 \WriteReg_reg[2]  ( .q(\WriteReg_Out<2> ), .d(n7), .clk(clk), .rst(
        n3) );
  dff_166 \rs_reg[0]  ( .q(\Rs_Out<0> ), .d(n8), .clk(clk), .rst(n3) );
  dff_167 \rs_reg[1]  ( .q(\Rs_Out<1> ), .d(n9), .clk(clk), .rst(n3) );
  dff_168 \rs_reg[2]  ( .q(\Rs_Out<2> ), .d(n10), .clk(clk), .rst(n3) );
  dff_163 \rt_reg[0]  ( .q(\Rt_Out<0> ), .d(n11), .clk(clk), .rst(n3) );
  dff_164 \rt_reg[1]  ( .q(\Rt_Out<1> ), .d(n12), .clk(clk), .rst(n2) );
  dff_165 \rt_reg[2]  ( .q(\Rt_Out<2> ), .d(n13), .clk(clk), .rst(n2) );
  dff_160 \rd_reg[0]  ( .q(\Rd_Out<0> ), .d(n14), .clk(clk), .rst(n2) );
  dff_161 \rd_reg[1]  ( .q(\Rd_Out<1> ), .d(n15), .clk(clk), .rst(n2) );
  dff_162 \rd_reg[2]  ( .q(\Rd_Out<2> ), .d(n16), .clk(clk), .rst(n2) );
  dff_173 rf_wr_en_reg ( .q(RegFileWrEn_Out), .d(n17), .clk(clk), .rst(n2) );
  dff_144 \executeout_reg[0]  ( .q(\ExecuteOut_Out<0> ), .d(n18), .clk(clk), 
        .rst(n2) );
  dff_145 \executeout_reg[1]  ( .q(\ExecuteOut_Out<1> ), .d(n35), .clk(clk), 
        .rst(n2) );
  dff_146 \executeout_reg[2]  ( .q(\ExecuteOut_Out<2> ), .d(n36), .clk(clk), 
        .rst(n2) );
  dff_147 \executeout_reg[3]  ( .q(\ExecuteOut_Out<3> ), .d(n37), .clk(clk), 
        .rst(n2) );
  dff_148 \executeout_reg[4]  ( .q(\ExecuteOut_Out<4> ), .d(n38), .clk(clk), 
        .rst(n2) );
  dff_149 \executeout_reg[5]  ( .q(\ExecuteOut_Out<5> ), .d(n39), .clk(clk), 
        .rst(n2) );
  dff_150 \executeout_reg[6]  ( .q(\ExecuteOut_Out<6> ), .d(n40), .clk(clk), 
        .rst(n2) );
  dff_151 \executeout_reg[7]  ( .q(\ExecuteOut_Out<7> ), .d(n41), .clk(clk), 
        .rst(n1) );
  dff_152 \executeout_reg[8]  ( .q(\ExecuteOut_Out<8> ), .d(n42), .clk(clk), 
        .rst(n1) );
  dff_153 \executeout_reg[9]  ( .q(\ExecuteOut_Out<9> ), .d(n43), .clk(clk), 
        .rst(n1) );
  dff_154 \executeout_reg[10]  ( .q(\ExecuteOut_Out<10> ), .d(n44), .clk(clk), 
        .rst(n1) );
  dff_155 \executeout_reg[11]  ( .q(\ExecuteOut_Out<11> ), .d(n45), .clk(clk), 
        .rst(n1) );
  dff_156 \executeout_reg[12]  ( .q(\ExecuteOut_Out<12> ), .d(n46), .clk(clk), 
        .rst(n1) );
  dff_157 \executeout_reg[13]  ( .q(\ExecuteOut_Out<13> ), .d(n47), .clk(clk), 
        .rst(n1) );
  dff_158 \executeout_reg[14]  ( .q(\ExecuteOut_Out<14> ), .d(n48), .clk(clk), 
        .rst(n1) );
  dff_159 \executeout_reg[15]  ( .q(\ExecuteOut_Out<15> ), .d(n95), .clk(clk), 
        .rst(n1) );
  dff_128 \memout_reg[0]  ( .q(\MemOut_Out<0> ), .d(n34), .clk(clk), .rst(n1)
         );
  dff_129 \memout_reg[1]  ( .q(\MemOut_Out<1> ), .d(n32), .clk(clk), .rst(n1)
         );
  dff_130 \memout_reg[2]  ( .q(\MemOut_Out<2> ), .d(n29), .clk(clk), .rst(n1)
         );
  dff_131 \memout_reg[3]  ( .q(\MemOut_Out<3> ), .d(n27), .clk(clk), .rst(n1)
         );
  dff_132 \memout_reg[4]  ( .q(\MemOut_Out<4> ), .d(n25), .clk(clk), .rst(n3)
         );
  dff_133 \memout_reg[5]  ( .q(\MemOut_Out<5> ), .d(n23), .clk(clk), .rst(n3)
         );
  dff_134 \memout_reg[6]  ( .q(\MemOut_Out<6> ), .d(n21), .clk(clk), .rst(n3)
         );
  dff_135 \memout_reg[7]  ( .q(\MemOut_Out<7> ), .d(n19), .clk(clk), .rst(n3)
         );
  dff_136 \memout_reg[8]  ( .q(\MemOut_Out<8> ), .d(n33), .clk(clk), .rst(n3)
         );
  dff_137 \memout_reg[9]  ( .q(\MemOut_Out<9> ), .d(n31), .clk(clk), .rst(n3)
         );
  dff_138 \memout_reg[10]  ( .q(\MemOut_Out<10> ), .d(n30), .clk(clk), .rst(
        rst) );
  dff_139 \memout_reg[11]  ( .q(\MemOut_Out<11> ), .d(n28), .clk(clk), .rst(
        rst) );
  dff_140 \memout_reg[12]  ( .q(\MemOut_Out<12> ), .d(n26), .clk(clk), .rst(
        rst) );
  dff_141 \memout_reg[13]  ( .q(\MemOut_Out<13> ), .d(n24), .clk(clk), .rst(
        rst) );
  dff_142 \memout_reg[14]  ( .q(\MemOut_Out<14> ), .d(n22), .clk(clk), .rst(
        rst) );
  dff_143 \memout_reg[15]  ( .q(\MemOut_Out<15> ), .d(n20), .clk(clk), .rst(
        rst) );
  dff_172 memtoreg_reg ( .q(MemToReg_Out), .d(n96), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(Stall), .Y(n97) );
  INVX1 U2 ( .A(rst), .Y(n4) );
  INVX1 U3 ( .A(n4), .Y(n1) );
  INVX1 U4 ( .A(n4), .Y(n2) );
  INVX1 U5 ( .A(n4), .Y(n3) );
  INVX1 U6 ( .A(n94), .Y(n18) );
  INVX1 U7 ( .A(n93), .Y(n44) );
  INVX1 U8 ( .A(n92), .Y(n45) );
  INVX1 U9 ( .A(n91), .Y(n46) );
  INVX1 U10 ( .A(n90), .Y(n47) );
  INVX1 U11 ( .A(n89), .Y(n48) );
  INVX1 U12 ( .A(n88), .Y(n95) );
  INVX1 U13 ( .A(n87), .Y(n35) );
  INVX1 U14 ( .A(n86), .Y(n36) );
  INVX1 U15 ( .A(n85), .Y(n37) );
  INVX1 U16 ( .A(n84), .Y(n38) );
  INVX1 U17 ( .A(n83), .Y(n39) );
  INVX1 U18 ( .A(n82), .Y(n40) );
  INVX1 U19 ( .A(n81), .Y(n41) );
  INVX1 U20 ( .A(n80), .Y(n42) );
  INVX1 U21 ( .A(n79), .Y(n43) );
  INVX1 U22 ( .A(n78), .Y(n34) );
  INVX1 U23 ( .A(n77), .Y(n30) );
  INVX1 U24 ( .A(n76), .Y(n28) );
  INVX1 U25 ( .A(n75), .Y(n26) );
  INVX1 U26 ( .A(n74), .Y(n24) );
  INVX1 U27 ( .A(n73), .Y(n22) );
  INVX1 U28 ( .A(n72), .Y(n20) );
  INVX1 U29 ( .A(n71), .Y(n32) );
  INVX1 U30 ( .A(n70), .Y(n29) );
  INVX1 U31 ( .A(n69), .Y(n27) );
  INVX1 U32 ( .A(n68), .Y(n25) );
  INVX1 U33 ( .A(n67), .Y(n23) );
  INVX1 U34 ( .A(n66), .Y(n21) );
  INVX1 U35 ( .A(n65), .Y(n19) );
  INVX1 U36 ( .A(n64), .Y(n33) );
  INVX1 U37 ( .A(n63), .Y(n31) );
  INVX1 U38 ( .A(n62), .Y(n96) );
  INVX1 U39 ( .A(n61), .Y(n14) );
  INVX1 U40 ( .A(n60), .Y(n15) );
  INVX1 U41 ( .A(n59), .Y(n16) );
  INVX1 U42 ( .A(n58), .Y(n17) );
  INVX1 U43 ( .A(n57), .Y(n8) );
  INVX1 U44 ( .A(n56), .Y(n9) );
  INVX1 U45 ( .A(n55), .Y(n10) );
  INVX1 U46 ( .A(n54), .Y(n11) );
  INVX1 U47 ( .A(n53), .Y(n12) );
  INVX1 U94 ( .A(n52), .Y(n13) );
  INVX1 U95 ( .A(n51), .Y(n5) );
  INVX1 U96 ( .A(n50), .Y(n6) );
  INVX1 U97 ( .A(n49), .Y(n7) );
endmodule


module writeback ( .ExecuteOut({\ExecuteOut<15> , \ExecuteOut<14> , 
        \ExecuteOut<13> , \ExecuteOut<12> , \ExecuteOut<11> , \ExecuteOut<10> , 
        \ExecuteOut<9> , \ExecuteOut<8> , \ExecuteOut<7> , \ExecuteOut<6> , 
        \ExecuteOut<5> , \ExecuteOut<4> , \ExecuteOut<3> , \ExecuteOut<2> , 
        \ExecuteOut<1> , \ExecuteOut<0> }), .MemOut({\MemOut<15> , 
        \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> , \MemOut<10> , 
        \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> , \MemOut<5> , 
        \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> , \MemOut<0> }), 
        MemToReg, .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }) );
  input \ExecuteOut<15> , \ExecuteOut<14> , \ExecuteOut<13> , \ExecuteOut<12> ,
         \ExecuteOut<11> , \ExecuteOut<10> , \ExecuteOut<9> , \ExecuteOut<8> ,
         \ExecuteOut<7> , \ExecuteOut<6> , \ExecuteOut<5> , \ExecuteOut<4> ,
         \ExecuteOut<3> , \ExecuteOut<2> , \ExecuteOut<1> , \ExecuteOut<0> ,
         \MemOut<15> , \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> ,
         \MemOut<10> , \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> ,
         \MemOut<5> , \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> ,
         \MemOut<0> , MemToReg;
  output \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n17;

  AOI22X1 U18 ( .A(\ExecuteOut<9> ), .B(n17), .C(MemToReg), .D(\MemOut<9> ), 
        .Y(n19) );
  AOI22X1 U19 ( .A(\ExecuteOut<8> ), .B(n17), .C(\MemOut<8> ), .D(MemToReg), 
        .Y(n20) );
  AOI22X1 U20 ( .A(\ExecuteOut<7> ), .B(n17), .C(\MemOut<7> ), .D(MemToReg), 
        .Y(n21) );
  AOI22X1 U21 ( .A(\ExecuteOut<6> ), .B(n17), .C(\MemOut<6> ), .D(MemToReg), 
        .Y(n22) );
  AOI22X1 U22 ( .A(\ExecuteOut<5> ), .B(n17), .C(\MemOut<5> ), .D(MemToReg), 
        .Y(n23) );
  AOI22X1 U23 ( .A(\ExecuteOut<4> ), .B(n17), .C(\MemOut<4> ), .D(MemToReg), 
        .Y(n24) );
  AOI22X1 U24 ( .A(\ExecuteOut<3> ), .B(n17), .C(\MemOut<3> ), .D(MemToReg), 
        .Y(n25) );
  AOI22X1 U25 ( .A(\ExecuteOut<2> ), .B(n17), .C(\MemOut<2> ), .D(MemToReg), 
        .Y(n26) );
  AOI22X1 U26 ( .A(\ExecuteOut<1> ), .B(n17), .C(\MemOut<1> ), .D(MemToReg), 
        .Y(n27) );
  AOI22X1 U27 ( .A(\ExecuteOut<15> ), .B(n17), .C(\MemOut<15> ), .D(MemToReg), 
        .Y(n28) );
  AOI22X1 U28 ( .A(\ExecuteOut<14> ), .B(n17), .C(\MemOut<14> ), .D(MemToReg), 
        .Y(n29) );
  AOI22X1 U29 ( .A(\ExecuteOut<13> ), .B(n17), .C(\MemOut<13> ), .D(MemToReg), 
        .Y(n30) );
  AOI22X1 U30 ( .A(\ExecuteOut<12> ), .B(n17), .C(\MemOut<12> ), .D(MemToReg), 
        .Y(n31) );
  AOI22X1 U31 ( .A(\ExecuteOut<11> ), .B(n17), .C(\MemOut<11> ), .D(MemToReg), 
        .Y(n32) );
  AOI22X1 U32 ( .A(\ExecuteOut<10> ), .B(n17), .C(\MemOut<10> ), .D(MemToReg), 
        .Y(n33) );
  AOI22X1 U33 ( .A(\ExecuteOut<0> ), .B(n17), .C(\MemOut<0> ), .D(MemToReg), 
        .Y(n34) );
  INVX1 U1 ( .A(n34), .Y(\WriteData<0> ) );
  INVX1 U2 ( .A(n33), .Y(\WriteData<10> ) );
  INVX1 U3 ( .A(n32), .Y(\WriteData<11> ) );
  INVX1 U4 ( .A(n31), .Y(\WriteData<12> ) );
  INVX1 U5 ( .A(n30), .Y(\WriteData<13> ) );
  INVX1 U6 ( .A(n29), .Y(\WriteData<14> ) );
  INVX1 U7 ( .A(n28), .Y(\WriteData<15> ) );
  INVX1 U8 ( .A(n27), .Y(\WriteData<1> ) );
  INVX1 U9 ( .A(n26), .Y(\WriteData<2> ) );
  INVX1 U10 ( .A(n25), .Y(\WriteData<3> ) );
  INVX1 U11 ( .A(n24), .Y(\WriteData<4> ) );
  INVX1 U12 ( .A(n23), .Y(\WriteData<5> ) );
  INVX1 U13 ( .A(n22), .Y(\WriteData<6> ) );
  INVX1 U14 ( .A(n21), .Y(\WriteData<7> ) );
  INVX1 U15 ( .A(n20), .Y(\WriteData<8> ) );
  INVX1 U16 ( .A(n19), .Y(\WriteData<9> ) );
  INVX1 U17 ( .A(MemToReg), .Y(n17) );
endmodule


module proc ( err, clk, rst );
  input clk, rst;
  output err;
  wire   M_Err, E_BranchJumpTaken, M_DataMemStall, D_RsValid, PDE_RegFileWrEn,
         \PDE_WriteReg<2> , \PDE_WriteReg<1> , \PDE_WriteReg<0> , \D_Rs<2> ,
         \D_Rs<1> , \D_Rs<0> , D_RtValid, \D_Rt<2> , \D_Rt<1> , \D_Rt<0> ,
         PEM_RegFileWrEn, \PEM_WriteReg<2> , \PEM_WriteReg<1> ,
         \PEM_WriteReg<0> , D_RdValid, D_Store, \D_Rd<2> , \D_Rd<1> ,
         \D_Rd<0> , \E_BranchPC<15> , \E_BranchPC<14> , \E_BranchPC<13> ,
         \E_BranchPC<12> , \E_BranchPC<11> , \E_BranchPC<10> , \E_BranchPC<9> ,
         \E_BranchPC<8> , \E_BranchPC<7> , \E_BranchPC<6> , \E_BranchPC<5> ,
         \E_BranchPC<4> , \E_BranchPC<3> , \E_BranchPC<2> , \E_BranchPC<1> ,
         \E_BranchPC<0> , PEM_Halt, D_Exception, D_Rti, \F_Instr<15> ,
         \F_Instr<14> , \F_Instr<13> , \F_Instr<12> , \F_Instr<11> ,
         \F_Instr<10> , \F_Instr<9> , \F_Instr<8> , \F_Instr<7> , \F_Instr<6> ,
         \F_Instr<5> , \F_Instr<4> , \F_Instr<3> , \F_Instr<2> , \F_Instr<1> ,
         \F_Instr<0> , \F_IncPC<15> , \F_IncPC<14> , \F_IncPC<13> ,
         \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , \F_IncPC<9> ,
         \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , \F_IncPC<4> ,
         \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> ,
         \PFD_Instr<15> , \PFD_Instr<14> , \PFD_Instr<13> , \PFD_Instr<12> ,
         \PFD_Instr<11> , \PFD_Instr<10> , \PFD_Instr<9> , \PFD_Instr<8> ,
         \PFD_Instr<7> , \PFD_Instr<6> , \PFD_Instr<5> , \PFD_Instr<4> ,
         \PFD_Instr<3> , \PFD_Instr<2> , \PFD_Instr<1> , \PFD_Instr<0> ,
         \PFD_IncPC<15> , \PFD_IncPC<14> , \PFD_IncPC<13> , \PFD_IncPC<12> ,
         \PFD_IncPC<11> , \PFD_IncPC<10> , \PFD_IncPC<9> , \PFD_IncPC<8> ,
         \PFD_IncPC<7> , \PFD_IncPC<6> , \PFD_IncPC<5> , \PFD_IncPC<4> ,
         \PFD_IncPC<3> , \PFD_IncPC<2> , \PFD_IncPC<1> , \PFD_IncPC<0> ,
         PFD_CPUActive, _3_net_, \W_WriteData<15> , \W_WriteData<14> ,
         \W_WriteData<13> , \W_WriteData<12> , \W_WriteData<11> ,
         \W_WriteData<10> , \W_WriteData<9> , \W_WriteData<8> ,
         \W_WriteData<7> , \W_WriteData<6> , \W_WriteData<5> ,
         \W_WriteData<4> , \W_WriteData<3> , \W_WriteData<2> ,
         \W_WriteData<1> , \W_WriteData<0> , \D_ALUOp1<15> , \D_ALUOp1<14> ,
         \D_ALUOp1<13> , \D_ALUOp1<12> , \D_ALUOp1<11> , \D_ALUOp1<10> ,
         \D_ALUOp1<9> , \D_ALUOp1<8> , \D_ALUOp1<7> , \D_ALUOp1<6> ,
         \D_ALUOp1<5> , \D_ALUOp1<4> , \D_ALUOp1<3> , \D_ALUOp1<2> ,
         \D_ALUOp1<1> , \D_ALUOp1<0> , \D_ALUOp2<15> , \D_ALUOp2<14> ,
         \D_ALUOp2<13> , \D_ALUOp2<12> , \D_ALUOp2<11> , \D_ALUOp2<10> ,
         \D_ALUOp2<9> , \D_ALUOp2<8> , \D_ALUOp2<7> , \D_ALUOp2<6> ,
         \D_ALUOp2<5> , \D_ALUOp2<4> , \D_ALUOp2<3> , \D_ALUOp2<2> ,
         \D_ALUOp2<1> , \D_ALUOp2<0> , D_ALUSrc, D_Branch, D_Jump, D_JumpReg,
         D_Set, D_Btr, \D_ALUOpcode<2> , \D_ALUOpcode<1> , \D_ALUOpcode<0> ,
         \D_Func<1> , \D_Func<0> , D_MemWrite, D_MemRead, D_MemToReg, D_Halt,
         \D_Immediate<15> , \D_Immediate<14> , \D_Immediate<13> ,
         \D_Immediate<12> , \D_Immediate<11> , \D_Immediate<10> ,
         \D_Immediate<9> , \D_Immediate<8> , \D_Immediate<7> ,
         \D_Immediate<6> , \D_Immediate<5> , \D_Immediate<4> ,
         \D_Immediate<3> , \D_Immediate<2> , \D_Immediate<1> ,
         \D_Immediate<0> , D_InvA, D_InvB, D_Cin, PMW_RegFileWrEn,
         D_RegFileWrEn, \PMW_WriteReg<2> , \PMW_WriteReg<1> ,
         \PMW_WriteReg<0> , \D_WriteReg<2> , \D_WriteReg<1> , \D_WriteReg<0> ,
         D_Link, _4_net_, \_5_net_<0> , _6_net_, _7_net_, _8_net_, _9_net_,
         _10_net_, _11_net_, _12_net_, _13_net_, _14_net_, _15_net_, _16_net_,
         _17_net_, _18_net_, \PDE_IncPC<15> , \PDE_IncPC<14> , \PDE_IncPC<13> ,
         \PDE_IncPC<12> , \PDE_IncPC<11> , \PDE_IncPC<10> , \PDE_IncPC<9> ,
         \PDE_IncPC<8> , \PDE_IncPC<7> , \PDE_IncPC<6> , \PDE_IncPC<5> ,
         \PDE_IncPC<4> , \PDE_IncPC<3> , \PDE_IncPC<2> , \PDE_IncPC<1> ,
         \PDE_IncPC<0> , \PDE_ALUOp1<15> , \PDE_ALUOp1<14> , \PDE_ALUOp1<13> ,
         \PDE_ALUOp1<12> , \PDE_ALUOp1<11> , \PDE_ALUOp1<10> , \PDE_ALUOp1<9> ,
         \PDE_ALUOp1<8> , \PDE_ALUOp1<7> , \PDE_ALUOp1<6> , \PDE_ALUOp1<5> ,
         \PDE_ALUOp1<4> , \PDE_ALUOp1<3> , \PDE_ALUOp1<2> , \PDE_ALUOp1<1> ,
         \PDE_ALUOp1<0> , \PDE_ALUOp2<15> , \PDE_ALUOp2<14> , \PDE_ALUOp2<13> ,
         \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , \PDE_ALUOp2<10> , \PDE_ALUOp2<9> ,
         \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , \PDE_ALUOp2<6> , \PDE_ALUOp2<5> ,
         \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , \PDE_ALUOp2<2> , \PDE_ALUOp2<1> ,
         \PDE_ALUOp2<0> , \PDE_Immediate<15> , \PDE_Immediate<14> ,
         \PDE_Immediate<13> , \PDE_Immediate<12> , \PDE_Immediate<11> ,
         \PDE_Immediate<10> , \PDE_Immediate<9> , \PDE_Immediate<8> ,
         \PDE_Immediate<7> , \PDE_Immediate<6> , \PDE_Immediate<5> ,
         \PDE_Immediate<4> , \PDE_Immediate<3> , \PDE_Immediate<2> ,
         \PDE_Immediate<1> , \PDE_Immediate<0> , \PDE_ALUOpcode<2> ,
         \PDE_ALUOpcode<1> , \PDE_ALUOpcode<0> , \PDE_Func<1> , \PDE_Func<0> ,
         PDE_ALUSrc, PDE_Branch, PDE_Jump, PDE_JumpReg, PDE_Set, PDE_Btr,
         PDE_MemWrite, PDE_MemRead, PDE_MemToReg, PDE_Halt, PDE_InvA, PDE_InvB,
         PDE_Cin, _19_net_, \PDE_Rs<2> , \PDE_Rs<1> , \PDE_Rs<0> , \PDE_Rt<2> ,
         \PDE_Rt<1> , \PDE_Rt<0> , \PDE_Rd<2> , \PDE_Rd<1> , \PDE_Rd<0> ,
         _20_net_, \PDE_DecodeIncPC<15> , \PDE_DecodeIncPC<14> ,
         \PDE_DecodeIncPC<13> , \PDE_DecodeIncPC<12> , \PDE_DecodeIncPC<11> ,
         \PDE_DecodeIncPC<10> , \PDE_DecodeIncPC<9> , \PDE_DecodeIncPC<8> ,
         \PDE_DecodeIncPC<7> , \PDE_DecodeIncPC<6> , \PDE_DecodeIncPC<5> ,
         \PDE_DecodeIncPC<4> , \PDE_DecodeIncPC<3> , \PDE_DecodeIncPC<2> ,
         \PDE_DecodeIncPC<1> , \PDE_DecodeIncPC<0> , PDE_Link,
         \E_ExecuteResult<15> , \E_ExecuteResult<14> , \E_ExecuteResult<13> ,
         \E_ExecuteResult<12> , \E_ExecuteResult<11> , \E_ExecuteResult<10> ,
         \E_ExecuteResult<9> , \E_ExecuteResult<8> , \E_ExecuteResult<7> ,
         \E_ExecuteResult<6> , \E_ExecuteResult<5> , \E_ExecuteResult<4> ,
         \E_ExecuteResult<3> , \E_ExecuteResult<2> , \E_ExecuteResult<1> ,
         \E_ExecuteResult<0> , \PEM_Address<15> , \PEM_Address<14> ,
         \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> ,
         \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> ,
         \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> ,
         \PEM_Address<4> , \PEM_Address<3> , \PEM_Address<2> ,
         \PEM_Address<1> , \PEM_Address<0> , \PMW_ExecuteOut<15> ,
         \PMW_ExecuteOut<14> , \PMW_ExecuteOut<13> , \PMW_ExecuteOut<12> ,
         \PMW_ExecuteOut<11> , \PMW_ExecuteOut<10> , \PMW_ExecuteOut<9> ,
         \PMW_ExecuteOut<8> , \PMW_ExecuteOut<7> , \PMW_ExecuteOut<6> ,
         \PMW_ExecuteOut<5> , \PMW_ExecuteOut<4> , \PMW_ExecuteOut<3> ,
         \PMW_ExecuteOut<2> , \PMW_ExecuteOut<1> , \PMW_ExecuteOut<0> ,
         PEM_MemRead, PEM_MemWrite, PEM_MemToReg, \PEM_WriteData<15> ,
         \PEM_WriteData<14> , \PEM_WriteData<13> , \PEM_WriteData<12> ,
         \PEM_WriteData<11> , \PEM_WriteData<10> , \PEM_WriteData<9> ,
         \PEM_WriteData<8> , \PEM_WriteData<7> , \PEM_WriteData<6> ,
         \PEM_WriteData<5> , \PEM_WriteData<4> , \PEM_WriteData<3> ,
         \PEM_WriteData<2> , \PEM_WriteData<1> , \PEM_WriteData<0> ,
         \PEM_Rs<2> , \PEM_Rs<1> , \PEM_Rs<0> , \PEM_Rt<2> , \PEM_Rt<1> ,
         \PEM_Rt<0> , \PEM_Rd<2> , \PEM_Rd<1> , \PEM_Rd<0> , \M_ReadData<15> ,
         \M_ReadData<14> , \M_ReadData<13> , \M_ReadData<12> ,
         \M_ReadData<11> , \M_ReadData<10> , \M_ReadData<9> , \M_ReadData<8> ,
         \M_ReadData<7> , \M_ReadData<6> , \M_ReadData<5> , \M_ReadData<4> ,
         \M_ReadData<3> , \M_ReadData<2> , \M_ReadData<1> , \M_ReadData<0> ,
         _22_net_, \PMW_MemOut<15> , \PMW_MemOut<14> , \PMW_MemOut<13> ,
         \PMW_MemOut<12> , \PMW_MemOut<11> , \PMW_MemOut<10> , \PMW_MemOut<9> ,
         \PMW_MemOut<8> , \PMW_MemOut<7> , \PMW_MemOut<6> , \PMW_MemOut<5> ,
         \PMW_MemOut<4> , \PMW_MemOut<3> , \PMW_MemOut<2> , \PMW_MemOut<1> ,
         \PMW_MemOut<0> , PMW_MemToReg, n8, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;

  AND2X2 U10 ( .A(n67), .B(D_RtValid), .Y(_19_net_) );
  NOR3X1 U27 ( .A(_3_net_), .B(n65), .C(n69), .Y(_15_net_) );
  OAI21X1 U28 ( .A(n63), .B(n8), .C(n62), .Y(_3_net_) );
  AOI22X1 U29 ( .A(PDE_RegFileWrEn), .B(n43), .C(PEM_RegFileWrEn), .D(n44), 
        .Y(n8) );
  NAND3X1 U30 ( .A(n52), .B(n54), .C(n46), .Y(n11) );
  NAND3X1 U31 ( .A(n15), .B(n16), .C(n50), .Y(n14) );
  XOR2X1 U33 ( .A(\PEM_WriteReg<2> ), .B(\D_Rs<2> ), .Y(n18) );
  XNOR2X1 U34 ( .A(\D_Rs<1> ), .B(\PEM_WriteReg<1> ), .Y(n16) );
  XNOR2X1 U35 ( .A(\D_Rs<0> ), .B(\PEM_WriteReg<0> ), .Y(n15) );
  NAND3X1 U36 ( .A(n19), .B(n20), .C(n21), .Y(n13) );
  NOR3X1 U37 ( .A(n22), .B(n70), .C(n72), .Y(n21) );
  XOR2X1 U38 ( .A(\PEM_WriteReg<2> ), .B(\D_Rd<2> ), .Y(n22) );
  XNOR2X1 U39 ( .A(\D_Rd<1> ), .B(\PEM_WriteReg<1> ), .Y(n20) );
  XNOR2X1 U40 ( .A(\D_Rd<0> ), .B(\PEM_WriteReg<0> ), .Y(n19) );
  NAND3X1 U41 ( .A(n23), .B(n24), .C(n60), .Y(n12) );
  XOR2X1 U43 ( .A(\PEM_WriteReg<2> ), .B(\D_Rt<2> ), .Y(n26) );
  XNOR2X1 U44 ( .A(\D_Rt<1> ), .B(\PEM_WriteReg<1> ), .Y(n24) );
  XNOR2X1 U45 ( .A(\D_Rt<0> ), .B(\PEM_WriteReg<0> ), .Y(n23) );
  NAND3X1 U46 ( .A(n42), .B(n51), .C(n45), .Y(n10) );
  NAND3X1 U47 ( .A(n30), .B(n56), .C(n31), .Y(n29) );
  XOR2X1 U49 ( .A(\PDE_WriteReg<2> ), .B(\D_Rs<2> ), .Y(n33) );
  XNOR2X1 U50 ( .A(\D_Rs<1> ), .B(\PDE_WriteReg<1> ), .Y(n31) );
  XNOR2X1 U51 ( .A(\D_Rs<0> ), .B(\PDE_WriteReg<0> ), .Y(n30) );
  NAND3X1 U52 ( .A(n34), .B(n35), .C(n36), .Y(n28) );
  NOR3X1 U53 ( .A(n37), .B(n70), .C(n72), .Y(n36) );
  XOR2X1 U54 ( .A(\PDE_WriteReg<2> ), .B(\D_Rd<2> ), .Y(n37) );
  XNOR2X1 U55 ( .A(\D_Rd<1> ), .B(\PDE_WriteReg<1> ), .Y(n35) );
  XNOR2X1 U56 ( .A(\D_Rd<0> ), .B(\PDE_WriteReg<0> ), .Y(n34) );
  NAND3X1 U57 ( .A(n38), .B(n39), .C(n58), .Y(n27) );
  XOR2X1 U59 ( .A(\PDE_WriteReg<2> ), .B(\D_Rt<2> ), .Y(n41) );
  XNOR2X1 U60 ( .A(\D_Rt<1> ), .B(\PDE_WriteReg<1> ), .Y(n39) );
  XNOR2X1 U61 ( .A(\D_Rt<0> ), .B(\PDE_WriteReg<0> ), .Y(n38) );
  fetch f ( .BranchPC({\E_BranchPC<15> , \E_BranchPC<14> , \E_BranchPC<13> , 
        \E_BranchPC<12> , \E_BranchPC<11> , \E_BranchPC<10> , \E_BranchPC<9> , 
        \E_BranchPC<8> , \E_BranchPC<7> , \E_BranchPC<6> , \E_BranchPC<5> , 
        \E_BranchPC<4> , \E_BranchPC<3> , \E_BranchPC<2> , \E_BranchPC<1> , 
        \E_BranchPC<0> }), .BranchJumpTaken(n48), .clk(clk), .rst(n65), .Halt(
        PEM_Halt), .Rti(D_Rti), .Exception(D_Exception), .Stall(_3_net_), 
        .Instr({\F_Instr<15> , \F_Instr<14> , \F_Instr<13> , \F_Instr<12> , 
        \F_Instr<11> , \F_Instr<10> , \F_Instr<9> , \F_Instr<8> , \F_Instr<7> , 
        \F_Instr<6> , \F_Instr<5> , \F_Instr<4> , \F_Instr<3> , \F_Instr<2> , 
        \F_Instr<1> , \F_Instr<0> }), .IncPC({\F_IncPC<15> , \F_IncPC<14> , 
        \F_IncPC<13> , \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , 
        \F_IncPC<9> , \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , 
        \F_IncPC<4> , \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> }), 
        .Err(), .CacheHit(), .InstrMemStall() );
  pipe_fd fd ( .Stall(_3_net_), .Flush(n63), .rst(n63), .clk(clk), .Instr({
        \F_Instr<15> , \F_Instr<14> , \F_Instr<13> , \F_Instr<12> , 
        \F_Instr<11> , \F_Instr<10> , \F_Instr<9> , \F_Instr<8> , \F_Instr<7> , 
        \F_Instr<6> , \F_Instr<5> , \F_Instr<4> , \F_Instr<3> , \F_Instr<2> , 
        \F_Instr<1> , \F_Instr<0> }), .IncPC({\F_IncPC<15> , \F_IncPC<14> , 
        \F_IncPC<13> , \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , 
        \F_IncPC<9> , \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , 
        \F_IncPC<4> , \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> }), 
        .Instr_Out({\PFD_Instr<15> , \PFD_Instr<14> , \PFD_Instr<13> , 
        \PFD_Instr<12> , \PFD_Instr<11> , \PFD_Instr<10> , \PFD_Instr<9> , 
        \PFD_Instr<8> , \PFD_Instr<7> , \PFD_Instr<6> , \PFD_Instr<5> , 
        \PFD_Instr<4> , \PFD_Instr<3> , \PFD_Instr<2> , \PFD_Instr<1> , 
        \PFD_Instr<0> }), .IncPC_Out({\PFD_IncPC<15> , \PFD_IncPC<14> , 
        \PFD_IncPC<13> , \PFD_IncPC<12> , \PFD_IncPC<11> , \PFD_IncPC<10> , 
        \PFD_IncPC<9> , \PFD_IncPC<8> , \PFD_IncPC<7> , \PFD_IncPC<6> , 
        \PFD_IncPC<5> , \PFD_IncPC<4> , \PFD_IncPC<3> , \PFD_IncPC<2> , 
        \PFD_IncPC<1> , \PFD_IncPC<0> }), .CPUActive(PFD_CPUActive) );
  decode d ( .clk(clk), .rst(n65), .Stall(_3_net_), .Instr({\PFD_Instr<15> , 
        \PFD_Instr<14> , \PFD_Instr<13> , \PFD_Instr<12> , \PFD_Instr<11> , 
        \PFD_Instr<10> , \PFD_Instr<9> , \PFD_Instr<8> , \PFD_Instr<7> , 
        \PFD_Instr<6> , \PFD_Instr<5> , \PFD_Instr<4> , \PFD_Instr<3> , 
        \PFD_Instr<2> , \PFD_Instr<1> , \PFD_Instr<0> }), .WriteData({
        \W_WriteData<15> , \W_WriteData<14> , \W_WriteData<13> , 
        \W_WriteData<12> , \W_WriteData<11> , \W_WriteData<10> , 
        \W_WriteData<9> , \W_WriteData<8> , \W_WriteData<7> , \W_WriteData<6> , 
        \W_WriteData<5> , \W_WriteData<4> , \W_WriteData<3> , \W_WriteData<2> , 
        \W_WriteData<1> , \W_WriteData<0> }), .IncPC({\PFD_IncPC<15> , 
        \PFD_IncPC<14> , \PFD_IncPC<13> , \PFD_IncPC<12> , \PFD_IncPC<11> , 
        \PFD_IncPC<10> , \PFD_IncPC<9> , \PFD_IncPC<8> , \PFD_IncPC<7> , 
        \PFD_IncPC<6> , \PFD_IncPC<5> , \PFD_IncPC<4> , \PFD_IncPC<3> , 
        \PFD_IncPC<2> , \PFD_IncPC<1> , \PFD_IncPC<0> }), .ALUOp1({
        \D_ALUOp1<15> , \D_ALUOp1<14> , \D_ALUOp1<13> , \D_ALUOp1<12> , 
        \D_ALUOp1<11> , \D_ALUOp1<10> , \D_ALUOp1<9> , \D_ALUOp1<8> , 
        \D_ALUOp1<7> , \D_ALUOp1<6> , \D_ALUOp1<5> , \D_ALUOp1<4> , 
        \D_ALUOp1<3> , \D_ALUOp1<2> , \D_ALUOp1<1> , \D_ALUOp1<0> }), .ALUOp2(
        {\D_ALUOp2<15> , \D_ALUOp2<14> , \D_ALUOp2<13> , \D_ALUOp2<12> , 
        \D_ALUOp2<11> , \D_ALUOp2<10> , \D_ALUOp2<9> , \D_ALUOp2<8> , 
        \D_ALUOp2<7> , \D_ALUOp2<6> , \D_ALUOp2<5> , \D_ALUOp2<4> , 
        \D_ALUOp2<3> , \D_ALUOp2<2> , \D_ALUOp2<1> , \D_ALUOp2<0> }), .ALUSrc(
        D_ALUSrc), .Immediate({\D_Immediate<15> , \D_Immediate<14> , 
        \D_Immediate<13> , \D_Immediate<12> , \D_Immediate<11> , 
        \D_Immediate<10> , \D_Immediate<9> , \D_Immediate<8> , 
        \D_Immediate<7> , \D_Immediate<6> , \D_Immediate<5> , \D_Immediate<4> , 
        \D_Immediate<3> , \D_Immediate<2> , \D_Immediate<1> , \D_Immediate<0> }), .Branch(D_Branch), .Jump(D_Jump), .JumpReg(D_JumpReg), .Set(D_Set), .Btr(
        D_Btr), .InvA(D_InvA), .InvB(D_InvB), .Cin(D_Cin), .ALUOpcode({
        \D_ALUOpcode<2> , \D_ALUOpcode<1> , \D_ALUOpcode<0> }), .Func({
        \D_Func<1> , \D_Func<0> }), .MemWrite(D_MemWrite), .MemRead(D_MemRead), 
        .MemToReg(D_MemToReg), .Halt(D_Halt), .Exception(D_Exception), .Err(), 
        .Rti(D_Rti), .Rs({\D_Rs<2> , \D_Rs<1> , \D_Rs<0> }), .Rt({\D_Rt<2> , 
        \D_Rt<1> , \D_Rt<0> }), .Rd({\D_Rd<2> , \D_Rd<1> , \D_Rd<0> }), 
        .RegFileWrEn(PMW_RegFileWrEn), .RegFileWrEn_Out(D_RegFileWrEn), 
        .WriteReg({\PMW_WriteReg<2> , \PMW_WriteReg<1> , \PMW_WriteReg<0> }), 
        .WriteReg_Out({\D_WriteReg<2> , \D_WriteReg<1> , \D_WriteReg<0> }), 
        .RtValid(D_RtValid), .RsValid(D_RsValid), .RdValid(D_RdValid), .Link(
        D_Link), .Store(D_Store) );
  pipe_de pde ( .clk(clk), .rst(n63), .Stall(n61), .Flush(n63), .ALUOp1({
        \D_ALUOp1<15> , \D_ALUOp1<14> , \D_ALUOp1<13> , \D_ALUOp1<12> , 
        \D_ALUOp1<11> , \D_ALUOp1<10> , \D_ALUOp1<9> , \D_ALUOp1<8> , 
        \D_ALUOp1<7> , \D_ALUOp1<6> , \D_ALUOp1<5> , \D_ALUOp1<4> , 
        \D_ALUOp1<3> , \D_ALUOp1<2> , \D_ALUOp1<1> , \D_ALUOp1<0> }), .ALUOp2(
        {\D_ALUOp2<15> , \D_ALUOp2<14> , \D_ALUOp2<13> , \D_ALUOp2<12> , 
        \D_ALUOp2<11> , \D_ALUOp2<10> , \D_ALUOp2<9> , \D_ALUOp2<8> , 
        \D_ALUOp2<7> , \D_ALUOp2<6> , \D_ALUOp2<5> , \D_ALUOp2<4> , 
        \D_ALUOp2<3> , \D_ALUOp2<2> , \D_ALUOp2<1> , \D_ALUOp2<0> }), 
        .Immediate({\D_Immediate<15> , \D_Immediate<14> , \D_Immediate<13> , 
        \D_Immediate<12> , \D_Immediate<11> , \D_Immediate<10> , 
        \D_Immediate<9> , \D_Immediate<8> , \D_Immediate<7> , \D_Immediate<6> , 
        \D_Immediate<5> , \D_Immediate<4> , \D_Immediate<3> , \D_Immediate<2> , 
        \D_Immediate<1> , \D_Immediate<0> }), .ALUOpcode({\D_ALUOpcode<2> , 
        \D_ALUOpcode<1> , \D_ALUOpcode<0> }), .Func({\D_Func<1> , \_5_net_<0> }), .ALUSrc(_6_net_), .Branch(_7_net_), .Jump(_8_net_), .JumpReg(_9_net_), 
        .Set(_10_net_), .Btr(_11_net_), .MemWrite(_12_net_), .MemRead(_13_net_), .MemToReg(_14_net_), .Halt(_15_net_), .InvA(_16_net_), .InvB(_17_net_), 
        .Cin(_18_net_), .IncPC({\F_IncPC<15> , \F_IncPC<14> , \F_IncPC<13> , 
        \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , \F_IncPC<9> , 
        \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , \F_IncPC<4> , 
        \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> }), .CPUActive(
        PFD_CPUActive), .ALUOp1_Out({\PDE_ALUOp1<15> , \PDE_ALUOp1<14> , 
        \PDE_ALUOp1<13> , \PDE_ALUOp1<12> , \PDE_ALUOp1<11> , \PDE_ALUOp1<10> , 
        \PDE_ALUOp1<9> , \PDE_ALUOp1<8> , \PDE_ALUOp1<7> , \PDE_ALUOp1<6> , 
        \PDE_ALUOp1<5> , \PDE_ALUOp1<4> , \PDE_ALUOp1<3> , \PDE_ALUOp1<2> , 
        \PDE_ALUOp1<1> , \PDE_ALUOp1<0> }), .ALUOp2_Out({\PDE_ALUOp2<15> , 
        \PDE_ALUOp2<14> , \PDE_ALUOp2<13> , \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , 
        \PDE_ALUOp2<10> , \PDE_ALUOp2<9> , \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , 
        \PDE_ALUOp2<6> , \PDE_ALUOp2<5> , \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , 
        \PDE_ALUOp2<2> , \PDE_ALUOp2<1> , \PDE_ALUOp2<0> }), .Immediate_Out({
        \PDE_Immediate<15> , \PDE_Immediate<14> , \PDE_Immediate<13> , 
        \PDE_Immediate<12> , \PDE_Immediate<11> , \PDE_Immediate<10> , 
        \PDE_Immediate<9> , \PDE_Immediate<8> , \PDE_Immediate<7> , 
        \PDE_Immediate<6> , \PDE_Immediate<5> , \PDE_Immediate<4> , 
        \PDE_Immediate<3> , \PDE_Immediate<2> , \PDE_Immediate<1> , 
        \PDE_Immediate<0> }), .ALUOpcode_Out({\PDE_ALUOpcode<2> , 
        \PDE_ALUOpcode<1> , \PDE_ALUOpcode<0> }), .Func_Out({\PDE_Func<1> , 
        \PDE_Func<0> }), .ALUSrc_Out(PDE_ALUSrc), .Branch_Out(PDE_Branch), 
        .Jump_Out(PDE_Jump), .JumpReg_Out(PDE_JumpReg), .Set_Out(PDE_Set), 
        .Btr_Out(PDE_Btr), .MemWrite_Out(PDE_MemWrite), .MemRead_Out(
        PDE_MemRead), .MemToReg_Out(PDE_MemToReg), .Halt_Out(PDE_Halt), 
        .InvA_Out(PDE_InvA), .InvB_Out(PDE_InvB), .Cin_Out(PDE_Cin), .Rs({
        \D_Rs<2> , \D_Rs<1> , \D_Rs<0> }), .Rt({\D_Rt<2> , \D_Rt<1> , 
        \D_Rt<0> }), .Rd({\D_Rd<2> , \D_Rd<1> , \D_Rd<0> }), .Rs_Out({
        \PDE_Rs<2> , \PDE_Rs<1> , \PDE_Rs<0> }), .Rt_Out({\PDE_Rt<2> , 
        \PDE_Rt<1> , \PDE_Rt<0> }), .Rd_Out({\PDE_Rd<2> , \PDE_Rd<1> , 
        \PDE_Rd<0> }), .RegFileWrEn(_20_net_), .RegFileWrEn_Out(
        PDE_RegFileWrEn), .IncPC_Out({\PDE_IncPC<15> , \PDE_IncPC<14> , 
        \PDE_IncPC<13> , \PDE_IncPC<12> , \PDE_IncPC<11> , \PDE_IncPC<10> , 
        \PDE_IncPC<9> , \PDE_IncPC<8> , \PDE_IncPC<7> , \PDE_IncPC<6> , 
        \PDE_IncPC<5> , \PDE_IncPC<4> , \PDE_IncPC<3> , \PDE_IncPC<2> , 
        \PDE_IncPC<1> , \PDE_IncPC<0> }), .WriteReg({\D_WriteReg<2> , 
        \D_WriteReg<1> , \D_WriteReg<0> }), .WriteReg_Out({\PDE_WriteReg<2> , 
        \PDE_WriteReg<1> , \PDE_WriteReg<0> }), .RtValid(_19_net_), 
        .RtValid_Out(), .CPUActive_Out(), .RsValid(D_RsValid), .RdValid(
        D_RdValid), .RsValid_Out(), .RdValid_Out(), .DecodeIncPC({
        \PFD_IncPC<15> , \PFD_IncPC<14> , \PFD_IncPC<13> , \PFD_IncPC<12> , 
        \PFD_IncPC<11> , \PFD_IncPC<10> , \PFD_IncPC<9> , \PFD_IncPC<8> , 
        \PFD_IncPC<7> , \PFD_IncPC<6> , \PFD_IncPC<5> , \PFD_IncPC<4> , 
        \PFD_IncPC<3> , \PFD_IncPC<2> , \PFD_IncPC<1> , \PFD_IncPC<0> }), 
        .DecodeIncPC_Out({\PDE_DecodeIncPC<15> , \PDE_DecodeIncPC<14> , 
        \PDE_DecodeIncPC<13> , \PDE_DecodeIncPC<12> , \PDE_DecodeIncPC<11> , 
        \PDE_DecodeIncPC<10> , \PDE_DecodeIncPC<9> , \PDE_DecodeIncPC<8> , 
        \PDE_DecodeIncPC<7> , \PDE_DecodeIncPC<6> , \PDE_DecodeIncPC<5> , 
        \PDE_DecodeIncPC<4> , \PDE_DecodeIncPC<3> , \PDE_DecodeIncPC<2> , 
        \PDE_DecodeIncPC<1> , \PDE_DecodeIncPC<0> }), .Link(D_Link), 
        .Link_Out(PDE_Link) );
  execute e ( .ALUOp1({\PDE_ALUOp1<15> , \PDE_ALUOp1<14> , \PDE_ALUOp1<13> , 
        \PDE_ALUOp1<12> , \PDE_ALUOp1<11> , \PDE_ALUOp1<10> , \PDE_ALUOp1<9> , 
        \PDE_ALUOp1<8> , \PDE_ALUOp1<7> , \PDE_ALUOp1<6> , \PDE_ALUOp1<5> , 
        \PDE_ALUOp1<4> , \PDE_ALUOp1<3> , \PDE_ALUOp1<2> , \PDE_ALUOp1<1> , 
        \PDE_ALUOp1<0> }), .ALUOp2({\PDE_ALUOp2<15> , \PDE_ALUOp2<14> , 
        \PDE_ALUOp2<13> , \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , \PDE_ALUOp2<10> , 
        \PDE_ALUOp2<9> , \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , \PDE_ALUOp2<6> , 
        \PDE_ALUOp2<5> , \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , \PDE_ALUOp2<2> , 
        \PDE_ALUOp2<1> , \PDE_ALUOp2<0> }), .Opcode({\PDE_ALUOpcode<2> , 
        \PDE_ALUOpcode<1> , \PDE_ALUOpcode<0> }), .IncPC({\PDE_IncPC<15> , 
        \PDE_IncPC<14> , \PDE_IncPC<13> , \PDE_IncPC<12> , \PDE_IncPC<11> , 
        \PDE_IncPC<10> , \PDE_IncPC<9> , \PDE_IncPC<8> , \PDE_IncPC<7> , 
        \PDE_IncPC<6> , \PDE_IncPC<5> , \PDE_IncPC<4> , \PDE_IncPC<3> , 
        \PDE_IncPC<2> , \PDE_IncPC<1> , \PDE_IncPC<0> }), .Jump(PDE_Jump), 
        .Branch(PDE_Branch), .JumpReg(PDE_JumpReg), .Set(PDE_Set), .InvA(
        PDE_InvA), .InvB(PDE_InvB), .Cin(PDE_Cin), .Btr(PDE_Btr), .Func({
        \PDE_Func<1> , \PDE_Func<0> }), .Imm({\PDE_Immediate<15> , 
        \PDE_Immediate<14> , \PDE_Immediate<13> , \PDE_Immediate<12> , 
        \PDE_Immediate<11> , \PDE_Immediate<10> , \PDE_Immediate<9> , 
        \PDE_Immediate<8> , \PDE_Immediate<7> , \PDE_Immediate<6> , 
        \PDE_Immediate<5> , \PDE_Immediate<4> , \PDE_Immediate<3> , 
        \PDE_Immediate<2> , \PDE_Immediate<1> , \PDE_Immediate<0> }), .ALUSrc(
        PDE_ALUSrc), .Result({\E_ExecuteResult<15> , \E_ExecuteResult<14> , 
        \E_ExecuteResult<13> , \E_ExecuteResult<12> , \E_ExecuteResult<11> , 
        \E_ExecuteResult<10> , \E_ExecuteResult<9> , \E_ExecuteResult<8> , 
        \E_ExecuteResult<7> , \E_ExecuteResult<6> , \E_ExecuteResult<5> , 
        \E_ExecuteResult<4> , \E_ExecuteResult<3> , \E_ExecuteResult<2> , 
        \E_ExecuteResult<1> , \E_ExecuteResult<0> }), .NextPC({
        \E_BranchPC<15> , \E_BranchPC<14> , \E_BranchPC<13> , \E_BranchPC<12> , 
        \E_BranchPC<11> , \E_BranchPC<10> , \E_BranchPC<9> , \E_BranchPC<8> , 
        \E_BranchPC<7> , \E_BranchPC<6> , \E_BranchPC<5> , \E_BranchPC<4> , 
        \E_BranchPC<3> , \E_BranchPC<2> , \E_BranchPC<1> , \E_BranchPC<0> }), 
        .Err(), .BranchJumpTaken(E_BranchJumpTaken), .rst(n65), .DecodeIncPC({
        \PDE_DecodeIncPC<15> , \PDE_DecodeIncPC<14> , \PDE_DecodeIncPC<13> , 
        \PDE_DecodeIncPC<12> , \PDE_DecodeIncPC<11> , \PDE_DecodeIncPC<10> , 
        \PDE_DecodeIncPC<9> , \PDE_DecodeIncPC<8> , \PDE_DecodeIncPC<7> , 
        \PDE_DecodeIncPC<6> , \PDE_DecodeIncPC<5> , \PDE_DecodeIncPC<4> , 
        \PDE_DecodeIncPC<3> , \PDE_DecodeIncPC<2> , \PDE_DecodeIncPC<1> , 
        \PDE_DecodeIncPC<0> }), .Link(PDE_Link), .ForwardALUOp1({1'b0, 1'b0}), 
        .ForwardALUOp2({1'b0, 1'b0}), .PipeMW_Result({\PMW_ExecuteOut<15> , 
        \PMW_ExecuteOut<14> , \PMW_ExecuteOut<13> , \PMW_ExecuteOut<12> , 
        \PMW_ExecuteOut<11> , \PMW_ExecuteOut<10> , \PMW_ExecuteOut<9> , 
        \PMW_ExecuteOut<8> , \PMW_ExecuteOut<7> , \PMW_ExecuteOut<6> , 
        \PMW_ExecuteOut<5> , \PMW_ExecuteOut<4> , \PMW_ExecuteOut<3> , 
        \PMW_ExecuteOut<2> , \PMW_ExecuteOut<1> , \PMW_ExecuteOut<0> }), 
        .PipeEM_Result({\PEM_Address<15> , \PEM_Address<14> , 
        \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> , 
        \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> , 
        \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> , \PEM_Address<4> , 
        \PEM_Address<3> , \PEM_Address<2> , \PEM_Address<1> , \PEM_Address<0> }) );
  pipe_em pem ( .Stall(M_DataMemStall), .rst(n65), .clk(clk), .Result({
        \E_ExecuteResult<15> , \E_ExecuteResult<14> , \E_ExecuteResult<13> , 
        \E_ExecuteResult<12> , \E_ExecuteResult<11> , \E_ExecuteResult<10> , 
        \E_ExecuteResult<9> , \E_ExecuteResult<8> , \E_ExecuteResult<7> , 
        \E_ExecuteResult<6> , \E_ExecuteResult<5> , \E_ExecuteResult<4> , 
        \E_ExecuteResult<3> , \E_ExecuteResult<2> , \E_ExecuteResult<1> , 
        \E_ExecuteResult<0> }), .MemRead(PDE_MemRead), .MemWrite(PDE_MemWrite), 
        .MemToReg(PDE_MemToReg), .Halt(PDE_Halt), .ALUOp2({\PDE_ALUOp2<15> , 
        \PDE_ALUOp2<14> , \PDE_ALUOp2<13> , \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , 
        \PDE_ALUOp2<10> , \PDE_ALUOp2<9> , \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , 
        \PDE_ALUOp2<6> , \PDE_ALUOp2<5> , \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , 
        \PDE_ALUOp2<2> , \PDE_ALUOp2<1> , \PDE_ALUOp2<0> }), .RegFileWrEn(
        PDE_RegFileWrEn), .Rs({\PDE_Rs<2> , \PDE_Rs<1> , \PDE_Rs<0> }), .Rt({
        \PDE_Rt<2> , \PDE_Rt<1> , \PDE_Rt<0> }), .Rd({\PDE_Rd<2> , \PDE_Rd<1> , 
        \PDE_Rd<0> }), .WriteReg({\PDE_WriteReg<2> , \PDE_WriteReg<1> , 
        \PDE_WriteReg<0> }), .Address({\PEM_Address<15> , \PEM_Address<14> , 
        \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> , 
        \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> , 
        \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> , \PEM_Address<4> , 
        \PEM_Address<3> , \PEM_Address<2> , \PEM_Address<1> , \PEM_Address<0> }), .MemRead_Out(PEM_MemRead), .MemWrite_Out(PEM_MemWrite), .MemToReg_Out(
        PEM_MemToReg), .Halt_Out(PEM_Halt), .WriteData({\PEM_WriteData<15> , 
        \PEM_WriteData<14> , \PEM_WriteData<13> , \PEM_WriteData<12> , 
        \PEM_WriteData<11> , \PEM_WriteData<10> , \PEM_WriteData<9> , 
        \PEM_WriteData<8> , \PEM_WriteData<7> , \PEM_WriteData<6> , 
        \PEM_WriteData<5> , \PEM_WriteData<4> , \PEM_WriteData<3> , 
        \PEM_WriteData<2> , \PEM_WriteData<1> , \PEM_WriteData<0> }), 
        .RegFileWrEn_Out(PEM_RegFileWrEn), .Rs_Out({\PEM_Rs<2> , \PEM_Rs<1> , 
        \PEM_Rs<0> }), .Rt_Out({\PEM_Rt<2> , \PEM_Rt<1> , \PEM_Rt<0> }), 
        .Rd_Out({\PEM_Rd<2> , \PEM_Rd<1> , \PEM_Rd<0> }), .WriteReg_Out({
        \PEM_WriteReg<2> , \PEM_WriteReg<1> , \PEM_WriteReg<0> }) );
  memory m ( .MemRead(PEM_MemRead), .MemWrite(PEM_MemWrite), .halt(PEM_Halt), 
        .clk(clk), .rst(n65), .Address({\PEM_Address<15> , \PEM_Address<14> , 
        \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> , 
        \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> , 
        \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> , \PEM_Address<4> , 
        \PEM_Address<3> , \PEM_Address<2> , \PEM_Address<1> , \PEM_Address<0> }), .WriteData({\PEM_WriteData<15> , \PEM_WriteData<14> , \PEM_WriteData<13> , 
        \PEM_WriteData<12> , \PEM_WriteData<11> , \PEM_WriteData<10> , 
        \PEM_WriteData<9> , \PEM_WriteData<8> , \PEM_WriteData<7> , 
        \PEM_WriteData<6> , \PEM_WriteData<5> , \PEM_WriteData<4> , 
        \PEM_WriteData<3> , \PEM_WriteData<2> , \PEM_WriteData<1> , 
        \PEM_WriteData<0> }), .ReadData({\M_ReadData<15> , \M_ReadData<14> , 
        \M_ReadData<13> , \M_ReadData<12> , \M_ReadData<11> , \M_ReadData<10> , 
        \M_ReadData<9> , \M_ReadData<8> , \M_ReadData<7> , \M_ReadData<6> , 
        \M_ReadData<5> , \M_ReadData<4> , \M_ReadData<3> , \M_ReadData<2> , 
        \M_ReadData<1> , \M_ReadData<0> }), .Err(M_Err), .DataMemStall(
        M_DataMemStall), .CacheHit() );
  pipe_mw pmw ( .Stall(1'b0), .rst(_22_net_), .clk(clk), .ExecuteOut({
        \PEM_Address<15> , \PEM_Address<14> , \PEM_Address<13> , 
        \PEM_Address<12> , \PEM_Address<11> , \PEM_Address<10> , 
        \PEM_Address<9> , \PEM_Address<8> , \PEM_Address<7> , \PEM_Address<6> , 
        \PEM_Address<5> , \PEM_Address<4> , \PEM_Address<3> , \PEM_Address<2> , 
        \PEM_Address<1> , \PEM_Address<0> }), .MemOut({\M_ReadData<15> , 
        \M_ReadData<14> , \M_ReadData<13> , \M_ReadData<12> , \M_ReadData<11> , 
        \M_ReadData<10> , \M_ReadData<9> , \M_ReadData<8> , \M_ReadData<7> , 
        \M_ReadData<6> , \M_ReadData<5> , \M_ReadData<4> , \M_ReadData<3> , 
        \M_ReadData<2> , \M_ReadData<1> , \M_ReadData<0> }), .MemToReg(
        PEM_MemToReg), .RegFileWrEn(PEM_RegFileWrEn), .Rs({\PEM_Rs<2> , 
        \PEM_Rs<1> , \PEM_Rs<0> }), .Rt({\PEM_Rt<2> , \PEM_Rt<1> , \PEM_Rt<0> }), .Rd({\PEM_Rd<2> , \PEM_Rd<1> , \PEM_Rd<0> }), .WriteReg({\PEM_WriteReg<2> , 
        \PEM_WriteReg<1> , \PEM_WriteReg<0> }), .ExecuteOut_Out({
        \PMW_ExecuteOut<15> , \PMW_ExecuteOut<14> , \PMW_ExecuteOut<13> , 
        \PMW_ExecuteOut<12> , \PMW_ExecuteOut<11> , \PMW_ExecuteOut<10> , 
        \PMW_ExecuteOut<9> , \PMW_ExecuteOut<8> , \PMW_ExecuteOut<7> , 
        \PMW_ExecuteOut<6> , \PMW_ExecuteOut<5> , \PMW_ExecuteOut<4> , 
        \PMW_ExecuteOut<3> , \PMW_ExecuteOut<2> , \PMW_ExecuteOut<1> , 
        \PMW_ExecuteOut<0> }), .MemOut_Out({\PMW_MemOut<15> , \PMW_MemOut<14> , 
        \PMW_MemOut<13> , \PMW_MemOut<12> , \PMW_MemOut<11> , \PMW_MemOut<10> , 
        \PMW_MemOut<9> , \PMW_MemOut<8> , \PMW_MemOut<7> , \PMW_MemOut<6> , 
        \PMW_MemOut<5> , \PMW_MemOut<4> , \PMW_MemOut<3> , \PMW_MemOut<2> , 
        \PMW_MemOut<1> , \PMW_MemOut<0> }), .MemToReg_Out(PMW_MemToReg), 
        .RegFileWrEn_Out(PMW_RegFileWrEn), .WriteReg_Out({\PMW_WriteReg<2> , 
        \PMW_WriteReg<1> , \PMW_WriteReg<0> }), .Rs_Out(), .Rt_Out(), 
        .Rd_Out() );
  writeback w ( .ExecuteOut({\PMW_ExecuteOut<15> , \PMW_ExecuteOut<14> , 
        \PMW_ExecuteOut<13> , \PMW_ExecuteOut<12> , \PMW_ExecuteOut<11> , 
        \PMW_ExecuteOut<10> , \PMW_ExecuteOut<9> , \PMW_ExecuteOut<8> , 
        \PMW_ExecuteOut<7> , \PMW_ExecuteOut<6> , \PMW_ExecuteOut<5> , 
        \PMW_ExecuteOut<4> , \PMW_ExecuteOut<3> , \PMW_ExecuteOut<2> , 
        \PMW_ExecuteOut<1> , \PMW_ExecuteOut<0> }), .MemOut({\PMW_MemOut<15> , 
        \PMW_MemOut<14> , \PMW_MemOut<13> , \PMW_MemOut<12> , \PMW_MemOut<11> , 
        \PMW_MemOut<10> , \PMW_MemOut<9> , \PMW_MemOut<8> , \PMW_MemOut<7> , 
        \PMW_MemOut<6> , \PMW_MemOut<5> , \PMW_MemOut<4> , \PMW_MemOut<3> , 
        \PMW_MemOut<2> , \PMW_MemOut<1> , \PMW_MemOut<0> }), .MemToReg(
        PMW_MemToReg), .WriteData({\W_WriteData<15> , \W_WriteData<14> , 
        \W_WriteData<13> , \W_WriteData<12> , \W_WriteData<11> , 
        \W_WriteData<10> , \W_WriteData<9> , \W_WriteData<8> , 
        \W_WriteData<7> , \W_WriteData<6> , \W_WriteData<5> , \W_WriteData<4> , 
        \W_WriteData<3> , \W_WriteData<2> , \W_WriteData<1> , \W_WriteData<0> }) );
  INVX1 U63 ( .A(n64), .Y(n63) );
  INVX1 U64 ( .A(_4_net_), .Y(n64) );
  OR2X1 U65 ( .A(n48), .B(n65), .Y(_4_net_) );
  INVX1 U66 ( .A(_3_net_), .Y(n67) );
  INVX1 U67 ( .A(rst), .Y(n66) );
  AND2X1 U68 ( .A(D_RegFileWrEn), .B(n67), .Y(_20_net_) );
  AND2X1 U69 ( .A(\D_Func<0> ), .B(n67), .Y(\_5_net_<0> ) );
  AND2X1 U70 ( .A(D_ALUSrc), .B(n67), .Y(_6_net_) );
  AND2X1 U71 ( .A(D_Branch), .B(n67), .Y(_7_net_) );
  AND2X1 U72 ( .A(D_Jump), .B(n67), .Y(_8_net_) );
  AND2X1 U73 ( .A(D_JumpReg), .B(n67), .Y(_9_net_) );
  AND2X1 U74 ( .A(D_Set), .B(n67), .Y(_10_net_) );
  AND2X1 U75 ( .A(D_Btr), .B(n67), .Y(_11_net_) );
  AND2X1 U76 ( .A(D_MemToReg), .B(n67), .Y(_14_net_) );
  AND2X1 U77 ( .A(D_InvA), .B(n67), .Y(_16_net_) );
  AND2X1 U78 ( .A(D_InvB), .B(n67), .Y(_17_net_) );
  AND2X1 U79 ( .A(D_Cin), .B(n67), .Y(_18_net_) );
  INVX1 U80 ( .A(D_RtValid), .Y(n71) );
  INVX1 U81 ( .A(D_Store), .Y(n72) );
  AND2X1 U82 ( .A(D_MemWrite), .B(n67), .Y(_12_net_) );
  AND2X1 U83 ( .A(D_MemRead), .B(n67), .Y(_13_net_) );
  INVX1 U84 ( .A(D_Halt), .Y(n69) );
  OR2X1 U85 ( .A(1'b0), .B(M_Err), .Y(err) );
  OR2X1 U86 ( .A(n65), .B(M_DataMemStall), .Y(_22_net_) );
  INVX1 U87 ( .A(n66), .Y(n65) );
  BUFX2 U88 ( .A(n28), .Y(n42) );
  BUFX2 U89 ( .A(n10), .Y(n43) );
  BUFX2 U90 ( .A(n11), .Y(n44) );
  BUFX2 U91 ( .A(n29), .Y(n45) );
  BUFX2 U92 ( .A(n14), .Y(n46) );
  INVX1 U93 ( .A(E_BranchJumpTaken), .Y(n47) );
  INVX1 U94 ( .A(n47), .Y(n48) );
  OR2X1 U95 ( .A(n68), .B(n18), .Y(n49) );
  INVX1 U96 ( .A(n49), .Y(n50) );
  BUFX2 U97 ( .A(n27), .Y(n51) );
  BUFX2 U98 ( .A(n12), .Y(n52) );
  INVX1 U99 ( .A(n13), .Y(n53) );
  INVX1 U100 ( .A(n53), .Y(n54) );
  OR2X2 U101 ( .A(n68), .B(n33), .Y(n55) );
  INVX1 U102 ( .A(n55), .Y(n56) );
  INVX1 U103 ( .A(D_RsValid), .Y(n68) );
  OR2X1 U104 ( .A(n71), .B(n41), .Y(n57) );
  INVX1 U105 ( .A(n57), .Y(n58) );
  OR2X1 U106 ( .A(n71), .B(n26), .Y(n59) );
  INVX1 U107 ( .A(n59), .Y(n60) );
  OR2X1 U108 ( .A(1'b0), .B(M_DataMemStall), .Y(n61) );
  INVX1 U109 ( .A(n61), .Y(n62) );
  INVX2 U112 ( .A(D_RdValid), .Y(n70) );
endmodule

