
module fulladder1_15 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3, n4;

  XOR2X1 U1 ( .A(n3), .B(A), .Y(P) );
  AND2X2 U2 ( .A(B), .B(A), .Y(G) );
  INVX1 U3 ( .A(Cin), .Y(n4) );
  INVX1 U4 ( .A(B), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(n3) );
  XNOR2X1 U6 ( .A(P), .B(n4), .Y(S) );
endmodule


module fulladder1_14 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3;

  INVX1 U1 ( .A(A), .Y(n2) );
  XNOR2X1 U2 ( .A(n2), .B(B), .Y(P) );
  BUFX2 U3 ( .A(P), .Y(n3) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n3), .Y(S) );
endmodule


module fulladder1_13 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(n3), .Y(n1) );
  XOR2X1 U2 ( .A(n5), .B(n6), .Y(n2) );
  XOR2X1 U3 ( .A(Cin), .B(n2), .Y(S) );
  INVX1 U4 ( .A(B), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  BUFX2 U6 ( .A(n4), .Y(n5) );
  BUFX2 U7 ( .A(A), .Y(n6) );
  AND2X2 U8 ( .A(n4), .B(A), .Y(G) );
  XOR2X1 U9 ( .A(n1), .B(A), .Y(P) );
endmodule


module fulladder1_12 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  BUFX2 U1 ( .A(P), .Y(n1) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  XOR2X1 U4 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module fulladder1_11 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  INVX1 U1 ( .A(A), .Y(n1) );
  XNOR2X1 U2 ( .A(n1), .B(B), .Y(P) );
  BUFX2 U3 ( .A(P), .Y(n2) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U5 ( .A(Cin), .B(n2), .Y(S) );
endmodule


module fulladder1_10 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  BUFX2 U1 ( .A(P), .Y(n1) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module fulladder1_9 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  BUFX2 U1 ( .A(P), .Y(n1) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(P) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U4 ( .A(Cin), .B(n1), .Y(S) );
endmodule


module fulladder1_8 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n3;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  XNOR2X1 U2 ( .A(Cin), .B(n3), .Y(S) );
  INVX1 U3 ( .A(P), .Y(n3) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_7 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  XOR2X1 U1 ( .A(Cin), .B(P), .Y(S) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  INVX2 U4 ( .A(n1), .Y(P) );
endmodule


module fulladder1_6 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1;

  INVX2 U1 ( .A(n1), .Y(P) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(P), .Y(S) );
endmodule


module fulladder1_5 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2, n4, n5, n6, n7;

  INVX1 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  XOR2X1 U3 ( .A(B), .B(A), .Y(P) );
  INVX1 U4 ( .A(A), .Y(n4) );
  INVX1 U5 ( .A(n4), .Y(n5) );
  BUFX2 U6 ( .A(Cin), .Y(n6) );
  BUFX2 U7 ( .A(P), .Y(n7) );
  AND2X2 U8 ( .A(n5), .B(n2), .Y(G) );
  XOR2X1 U9 ( .A(n6), .B(n7), .Y(S) );
endmodule


module fulladder1_4 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2, n3;

  XNOR2X1 U1 ( .A(n2), .B(n3), .Y(S) );
  BUFX2 U2 ( .A(Cin), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(P) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U5 ( .A(A), .B(B), .Y(n3) );
endmodule


module fulladder1_3 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XNOR2X1 U1 ( .A(Cin), .B(n2), .Y(S) );
  AND2X2 U2 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n2) );
  INVX2 U4 ( .A(n2), .Y(P) );
endmodule


module fulladder1_2 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  BUFX2 U1 ( .A(Cin), .Y(n1) );
  XNOR2X1 U2 ( .A(n1), .B(n2), .Y(S) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(B), .B(A), .Y(n2) );
  INVX2 U5 ( .A(n2), .Y(P) );
endmodule


module fulladder1_1 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n2;

  XOR2X1 U1 ( .A(A), .B(B), .Y(P) );
  INVX2 U2 ( .A(P), .Y(n2) );
  XNOR2X1 U3 ( .A(Cin), .B(n2), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_0 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;
  wire   n1, n2;

  BUFX2 U1 ( .A(Cin), .Y(n1) );
  XNOR2X1 U2 ( .A(n1), .B(n2), .Y(S) );
  AND2X2 U3 ( .A(A), .B(B), .Y(G) );
  XNOR2X1 U4 ( .A(A), .B(B), .Y(n2) );
  INVX2 U5 ( .A(n2), .Y(P) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module mux4to1_16_3 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module mux4to1_16_2 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module mux4to1_16_1 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module mux4to1_16_0 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n69), .C(\InB<9> ), .D(n70), .Y(n106) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n103), .C(\InD<9> ), .D(n102), .Y(n107) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n69), .C(\InB<8> ), .D(n70), .Y(n100) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n103), .C(\InD<8> ), .D(n102), .Y(n101) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n69), .C(\InB<7> ), .D(n70), .Y(n98) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n103), .C(\InD<7> ), .D(n102), .Y(n99) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n69), .C(\InB<6> ), .D(n70), .Y(n96) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n103), .C(\InD<6> ), .D(n102), .Y(n97) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n69), .C(\InB<5> ), .D(n70), .Y(n94) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n103), .C(\InD<5> ), .D(n102), .Y(n95) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n69), .C(\InB<4> ), .D(n70), .Y(n92) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n103), .C(\InD<4> ), .D(n102), .Y(n93) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n69), .C(\InB<3> ), .D(n70), .Y(n90) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n103), .C(\InD<3> ), .D(n102), .Y(n91) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n69), .C(\InB<2> ), .D(n70), .Y(n88) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n103), .C(\InD<2> ), .D(n102), .Y(n89) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n69), .C(\InB<1> ), .D(n70), .Y(n86) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n103), .C(\InD<1> ), .D(n102), .Y(n87) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n69), .C(\InB<15> ), .D(n70), .Y(n84) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n103), .C(\InD<15> ), .D(n102), .Y(n85) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n69), .C(\InB<14> ), .D(n70), .Y(n82) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n103), .C(\InD<14> ), .D(n102), .Y(n83) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n69), .C(\InB<13> ), .D(n70), .Y(n80) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n103), .C(\InD<13> ), .D(n102), .Y(n81) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n69), .C(\InB<12> ), .D(n70), .Y(n78) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n103), .C(\InD<12> ), .D(n102), .Y(n79) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n69), .C(\InB<11> ), .D(n70), .Y(n76) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n103), .C(\InD<11> ), .D(n102), .Y(n77) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n69), .C(\InB<10> ), .D(n70), .Y(n74) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n103), .C(\InD<10> ), .D(n102), .Y(n75) );
  AOI22X1 U50 ( .A(\InA<0> ), .B(n69), .C(\InB<0> ), .D(n70), .Y(n72) );
  NOR2X1 U51 ( .A(n71), .B(\S<1> ), .Y(n104) );
  NOR2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n105) );
  AOI22X1 U53 ( .A(\InC<0> ), .B(n103), .C(\InD<0> ), .D(n102), .Y(n73) );
  AND2X1 U1 ( .A(\S<1> ), .B(n71), .Y(n103) );
  AND2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n102) );
  INVX1 U3 ( .A(\S<0> ), .Y(n71) );
  BUFX2 U4 ( .A(n105), .Y(n69) );
  BUFX2 U7 ( .A(n104), .Y(n70) );
  AND2X2 U10 ( .A(n73), .B(n72), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(\Out<0> ) );
  AND2X2 U16 ( .A(n75), .B(n74), .Y(n39) );
  INVX1 U19 ( .A(n39), .Y(\Out<10> ) );
  AND2X2 U22 ( .A(n77), .B(n76), .Y(n41) );
  INVX1 U25 ( .A(n41), .Y(\Out<11> ) );
  AND2X2 U28 ( .A(n79), .B(n78), .Y(n43) );
  INVX1 U31 ( .A(n43), .Y(\Out<12> ) );
  AND2X2 U34 ( .A(n81), .B(n80), .Y(n45) );
  INVX1 U37 ( .A(n45), .Y(\Out<13> ) );
  AND2X2 U40 ( .A(n83), .B(n82), .Y(n47) );
  INVX1 U43 ( .A(n47), .Y(\Out<14> ) );
  AND2X2 U46 ( .A(n85), .B(n84), .Y(n49) );
  INVX1 U49 ( .A(n49), .Y(\Out<15> ) );
  AND2X2 U54 ( .A(n87), .B(n86), .Y(n51) );
  INVX1 U55 ( .A(n51), .Y(\Out<1> ) );
  AND2X2 U56 ( .A(n89), .B(n88), .Y(n53) );
  INVX1 U57 ( .A(n53), .Y(\Out<2> ) );
  AND2X2 U58 ( .A(n91), .B(n90), .Y(n55) );
  INVX1 U59 ( .A(n55), .Y(\Out<3> ) );
  AND2X2 U60 ( .A(n93), .B(n92), .Y(n57) );
  INVX1 U61 ( .A(n57), .Y(\Out<4> ) );
  AND2X2 U62 ( .A(n95), .B(n94), .Y(n59) );
  INVX1 U63 ( .A(n59), .Y(\Out<5> ) );
  AND2X2 U64 ( .A(n97), .B(n96), .Y(n61) );
  INVX1 U65 ( .A(n61), .Y(\Out<6> ) );
  AND2X2 U66 ( .A(n99), .B(n98), .Y(n63) );
  INVX1 U67 ( .A(n63), .Y(\Out<7> ) );
  AND2X2 U68 ( .A(n101), .B(n100), .Y(n65) );
  INVX1 U69 ( .A(n65), .Y(\Out<8> ) );
  AND2X2 U70 ( .A(n107), .B(n106), .Y(n67) );
  INVX1 U71 ( .A(n67), .Y(\Out<9> ) );
endmodule


module demux1to8_0 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_1 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_2 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_3 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_4 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_5 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  NOR3X1 U4 ( .A(n7), .B(n4), .C(n6), .Y(Out7) );
  NOR3X1 U5 ( .A(n7), .B(n5), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n6), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(n5), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n6), .C(n7), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(n5), .C(n7), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n6), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out0) );
  INVX1 U1 ( .A(n6), .Y(n5) );
  INVX1 U2 ( .A(n9), .Y(n8) );
  INVX1 U3 ( .A(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(\S<0> ), .Y(n6) );
  INVX1 U13 ( .A(\S<2> ), .Y(n9) );
  AND2X1 U14 ( .A(In), .B(n9), .Y(n1) );
  INVX1 U15 ( .A(n1), .Y(n2) );
  AND2X1 U16 ( .A(n8), .B(In), .Y(n3) );
  INVX1 U17 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_6 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  NOR3X1 U4 ( .A(n7), .B(n4), .C(n6), .Y(Out7) );
  NOR3X1 U5 ( .A(n7), .B(n5), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n6), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(n5), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n6), .C(n7), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(n5), .C(n7), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n6), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out0) );
  INVX1 U1 ( .A(n6), .Y(n5) );
  INVX1 U2 ( .A(n9), .Y(n8) );
  INVX1 U3 ( .A(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(\S<0> ), .Y(n6) );
  INVX1 U13 ( .A(\S<2> ), .Y(n9) );
  AND2X1 U14 ( .A(In), .B(n9), .Y(n1) );
  INVX1 U15 ( .A(n1), .Y(n2) );
  AND2X1 U16 ( .A(n8), .B(In), .Y(n3) );
  INVX1 U17 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_7 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_8 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_9 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_10 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_11 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_12 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_13 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_14 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to8_15 ( In, .S({\S<2> , \S<1> , \S<0> }), Out0, Out1, Out2, Out3, 
        Out4, Out5, Out6, Out7 );
  input In, \S<2> , \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3, Out4, Out5, Out6, Out7;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR3X1 U4 ( .A(n6), .B(n4), .C(n5), .Y(Out7) );
  NOR3X1 U5 ( .A(n6), .B(\S<0> ), .C(n4), .Y(Out6) );
  NOR3X1 U6 ( .A(n5), .B(\S<1> ), .C(n4), .Y(Out5) );
  NOR3X1 U7 ( .A(n4), .B(\S<1> ), .C(\S<0> ), .Y(Out4) );
  NOR3X1 U9 ( .A(n2), .B(n5), .C(n6), .Y(Out3) );
  NOR3X1 U10 ( .A(n2), .B(\S<0> ), .C(n6), .Y(Out2) );
  NOR3X1 U11 ( .A(n2), .B(\S<1> ), .C(n5), .Y(Out1) );
  NOR3X1 U12 ( .A(n2), .B(\S<1> ), .C(\S<0> ), .Y(Out0) );
  INVX1 U1 ( .A(\S<1> ), .Y(n6) );
  INVX1 U2 ( .A(\S<0> ), .Y(n5) );
  INVX1 U3 ( .A(\S<2> ), .Y(n7) );
  AND2X1 U8 ( .A(In), .B(n7), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X1 U14 ( .A(\S<2> ), .B(In), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
endmodule


module demux1to4_17 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<0> ), .Y(n3) );
  INVX1 U2 ( .A(\S<1> ), .Y(n4) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_18 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<0> ), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(\S<1> ), .Y(n3) );
  INVX1 U4 ( .A(In), .Y(n4) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n3), .B(n2), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n3), .B(n5), .C(n1), .Y(Out2) );
  NOR3X1 U8 ( .A(n2), .B(n5), .C(\S<1> ), .Y(Out1) );
  NOR3X1 U9 ( .A(\S<1> ), .B(n1), .C(n4), .Y(Out0) );
endmodule


module demux1to4_19 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4;

  INVX1 U1 ( .A(\S<0> ), .Y(n1) );
  INVX1 U2 ( .A(\S<1> ), .Y(n2) );
  INVX1 U3 ( .A(In), .Y(n3) );
  INVX1 U4 ( .A(In), .Y(n4) );
  NOR3X1 U5 ( .A(n2), .B(n1), .C(n3), .Y(Out3) );
  NOR3X1 U6 ( .A(n2), .B(n3), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U7 ( .A(n1), .B(n3), .C(\S<1> ), .Y(Out1) );
  NOR3X1 U8 ( .A(\S<1> ), .B(\S<0> ), .C(n4), .Y(Out0) );
endmodule


module demux1to4_20 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<0> ), .Y(n3) );
  INVX1 U2 ( .A(\S<1> ), .Y(n4) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_21 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  INVX1 U2 ( .A(In), .Y(n9) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  AND2X1 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(Out0) );
  INVX1 U10 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_22 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<0> ), .Y(n3) );
  INVX1 U2 ( .A(\S<1> ), .Y(n4) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_23 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5;

  INVX1 U1 ( .A(\S<1> ), .Y(n4) );
  INVX1 U2 ( .A(\S<0> ), .Y(n3) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(In), .Y(n5) );
  NOR3X1 U6 ( .A(n4), .B(n3), .C(n5), .Y(Out3) );
  NOR3X1 U7 ( .A(n4), .B(n5), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U8 ( .A(n3), .B(n5), .C(\S<1> ), .Y(Out1) );
  AND2X2 U9 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_24 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11;

  OR2X2 U1 ( .A(n4), .B(\S<0> ), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(Out0) );
  AND2X2 U3 ( .A(In), .B(n10), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  AND2X1 U5 ( .A(n9), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  OR2X2 U7 ( .A(n6), .B(n10), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(Out2) );
  INVX1 U9 ( .A(\S<0> ), .Y(n9) );
  INVX1 U10 ( .A(In), .Y(n11) );
  INVX1 U11 ( .A(\S<1> ), .Y(n10) );
  NOR3X1 U12 ( .A(n10), .B(n9), .C(n11), .Y(Out3) );
  NOR3X1 U13 ( .A(n9), .B(n11), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_25 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10;

  OR2X2 U1 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X1 U3 ( .A(n8), .B(n7), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  OR2X2 U5 ( .A(n4), .B(n9), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out2) );
  INVX1 U7 ( .A(n10), .Y(n7) );
  INVX1 U8 ( .A(\S<0> ), .Y(n8) );
  AND2X2 U9 ( .A(n2), .B(In), .Y(Out0) );
  INVX1 U10 ( .A(\S<1> ), .Y(n9) );
  INVX1 U11 ( .A(In), .Y(n10) );
  NOR3X1 U12 ( .A(n9), .B(n8), .C(n10), .Y(Out3) );
  NOR3X1 U13 ( .A(n8), .B(n10), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_26 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n6;

  INVX4 U1 ( .A(\S<1> ), .Y(n5) );
  AND2X2 U2 ( .A(In), .B(n1), .Y(Out0) );
  AND2X2 U3 ( .A(n5), .B(n3), .Y(n1) );
  INVX1 U4 ( .A(n5), .Y(n4) );
  INVX1 U5 ( .A(n3), .Y(n2) );
  INVX1 U6 ( .A(In), .Y(n6) );
  INVX8 U7 ( .A(\S<0> ), .Y(n3) );
  NOR3X1 U8 ( .A(n5), .B(n3), .C(n6), .Y(Out3) );
  NOR3X1 U9 ( .A(n5), .B(n6), .C(n2), .Y(Out2) );
  NOR3X1 U10 ( .A(n3), .B(n6), .C(n4), .Y(Out1) );
endmodule


module demux1to4_27 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13;

  OR2X1 U1 ( .A(n6), .B(n12), .Y(n7) );
  INVX1 U2 ( .A(n12), .Y(n11) );
  OR2X2 U3 ( .A(n4), .B(n11), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(Out0) );
  AND2X2 U5 ( .A(n10), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  AND2X1 U7 ( .A(n10), .B(n9), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  INVX1 U9 ( .A(n7), .Y(Out2) );
  INVX1 U10 ( .A(\S<0> ), .Y(n10) );
  INVX1 U11 ( .A(n13), .Y(n9) );
  INVX1 U12 ( .A(\S<1> ), .Y(n12) );
  INVX1 U13 ( .A(In), .Y(n13) );
  NOR3X1 U14 ( .A(n12), .B(n10), .C(n13), .Y(Out3) );
  NOR3X1 U15 ( .A(n10), .B(n13), .C(n11), .Y(Out1) );
endmodule


module demux1to4_28 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11;

  OR2X2 U1 ( .A(\S<0> ), .B(n9), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X1 U3 ( .A(n8), .B(n7), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  OR2X2 U5 ( .A(n4), .B(n10), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(Out2) );
  INVX1 U7 ( .A(n10), .Y(n9) );
  AND2X2 U8 ( .A(In), .B(n2), .Y(Out0) );
  INVX1 U9 ( .A(\S<0> ), .Y(n8) );
  INVX1 U10 ( .A(\S<1> ), .Y(n10) );
  INVX1 U11 ( .A(n11), .Y(n7) );
  INVX1 U12 ( .A(In), .Y(n11) );
  NOR3X1 U13 ( .A(n10), .B(n8), .C(n11), .Y(Out3) );
  NOR3X1 U14 ( .A(n8), .B(n11), .C(n9), .Y(Out1) );
endmodule


module demux1to4_29 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n6, n8, n9, n10;

  INVX1 U1 ( .A(\S<1> ), .Y(n9) );
  INVX1 U2 ( .A(In), .Y(n10) );
  INVX1 U3 ( .A(n2), .Y(n1) );
  AND2X2 U4 ( .A(n8), .B(In), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(n3) );
  OR2X2 U6 ( .A(n3), .B(n9), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(Out2) );
  OR2X2 U8 ( .A(n1), .B(\S<1> ), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(Out0) );
  INVX1 U10 ( .A(\S<0> ), .Y(n8) );
  NOR3X1 U11 ( .A(n9), .B(n8), .C(n10), .Y(Out3) );
  NOR3X1 U12 ( .A(n8), .B(n10), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_30 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n7, n8, n9;

  OR2X1 U1 ( .A(n2), .B(n8), .Y(n3) );
  INVX1 U2 ( .A(In), .Y(n9) );
  INVX1 U3 ( .A(\S<1> ), .Y(n8) );
  AND2X2 U4 ( .A(n7), .B(In), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  INVX1 U6 ( .A(n3), .Y(Out2) );
  OR2X2 U7 ( .A(n2), .B(\S<1> ), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out0) );
  INVX1 U9 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U10 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U11 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_31 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n6, n7, n8, n9;

  INVX1 U1 ( .A(In), .Y(n9) );
  BUFX2 U2 ( .A(n6), .Y(n1) );
  AND2X1 U3 ( .A(n7), .B(In), .Y(n2) );
  INVX1 U4 ( .A(n2), .Y(n3) );
  OR2X2 U5 ( .A(n3), .B(n8), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(Out2) );
  NAND3X1 U7 ( .A(In), .B(n7), .C(n8), .Y(n6) );
  INVX2 U8 ( .A(n1), .Y(Out0) );
  INVX1 U9 ( .A(\S<0> ), .Y(n7) );
  INVX1 U10 ( .A(\S<1> ), .Y(n8) );
  NOR3X1 U11 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U12 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_32 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  INVX1 U2 ( .A(In), .Y(n9) );
  OR2X1 U3 ( .A(n4), .B(n8), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(Out2) );
  AND2X1 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X2 U7 ( .A(n4), .B(\S<1> ), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out0) );
  INVX1 U9 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U10 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U11 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_15 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  AND2X2 U2 ( .A(In), .B(\S<1> ), .Y(n11) );
  AND2X2 U3 ( .A(In), .B(\S<0> ), .Y(n5) );
  OR2X1 U4 ( .A(n12), .B(n13), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(Out3) );
  OR2X1 U6 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(n4) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  OR2X2 U9 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(Out1) );
  OR2X1 U11 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Out2) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_14 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n5, n6, n7, n8, n10, n12, n13, n14;

  INVX1 U1 ( .A(\S<0> ), .Y(n14) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(\S<0> ), .B(n1), .Y(n6) );
  AND2X2 U4 ( .A(n1), .B(\S<1> ), .Y(n12) );
  OR2X1 U5 ( .A(n13), .B(n14), .Y(n2) );
  INVX1 U6 ( .A(n2), .Y(Out3) );
  OR2X1 U7 ( .A(\S<1> ), .B(\S<0> ), .Y(n4) );
  INVX1 U8 ( .A(n4), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(n7) );
  OR2X2 U10 ( .A(n7), .B(\S<1> ), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(Out1) );
  OR2X1 U12 ( .A(n13), .B(\S<0> ), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(Out2) );
  INVX1 U14 ( .A(n12), .Y(n13) );
  AND2X2 U15 ( .A(n5), .B(In), .Y(Out0) );
endmodule


module demux1to4_13 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n14, n15;

  INVX1 U1 ( .A(\S<0> ), .Y(n15) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X1 U3 ( .A(n14), .B(n15), .Y(n2) );
  INVX1 U4 ( .A(\S<1> ), .Y(n14) );
  OR2X1 U5 ( .A(n12), .B(n15), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(Out3) );
  AND2X2 U7 ( .A(n1), .B(\S<0> ), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  OR2X2 U9 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(Out1) );
  OR2X1 U11 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(Out2) );
  AND2X2 U13 ( .A(n1), .B(\S<1> ), .Y(n11) );
  INVX1 U14 ( .A(n11), .Y(n12) );
  AND2X2 U15 ( .A(In), .B(n2), .Y(Out0) );
endmodule


module demux1to4_12 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n5, n6, n7, n9, n11, n12, n13, n14, n15;

  INVX1 U1 ( .A(\S<1> ), .Y(n13) );
  INVX1 U2 ( .A(\S<0> ), .Y(n14) );
  BUFX2 U3 ( .A(In), .Y(n1) );
  AND2X2 U4 ( .A(n1), .B(\S<1> ), .Y(n11) );
  AND2X2 U5 ( .A(\S<0> ), .B(n1), .Y(n5) );
  AND2X2 U6 ( .A(n15), .B(In), .Y(Out0) );
  OR2X1 U7 ( .A(n12), .B(n14), .Y(n3) );
  INVX1 U8 ( .A(n3), .Y(Out3) );
  INVX1 U9 ( .A(n5), .Y(n6) );
  OR2X2 U10 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U11 ( .A(n7), .Y(Out1) );
  OR2X1 U12 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U13 ( .A(n9), .Y(Out2) );
  INVX1 U14 ( .A(n11), .Y(n12) );
  AND2X2 U15 ( .A(n13), .B(n14), .Y(n15) );
endmodule


module demux1to4_11 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  OR2X1 U2 ( .A(n12), .B(n13), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X1 U4 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  AND2X1 U6 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_10 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9, n10;

  INVX1 U1 ( .A(\S<0> ), .Y(n9) );
  INVX1 U2 ( .A(In), .Y(n10) );
  OR2X1 U3 ( .A(n8), .B(n9), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(Out3) );
  OR2X1 U5 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X1 U7 ( .A(n8), .B(\S<0> ), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  AND2X1 U9 ( .A(In), .B(\S<1> ), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(n8) );
  NOR3X1 U11 ( .A(n9), .B(\S<1> ), .C(n10), .Y(Out1) );
  AND2X2 U12 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_9 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  OR2X1 U2 ( .A(n12), .B(n13), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X1 U4 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  AND2X1 U6 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_8 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13, n14;

  INVX1 U1 ( .A(n14), .Y(n13) );
  OR2X1 U2 ( .A(n12), .B(n14), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X1 U4 ( .A(\S<1> ), .B(n13), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  AND2X1 U6 ( .A(n13), .B(In), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(n13), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  INVX1 U14 ( .A(\S<0> ), .Y(n14) );
  AND2X2 U15 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_7 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n6, n7, n9, n11, n12, n13;

  INVX1 U1 ( .A(\S<0> ), .Y(n13) );
  OR2X1 U2 ( .A(n12), .B(n13), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out3) );
  OR2X1 U4 ( .A(\S<1> ), .B(\S<0> ), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  AND2X1 U6 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  OR2X2 U8 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(Out1) );
  OR2X1 U10 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out2) );
  AND2X1 U12 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AND2X2 U14 ( .A(In), .B(n4), .Y(Out0) );
endmodule


module demux1to4_6 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15;

  BUFX2 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(n1), .B(\S<1> ), .Y(n12) );
  AND2X2 U3 ( .A(n1), .B(n14), .Y(n6) );
  OR2X1 U4 ( .A(n13), .B(n15), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(Out3) );
  OR2X1 U6 ( .A(\S<1> ), .B(n14), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n5) );
  INVX1 U8 ( .A(n6), .Y(n7) );
  OR2X2 U9 ( .A(n7), .B(\S<1> ), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(Out1) );
  OR2X1 U11 ( .A(n13), .B(n14), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(Out2) );
  INVX1 U13 ( .A(n12), .Y(n13) );
  INVX1 U14 ( .A(n15), .Y(n14) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
  AND2X2 U16 ( .A(n5), .B(In), .Y(Out0) );
endmodule


module demux1to4_5 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(\S<0> ), .Y(n4) );
  INVX1 U2 ( .A(\S<1> ), .Y(n5) );
  BUFX2 U3 ( .A(In), .Y(n1) );
  OR2X1 U4 ( .A(\S<0> ), .B(\S<1> ), .Y(n2) );
  INVX1 U5 ( .A(n2), .Y(n3) );
  INVX1 U6 ( .A(n1), .Y(n6) );
  NOR3X1 U7 ( .A(n5), .B(n4), .C(n6), .Y(Out3) );
  NOR3X1 U8 ( .A(n5), .B(n6), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U9 ( .A(n4), .B(n6), .C(\S<1> ), .Y(Out1) );
  AND2X2 U10 ( .A(n3), .B(In), .Y(Out0) );
endmodule


module demux1to4_4 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(\S<0> ), .Y(n4) );
  INVX1 U2 ( .A(\S<1> ), .Y(n5) );
  OR2X1 U3 ( .A(\S<0> ), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  BUFX2 U5 ( .A(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n6) );
  NOR3X1 U7 ( .A(n5), .B(n4), .C(n6), .Y(Out3) );
  NOR3X1 U8 ( .A(n5), .B(n6), .C(\S<0> ), .Y(Out2) );
  NOR3X1 U9 ( .A(n4), .B(n6), .C(\S<1> ), .Y(Out1) );
  AND2X2 U10 ( .A(n2), .B(In), .Y(Out0) );
endmodule


module demux1to4_3 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(\S<1> ), .Y(n8) );
  INVX1 U2 ( .A(In), .Y(n9) );
  OR2X2 U3 ( .A(n4), .B(\S<1> ), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(Out0) );
  AND2X2 U5 ( .A(n7), .B(In), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  OR2X1 U7 ( .A(n4), .B(n8), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(Out2) );
  INVX8 U9 ( .A(\S<0> ), .Y(n7) );
  NOR3X1 U10 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U11 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_2 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n7, n8, n9;

  INVX2 U1 ( .A(\S<0> ), .Y(n7) );
  INVX1 U2 ( .A(In), .Y(n9) );
  INVX1 U3 ( .A(\S<1> ), .Y(n8) );
  AND2X2 U4 ( .A(n7), .B(In), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  OR2X2 U6 ( .A(n2), .B(\S<1> ), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(Out0) );
  OR2X1 U8 ( .A(n2), .B(n8), .Y(n5) );
  INVX1 U9 ( .A(n5), .Y(Out2) );
  NOR3X1 U10 ( .A(n8), .B(n7), .C(n9), .Y(Out3) );
  NOR3X1 U11 ( .A(n7), .B(n9), .C(\S<1> ), .Y(Out1) );
endmodule


module demux1to4_1 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n3, n4, n5, n7, n8, n9, n11, n13, n14, n15;

  INVX1 U1 ( .A(\S<0> ), .Y(n15) );
  OR2X2 U2 ( .A(n4), .B(\S<1> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(Out0) );
  AND2X2 U4 ( .A(n15), .B(In), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  OR2X1 U6 ( .A(n14), .B(n15), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(Out3) );
  AND2X1 U8 ( .A(\S<0> ), .B(In), .Y(n7) );
  INVX1 U9 ( .A(n7), .Y(n8) );
  OR2X2 U10 ( .A(n8), .B(\S<1> ), .Y(n9) );
  INVX1 U11 ( .A(n9), .Y(Out1) );
  OR2X1 U12 ( .A(n14), .B(\S<0> ), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(Out2) );
  AND2X1 U14 ( .A(In), .B(\S<1> ), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(n14) );
endmodule


module demux1to4_0 ( In, .S({\S<1> , \S<0> }), Out0, Out1, Out2, Out3 );
  input In, \S<1> , \S<0> ;
  output Out0, Out1, Out2, Out3;
  wire   n1, n2, n3, n5, n6, n7, n9, n11, n12, n13, n15;

  AND2X2 U1 ( .A(n15), .B(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  OR2X1 U3 ( .A(n12), .B(n15), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(Out3) );
  AND2X2 U5 ( .A(\S<0> ), .B(In), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(n6) );
  OR2X2 U7 ( .A(n6), .B(\S<1> ), .Y(n7) );
  INVX1 U8 ( .A(n7), .Y(Out1) );
  OR2X1 U9 ( .A(n12), .B(\S<0> ), .Y(n9) );
  INVX1 U10 ( .A(n9), .Y(Out2) );
  AND2X1 U11 ( .A(In), .B(\S<1> ), .Y(n11) );
  INVX1 U12 ( .A(n11), .Y(n12) );
  OR2X2 U13 ( .A(n2), .B(\S<1> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(Out0) );
  INVX1 U15 ( .A(\S<0> ), .Y(n15) );
endmodule


module cla4_3 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79;

  fulladder1_15 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n76), .G(n72) );
  fulladder1_14 \fa[1]  ( .A(n54), .B(\B<1> ), .Cin(n37), .S(\S<1> ), .P(n77), 
        .G(n73) );
  fulladder1_13 \fa[2]  ( .A(n55), .B(\B<2> ), .Cin(n71), .S(\S<2> ), .P(n78), 
        .G(n74) );
  fulladder1_12 \fa[3]  ( .A(n7), .B(\B<3> ), .Cin(n70), .S(\S<3> ), .P(n79), 
        .G(n75) );
  BUFX2 U1 ( .A(n38), .Y(n1) );
  INVX1 U2 ( .A(n8), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
  AND2X2 U4 ( .A(n30), .B(n11), .Y(n4) );
  INVX1 U5 ( .A(n70), .Y(n67) );
  XNOR2X1 U6 ( .A(\B<1> ), .B(n49), .Y(n11) );
  INVX1 U7 ( .A(\A<0> ), .Y(n9) );
  INVX1 U8 ( .A(n59), .Y(n5) );
  XNOR2X1 U9 ( .A(n45), .B(n55), .Y(n57) );
  INVX1 U10 ( .A(n38), .Y(n6) );
  INVX8 U11 ( .A(n12), .Y(n7) );
  INVX4 U12 ( .A(\A<3> ), .Y(n12) );
  AND2X2 U13 ( .A(\B<0> ), .B(\A<0> ), .Y(n17) );
  XNOR2X1 U14 ( .A(n12), .B(\B<3> ), .Y(n52) );
  XNOR2X1 U15 ( .A(\B<0> ), .B(n9), .Y(n8) );
  INVX1 U16 ( .A(n11), .Y(n59) );
  INVX1 U17 ( .A(n16), .Y(n10) );
  INVX1 U18 ( .A(n71), .Y(n58) );
  INVX1 U19 ( .A(\B<2> ), .Y(n45) );
  AND2X2 U20 ( .A(\A<3> ), .B(\B<3> ), .Y(n32) );
  OR2X2 U21 ( .A(n18), .B(n20), .Y(n13) );
  INVX1 U22 ( .A(n13), .Y(PG) );
  AND2X2 U23 ( .A(n75), .B(n32), .Y(n15) );
  INVX1 U24 ( .A(n15), .Y(n16) );
  OR2X2 U25 ( .A(n22), .B(n21), .Y(n18) );
  AND2X2 U26 ( .A(n76), .B(n65), .Y(n19) );
  INVX1 U27 ( .A(n19), .Y(n20) );
  INVX1 U28 ( .A(n33), .Y(n21) );
  AND2X2 U29 ( .A(n77), .B(n5), .Y(n33) );
  BUFX2 U30 ( .A(n66), .Y(n22) );
  BUFX2 U31 ( .A(n62), .Y(n23) );
  BUFX2 U32 ( .A(n64), .Y(n24) );
  AND2X2 U33 ( .A(n29), .B(n6), .Y(n25) );
  INVX1 U34 ( .A(n25), .Y(n26) );
  AND2X2 U35 ( .A(n78), .B(n57), .Y(n27) );
  INVX1 U36 ( .A(n27), .Y(n28) );
  INVX1 U37 ( .A(n27), .Y(n29) );
  AND2X2 U38 ( .A(n17), .B(n72), .Y(n30) );
  INVX1 U39 ( .A(n30), .Y(n31) );
  INVX1 U40 ( .A(n60), .Y(n34) );
  INVX1 U41 ( .A(n34), .Y(n35) );
  AND2X2 U42 ( .A(n31), .B(n56), .Y(n36) );
  INVX1 U43 ( .A(n36), .Y(n37) );
  INVX1 U44 ( .A(n61), .Y(n38) );
  INVX1 U45 ( .A(n1), .Y(n39) );
  INVX1 U46 ( .A(n16), .Y(n40) );
  INVX1 U47 ( .A(n40), .Y(n41) );
  INVX1 U48 ( .A(n65), .Y(n42) );
  INVX1 U49 ( .A(n46), .Y(n43) );
  BUFX2 U50 ( .A(\B<1> ), .Y(n44) );
  INVX1 U51 ( .A(n77), .Y(n46) );
  INVX1 U52 ( .A(n55), .Y(n47) );
  INVX1 U53 ( .A(n47), .Y(n48) );
  INVX1 U54 ( .A(n54), .Y(n49) );
  INVX1 U55 ( .A(n49), .Y(n50) );
  BUFX2 U56 ( .A(\B<2> ), .Y(n51) );
  AND2X2 U57 ( .A(n52), .B(n79), .Y(n53) );
  INVX1 U58 ( .A(n53), .Y(n68) );
  BUFX4 U59 ( .A(\A<1> ), .Y(n54) );
  BUFX4 U60 ( .A(\A<2> ), .Y(n55) );
  INVX1 U61 ( .A(n28), .Y(n65) );
  NAND3X1 U62 ( .A(Cin), .B(n3), .C(n76), .Y(n56) );
  NAND3X1 U63 ( .A(n50), .B(n44), .C(n73), .Y(n60) );
  OAI21X1 U64 ( .A(n21), .B(n36), .C(n35), .Y(n71) );
  NAND3X1 U65 ( .A(n48), .B(n51), .C(n74), .Y(n61) );
  OAI21X1 U66 ( .A(n42), .B(n58), .C(n39), .Y(n70) );
  AOI21X1 U67 ( .A(n4), .B(n43), .C(n10), .Y(n64) );
  AND2X2 U68 ( .A(n39), .B(n35), .Y(n63) );
  AOI21X1 U69 ( .A(n26), .B(n53), .C(n40), .Y(n62) );
  AOI21X1 U70 ( .A(n63), .B(n24), .C(n23), .Y(GG) );
  NAND3X1 U71 ( .A(n52), .B(n8), .C(n79), .Y(n66) );
  OAI21X1 U72 ( .A(n68), .B(n67), .C(n41), .Y(Cout) );
endmodule


module cla4_2 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  fulladder1_11 \fa[0]  ( .A(n37), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(n73), 
        .G(n69) );
  fulladder1_10 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n9), .S(\S<1> ), .P(n74), .G(n70) );
  fulladder1_9 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n24), .S(\S<2> ), .P(n75), .G(n71) );
  fulladder1_8 \fa[3]  ( .A(n49), .B(\B<3> ), .Cin(n68), .S(\S<3> ), .P(n76), 
        .G(n72) );
  INVX1 U1 ( .A(n33), .Y(n54) );
  INVX1 U2 ( .A(\A<2> ), .Y(n3) );
  XOR2X1 U3 ( .A(n41), .B(\B<0> ), .Y(n1) );
  BUFX2 U4 ( .A(\B<2> ), .Y(n2) );
  XNOR2X1 U5 ( .A(n3), .B(\B<2> ), .Y(n50) );
  XNOR2X1 U6 ( .A(\B<1> ), .B(n42), .Y(n51) );
  INVX2 U7 ( .A(\A<1> ), .Y(n42) );
  BUFX2 U8 ( .A(n73), .Y(n4) );
  INVX1 U9 ( .A(n30), .Y(n5) );
  OR2X2 U10 ( .A(n13), .B(n17), .Y(n6) );
  INVX1 U11 ( .A(n6), .Y(PG) );
  AND2X2 U12 ( .A(n38), .B(n5), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  AND2X2 U14 ( .A(n47), .B(n31), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  AND2X2 U16 ( .A(n1), .B(n45), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  BUFX2 U18 ( .A(n62), .Y(n14) );
  AND2X2 U19 ( .A(n75), .B(n50), .Y(n15) );
  INVX1 U20 ( .A(n63), .Y(n16) );
  INVX1 U21 ( .A(n16), .Y(n17) );
  AND2X1 U22 ( .A(n15), .B(n36), .Y(n18) );
  AND2X1 U23 ( .A(n33), .B(n28), .Y(n19) );
  INVX1 U24 ( .A(n19), .Y(n20) );
  OR2X1 U25 ( .A(n54), .B(n58), .Y(n21) );
  INVX1 U26 ( .A(n21), .Y(n22) );
  INVX1 U27 ( .A(n67), .Y(n23) );
  INVX1 U28 ( .A(n23), .Y(n24) );
  INVX1 U29 ( .A(n53), .Y(n25) );
  INVX1 U30 ( .A(n25), .Y(n26) );
  INVX1 U31 ( .A(n56), .Y(n27) );
  INVX1 U32 ( .A(n27), .Y(n28) );
  BUFX2 U33 ( .A(n64), .Y(n29) );
  INVX1 U34 ( .A(n55), .Y(n30) );
  INVX1 U35 ( .A(n30), .Y(n31) );
  INVX1 U36 ( .A(n57), .Y(n32) );
  INVX1 U37 ( .A(n32), .Y(n33) );
  INVX1 U38 ( .A(n52), .Y(n34) );
  INVX1 U39 ( .A(n34), .Y(n35) );
  OAI21X1 U40 ( .A(n60), .B(n15), .C(n45), .Y(n61) );
  INVX1 U41 ( .A(n28), .Y(n60) );
  NAND3X1 U42 ( .A(n1), .B(n4), .C(Cin), .Y(n55) );
  AND2X2 U43 ( .A(n74), .B(n51), .Y(n36) );
  INVX1 U44 ( .A(n40), .Y(n37) );
  BUFX2 U45 ( .A(n26), .Y(n38) );
  INVX1 U46 ( .A(n40), .Y(n41) );
  INVX1 U47 ( .A(n36), .Y(n39) );
  INVX1 U48 ( .A(\A<0> ), .Y(n40) );
  INVX1 U49 ( .A(n42), .Y(n43) );
  BUFX2 U50 ( .A(\B<1> ), .Y(n44) );
  AND2X2 U51 ( .A(n76), .B(n59), .Y(n45) );
  INVX1 U52 ( .A(n45), .Y(n66) );
  AND2X2 U53 ( .A(n11), .B(n46), .Y(n68) );
  OR2X2 U54 ( .A(n34), .B(n18), .Y(n46) );
  AND2X2 U55 ( .A(n38), .B(n35), .Y(n47) );
  INVX1 U56 ( .A(n26), .Y(n58) );
  BUFX2 U57 ( .A(n68), .Y(n48) );
  BUFX4 U58 ( .A(\A<3> ), .Y(n49) );
  INVX1 U59 ( .A(n48), .Y(n65) );
  NAND3X1 U60 ( .A(n41), .B(\B<0> ), .C(n69), .Y(n53) );
  NAND3X1 U61 ( .A(n43), .B(n44), .C(n70), .Y(n57) );
  NAND3X1 U62 ( .A(\A<2> ), .B(n2), .C(n71), .Y(n56) );
  AOI21X1 U63 ( .A(n15), .B(n54), .C(n60), .Y(n52) );
  AOI22X1 U64 ( .A(n33), .B(n39), .C(n31), .D(n22), .Y(n67) );
  AOI21X1 U65 ( .A(n58), .B(n36), .C(n20), .Y(n62) );
  XOR2X1 U66 ( .A(n49), .B(\B<3> ), .Y(n59) );
  NAND3X1 U67 ( .A(n49), .B(\B<3> ), .C(n72), .Y(n64) );
  OAI21X1 U68 ( .A(n14), .B(n61), .C(n29), .Y(GG) );
  NAND3X1 U69 ( .A(n73), .B(n36), .C(n15), .Y(n63) );
  OAI21X1 U70 ( .A(n66), .B(n65), .C(n29), .Y(Cout) );
endmodule


module cla4_1 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97;

  fulladder1_7 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(n67), .S(\S<0> ), .P(n94), .G(n90) );
  fulladder1_6 \fa[1]  ( .A(n69), .B(\B<1> ), .Cin(n49), .S(\S<1> ), .P(n95), 
        .G(n91) );
  fulladder1_5 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n88), .S(\S<2> ), .P(n96), .G(n92) );
  fulladder1_4 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n89), .S(\S<3> ), .P(n97), .G(n93) );
  INVX1 U1 ( .A(n61), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U3 ( .A(n68), .B(n21), .Y(n3) );
  AND2X2 U4 ( .A(n94), .B(n79), .Y(n55) );
  INVX1 U5 ( .A(n66), .Y(n67) );
  NOR3X1 U6 ( .A(n5), .B(n12), .C(n76), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n80) );
  INVX8 U8 ( .A(n94), .Y(n5) );
  AND2X2 U9 ( .A(n8), .B(n30), .Y(n6) );
  OR2X2 U10 ( .A(n6), .B(n7), .Y(n14) );
  AND2X1 U11 ( .A(n53), .B(n50), .Y(n7) );
  AND2X1 U12 ( .A(n19), .B(n53), .Y(n8) );
  BUFX2 U13 ( .A(\B<2> ), .Y(n9) );
  INVX1 U14 ( .A(n16), .Y(n10) );
  XOR2X1 U15 ( .A(\B<2> ), .B(\A<2> ), .Y(n61) );
  INVX1 U16 ( .A(n74), .Y(n11) );
  INVX1 U17 ( .A(n68), .Y(n12) );
  INVX1 U18 ( .A(n12), .Y(n13) );
  INVX1 U19 ( .A(Cin), .Y(n74) );
  INVX1 U20 ( .A(n14), .Y(GG) );
  AND2X2 U21 ( .A(n38), .B(n91), .Y(n16) );
  AND2X2 U22 ( .A(n28), .B(n32), .Y(n17) );
  INVX1 U23 ( .A(n17), .Y(n18) );
  AND2X2 U24 ( .A(n52), .B(n26), .Y(n19) );
  AND2X2 U25 ( .A(\A<0> ), .B(\B<0> ), .Y(n20) );
  AND2X2 U26 ( .A(n20), .B(n90), .Y(n21) );
  INVX1 U27 ( .A(n21), .Y(n22) );
  AND2X2 U28 ( .A(n65), .B(n39), .Y(n23) );
  OR2X2 U29 ( .A(n34), .B(n80), .Y(n24) );
  INVX1 U30 ( .A(n24), .Y(PG) );
  BUFX2 U31 ( .A(n77), .Y(n26) );
  AND2X2 U32 ( .A(\B<1> ), .B(n59), .Y(n27) );
  INVX1 U33 ( .A(n27), .Y(n28) );
  AND2X2 U34 ( .A(n3), .B(n64), .Y(n29) );
  INVX1 U35 ( .A(n29), .Y(n30) );
  AND2X2 U36 ( .A(n60), .B(n69), .Y(n31) );
  INVX1 U37 ( .A(n31), .Y(n32) );
  AND2X2 U38 ( .A(n79), .B(n37), .Y(n33) );
  INVX1 U39 ( .A(n33), .Y(n34) );
  OR2X2 U40 ( .A(n21), .B(n67), .Y(n35) );
  INVX1 U41 ( .A(n35), .Y(n36) );
  AND2X2 U42 ( .A(n75), .B(n97), .Y(n37) );
  AND2X2 U43 ( .A(\B<1> ), .B(n69), .Y(n38) );
  AND2X2 U44 ( .A(n22), .B(n10), .Y(n39) );
  INVX1 U45 ( .A(n71), .Y(n40) );
  INVX1 U46 ( .A(n40), .Y(n41) );
  AND2X1 U47 ( .A(n10), .B(n12), .Y(n42) );
  INVX1 U48 ( .A(n42), .Y(n43) );
  BUFX2 U49 ( .A(n81), .Y(n44) );
  BUFX2 U50 ( .A(n86), .Y(n45) );
  AND2X1 U51 ( .A(n10), .B(n65), .Y(n46) );
  INVX1 U52 ( .A(n46), .Y(n47) );
  INVX1 U53 ( .A(n87), .Y(n48) );
  INVX1 U54 ( .A(n48), .Y(n49) );
  INVX1 U55 ( .A(n37), .Y(n50) );
  INVX1 U56 ( .A(n82), .Y(n51) );
  INVX1 U57 ( .A(n51), .Y(n52) );
  BUFX2 U58 ( .A(n85), .Y(n53) );
  INVX1 U59 ( .A(n39), .Y(n54) );
  INVX1 U60 ( .A(n55), .Y(n56) );
  INVX1 U61 ( .A(n76), .Y(n57) );
  INVX1 U62 ( .A(n78), .Y(n58) );
  INVX1 U63 ( .A(n69), .Y(n59) );
  INVX1 U64 ( .A(\B<1> ), .Y(n60) );
  XNOR2X1 U65 ( .A(n62), .B(\A<3> ), .Y(n75) );
  INVX1 U66 ( .A(\B<3> ), .Y(n62) );
  INVX1 U67 ( .A(n62), .Y(n63) );
  AND2X2 U68 ( .A(n96), .B(n2), .Y(n64) );
  INVX1 U69 ( .A(n64), .Y(n76) );
  BUFX2 U70 ( .A(n52), .Y(n65) );
  INVX1 U71 ( .A(Cin), .Y(n66) );
  INVX1 U72 ( .A(n65), .Y(n83) );
  INVX1 U73 ( .A(n50), .Y(n78) );
  AND2X2 U74 ( .A(n18), .B(n95), .Y(n68) );
  BUFX4 U75 ( .A(\A<1> ), .Y(n69) );
  NAND3X1 U76 ( .A(n9), .B(\A<2> ), .C(n92), .Y(n82) );
  XNOR2X1 U77 ( .A(\A<0> ), .B(\B<0> ), .Y(n70) );
  INVX2 U78 ( .A(n70), .Y(n79) );
  AOI22X1 U79 ( .A(n65), .B(n76), .C(n23), .D(n56), .Y(n71) );
  OAI21X1 U80 ( .A(n13), .B(n47), .C(n41), .Y(n72) );
  AOI21X1 U81 ( .A(n74), .B(n23), .C(n72), .Y(n89) );
  OAI21X1 U82 ( .A(n55), .B(n54), .C(n43), .Y(n73) );
  AOI21X1 U83 ( .A(n74), .B(n39), .C(n73), .Y(n88) );
  AOI21X1 U84 ( .A(n22), .B(n56), .C(n36), .Y(n87) );
  NAND3X1 U85 ( .A(\A<3> ), .B(n63), .C(n93), .Y(n85) );
  NAND3X1 U86 ( .A(n61), .B(n16), .C(n96), .Y(n77) );
  AOI21X1 U87 ( .A(n11), .B(n55), .C(n21), .Y(n81) );
  OAI21X1 U88 ( .A(n44), .B(n12), .C(n10), .Y(n84) );
  AOI21X1 U89 ( .A(n57), .B(n84), .C(n83), .Y(n86) );
  OAI21X1 U90 ( .A(n45), .B(n58), .C(n53), .Y(Cout) );
endmodule


module cla4_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  fulladder1_3 \fa[0]  ( .A(\A<0> ), .B(n43), .Cin(n48), .S(\S<0> ), .P(n74), 
        .G(n70) );
  fulladder1_2 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n68), .S(\S<1> ), .P(n75), .G(n71) );
  fulladder1_1 \fa[2]  ( .A(\A<2> ), .B(n47), .Cin(n1), .S(\S<2> ), .P(n76), 
        .G(n72) );
  fulladder1_0 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n69), .S(\S<3> ), .P(n77), .G(n73) );
  INVX1 U1 ( .A(n21), .Y(n1) );
  INVX1 U2 ( .A(n54), .Y(n2) );
  AND2X2 U3 ( .A(n74), .B(n61), .Y(n38) );
  INVX2 U4 ( .A(n46), .Y(n47) );
  OR2X2 U5 ( .A(n11), .B(n26), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(PG) );
  AND2X2 U7 ( .A(n37), .B(n32), .Y(n5) );
  INVX1 U8 ( .A(n5), .Y(n6) );
  AND2X2 U9 ( .A(n75), .B(n51), .Y(n7) );
  AND2X2 U10 ( .A(Cin), .B(n13), .Y(n8) );
  INVX1 U11 ( .A(n8), .Y(n9) );
  AND2X2 U12 ( .A(n61), .B(n34), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(n11) );
  OR2X2 U14 ( .A(n39), .B(n42), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(n13) );
  OR2X2 U16 ( .A(n2), .B(n40), .Y(n14) );
  INVX1 U17 ( .A(n14), .Y(n15) );
  AND2X2 U18 ( .A(n44), .B(n6), .Y(n16) );
  INVX1 U19 ( .A(n16), .Y(n17) );
  INVX1 U20 ( .A(n16), .Y(n18) );
  AND2X2 U21 ( .A(n41), .B(n17), .Y(n19) );
  INVX1 U22 ( .A(n19), .Y(n20) );
  AND2X2 U23 ( .A(n56), .B(n9), .Y(n21) );
  INVX1 U24 ( .A(n21), .Y(n22) );
  AND2X2 U25 ( .A(n34), .B(n66), .Y(n23) );
  INVX1 U26 ( .A(n23), .Y(n24) );
  INVX1 U27 ( .A(n63), .Y(n25) );
  INVX1 U28 ( .A(n25), .Y(n26) );
  INVX1 U29 ( .A(n60), .Y(n27) );
  INVX1 U30 ( .A(n27), .Y(n28) );
  INVX1 U31 ( .A(n55), .Y(n29) );
  INVX1 U32 ( .A(n29), .Y(n30) );
  AND2X1 U33 ( .A(n76), .B(n49), .Y(n31) );
  INVX1 U34 ( .A(n31), .Y(n32) );
  BUFX2 U35 ( .A(n67), .Y(n33) );
  AND2X1 U36 ( .A(n77), .B(n59), .Y(n34) );
  INVX1 U37 ( .A(n34), .Y(n35) );
  INVX1 U38 ( .A(n64), .Y(n36) );
  INVX1 U39 ( .A(n36), .Y(n37) );
  INVX1 U40 ( .A(n38), .Y(n39) );
  INVX1 U41 ( .A(n41), .Y(n40) );
  BUFX2 U42 ( .A(n57), .Y(n41) );
  INVX1 U43 ( .A(n7), .Y(n42) );
  BUFX4 U44 ( .A(\B<0> ), .Y(n43) );
  OR2X1 U45 ( .A(n29), .B(n36), .Y(n44) );
  INVX1 U46 ( .A(n62), .Y(n45) );
  INVX1 U47 ( .A(\B<2> ), .Y(n46) );
  INVX1 U48 ( .A(n32), .Y(n62) );
  INVX1 U49 ( .A(n54), .Y(n48) );
  INVX1 U50 ( .A(Cin), .Y(n54) );
  INVX1 U51 ( .A(n22), .Y(n65) );
  NAND3X1 U52 ( .A(\A<1> ), .B(\B<1> ), .C(n71), .Y(n55) );
  NAND3X1 U53 ( .A(\A<2> ), .B(n47), .C(n72), .Y(n64) );
  XOR2X1 U54 ( .A(n47), .B(\A<2> ), .Y(n49) );
  NAND3X1 U55 ( .A(\A<0> ), .B(n43), .C(n70), .Y(n57) );
  XNOR2X1 U56 ( .A(\A<0> ), .B(n43), .Y(n50) );
  INVX2 U57 ( .A(n50), .Y(n61) );
  XOR2X1 U58 ( .A(\B<1> ), .B(\A<1> ), .Y(n51) );
  OAI21X1 U59 ( .A(n42), .B(n5), .C(n18), .Y(n52) );
  OAI21X1 U60 ( .A(n20), .B(n38), .C(n52), .Y(n53) );
  AOI21X1 U61 ( .A(n54), .B(n19), .C(n53), .Y(n69) );
  OAI21X1 U62 ( .A(n41), .B(n42), .C(n30), .Y(n58) );
  INVX2 U63 ( .A(n58), .Y(n56) );
  AOI21X1 U64 ( .A(n41), .B(n39), .C(n15), .Y(n68) );
  AOI21X1 U65 ( .A(n62), .B(n58), .C(n36), .Y(n60) );
  XOR2X1 U66 ( .A(\B<3> ), .B(\A<3> ), .Y(n59) );
  NAND3X1 U67 ( .A(\A<3> ), .B(\B<3> ), .C(n73), .Y(n67) );
  OAI21X1 U68 ( .A(n28), .B(n35), .C(n33), .Y(GG) );
  NAND3X1 U69 ( .A(n74), .B(n7), .C(n62), .Y(n63) );
  OAI21X1 U70 ( .A(n45), .B(n65), .C(n37), .Y(n66) );
  NAND2X1 U71 ( .A(n33), .B(n24), .Y(Cout) );
endmodule


module fulladder1_44 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_45 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_46 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_47 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_43 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_42 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_41 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_40 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_39 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_38 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_37 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_36 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_35 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_34 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_33 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module fulladder1_32 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module register16_0 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n35;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n19) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n20) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n21) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n22) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n23) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n24) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n25) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n26) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n27) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n28) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n29) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n30) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n31) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n32) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n33) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n34) );
  dff_15 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_14 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_13 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_12 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_11 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_10 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_9 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_8 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_7 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_6 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_5 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_4 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_3 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_2 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_1 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_0 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n34), .Y(n18) );
  INVX1 U5 ( .A(n33), .Y(n12) );
  INVX1 U6 ( .A(n32), .Y(n13) );
  INVX1 U7 ( .A(n31), .Y(n14) );
  INVX1 U8 ( .A(n30), .Y(n15) );
  INVX1 U9 ( .A(n29), .Y(n16) );
  INVX1 U10 ( .A(n28), .Y(n17) );
  INVX1 U11 ( .A(n27), .Y(n3) );
  INVX1 U12 ( .A(n26), .Y(n4) );
  INVX1 U13 ( .A(n25), .Y(n5) );
  INVX1 U14 ( .A(n24), .Y(n6) );
  INVX1 U15 ( .A(n23), .Y(n7) );
  INVX1 U16 ( .A(n22), .Y(n8) );
  INVX1 U17 ( .A(n21), .Y(n9) );
  INVX1 U34 ( .A(n20), .Y(n10) );
  INVX1 U35 ( .A(n19), .Y(n11) );
endmodule


module register16_1 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_31 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_30 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_29 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_28 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_27 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_26 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_25 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_24 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_23 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_22 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_21 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_20 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_19 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_18 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_17 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_16 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_2 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_47 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_46 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_45 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_44 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_43 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_42 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_41 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_40 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_39 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_38 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_37 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_36 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_35 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_34 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_33 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_32 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_3 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_63 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_62 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_61 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_60 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_59 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_58 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_57 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_56 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_55 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_54 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_53 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_52 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_51 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_50 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_49 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_48 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_4 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_79 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_78 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_77 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_76 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_75 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_74 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_73 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_72 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_71 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_70 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_69 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_68 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_67 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_66 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_65 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_64 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_5 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_95 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_94 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_93 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_92 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_91 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_90 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_89 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_88 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_87 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_86 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_85 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_84 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_83 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_82 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_81 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_80 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_6 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_111 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_110 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_109 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_108 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_107 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_106 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_105 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_104 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_103 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_102 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_101 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_100 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_99 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_98 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_97 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_96 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module register16_7 ( .d({\d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , 
        \d<9> , \d<8> , \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , 
        \d<0> }), clk, wr_en, rst, .q({\q<15> , \q<14> , \q<13> , \q<12> , 
        \q<11> , \q<10> , \q<9> , \q<8> , \q<7> , \q<6> , \q<5> , \q<4> , 
        \q<3> , \q<2> , \q<1> , \q<0> }) );
  input \d<15> , \d<14> , \d<13> , \d<12> , \d<11> , \d<10> , \d<9> , \d<8> ,
         \d<7> , \d<6> , \d<5> , \d<4> , \d<3> , \d<2> , \d<1> , \d<0> , clk,
         wr_en, rst;
  output \q<15> , \q<14> , \q<13> , \q<12> , \q<11> , \q<10> , \q<9> , \q<8> ,
         \q<7> , \q<6> , \q<5> , \q<4> , \q<3> , \q<2> , \q<1> , \q<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  AOI22X1 U18 ( .A(n1), .B(\d<9> ), .C(\q<9> ), .D(n35), .Y(n51) );
  AOI22X1 U19 ( .A(\d<8> ), .B(n1), .C(\q<8> ), .D(n35), .Y(n50) );
  AOI22X1 U20 ( .A(\d<7> ), .B(n1), .C(\q<7> ), .D(n35), .Y(n49) );
  AOI22X1 U21 ( .A(\d<6> ), .B(n1), .C(\q<6> ), .D(n35), .Y(n48) );
  AOI22X1 U22 ( .A(\d<5> ), .B(n1), .C(\q<5> ), .D(n35), .Y(n47) );
  AOI22X1 U23 ( .A(\d<4> ), .B(n1), .C(\q<4> ), .D(n35), .Y(n46) );
  AOI22X1 U24 ( .A(\d<3> ), .B(n1), .C(\q<3> ), .D(n35), .Y(n45) );
  AOI22X1 U25 ( .A(\d<2> ), .B(n1), .C(\q<2> ), .D(n35), .Y(n44) );
  AOI22X1 U26 ( .A(\d<1> ), .B(n2), .C(\q<1> ), .D(n35), .Y(n43) );
  AOI22X1 U27 ( .A(\d<15> ), .B(n2), .C(\q<15> ), .D(n35), .Y(n42) );
  AOI22X1 U28 ( .A(\d<14> ), .B(n2), .C(\q<14> ), .D(n35), .Y(n41) );
  AOI22X1 U29 ( .A(\d<13> ), .B(n2), .C(\q<13> ), .D(n35), .Y(n40) );
  AOI22X1 U30 ( .A(\d<12> ), .B(n2), .C(\q<12> ), .D(n35), .Y(n39) );
  AOI22X1 U31 ( .A(\d<11> ), .B(n2), .C(\q<11> ), .D(n35), .Y(n38) );
  AOI22X1 U32 ( .A(\d<10> ), .B(n2), .C(\q<10> ), .D(n35), .Y(n37) );
  AOI22X1 U33 ( .A(\d<0> ), .B(n2), .C(\q<0> ), .D(n35), .Y(n36) );
  dff_112 \dff_arr[0]  ( .q(\q<0> ), .d(n18), .clk(clk), .rst(rst) );
  dff_113 \dff_arr[1]  ( .q(\q<1> ), .d(n3), .clk(clk), .rst(rst) );
  dff_114 \dff_arr[2]  ( .q(\q<2> ), .d(n4), .clk(clk), .rst(rst) );
  dff_115 \dff_arr[3]  ( .q(\q<3> ), .d(n5), .clk(clk), .rst(rst) );
  dff_116 \dff_arr[4]  ( .q(\q<4> ), .d(n6), .clk(clk), .rst(rst) );
  dff_117 \dff_arr[5]  ( .q(\q<5> ), .d(n7), .clk(clk), .rst(rst) );
  dff_118 \dff_arr[6]  ( .q(\q<6> ), .d(n8), .clk(clk), .rst(rst) );
  dff_119 \dff_arr[7]  ( .q(\q<7> ), .d(n9), .clk(clk), .rst(rst) );
  dff_120 \dff_arr[8]  ( .q(\q<8> ), .d(n10), .clk(clk), .rst(rst) );
  dff_121 \dff_arr[9]  ( .q(\q<9> ), .d(n11), .clk(clk), .rst(rst) );
  dff_122 \dff_arr[10]  ( .q(\q<10> ), .d(n12), .clk(clk), .rst(rst) );
  dff_123 \dff_arr[11]  ( .q(\q<11> ), .d(n13), .clk(clk), .rst(rst) );
  dff_124 \dff_arr[12]  ( .q(\q<12> ), .d(n14), .clk(clk), .rst(rst) );
  dff_125 \dff_arr[13]  ( .q(\q<13> ), .d(n15), .clk(clk), .rst(rst) );
  dff_126 \dff_arr[14]  ( .q(\q<14> ), .d(n16), .clk(clk), .rst(rst) );
  dff_127 \dff_arr[15]  ( .q(\q<15> ), .d(n17), .clk(clk), .rst(rst) );
  BUFX2 U1 ( .A(wr_en), .Y(n1) );
  BUFX2 U2 ( .A(wr_en), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n35) );
  INVX1 U4 ( .A(n36), .Y(n18) );
  INVX1 U5 ( .A(n37), .Y(n12) );
  INVX1 U6 ( .A(n38), .Y(n13) );
  INVX1 U7 ( .A(n39), .Y(n14) );
  INVX1 U8 ( .A(n40), .Y(n15) );
  INVX1 U9 ( .A(n41), .Y(n16) );
  INVX1 U10 ( .A(n42), .Y(n17) );
  INVX1 U11 ( .A(n43), .Y(n3) );
  INVX1 U12 ( .A(n44), .Y(n4) );
  INVX1 U13 ( .A(n45), .Y(n5) );
  INVX1 U14 ( .A(n46), .Y(n6) );
  INVX1 U15 ( .A(n47), .Y(n7) );
  INVX1 U16 ( .A(n48), .Y(n8) );
  INVX1 U17 ( .A(n49), .Y(n9) );
  INVX1 U34 ( .A(n50), .Y(n10) );
  INVX1 U35 ( .A(n51), .Y(n11) );
endmodule


module decoder3to8 ( .In({\In<2> , \In<1> , \In<0> }), .Out({\Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<2> , \In<1> , \In<0> ;
  output \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> ,
         \Out<0> ;
  wire   n1, n2, n3;

  NOR3X1 U4 ( .A(n3), .B(n1), .C(n2), .Y(\Out<7> ) );
  NOR3X1 U5 ( .A(n3), .B(\In<0> ), .C(n2), .Y(\Out<6> ) );
  NOR3X1 U6 ( .A(n3), .B(\In<1> ), .C(n1), .Y(\Out<5> ) );
  NOR3X1 U7 ( .A(n3), .B(\In<1> ), .C(\In<0> ), .Y(\Out<4> ) );
  NOR3X1 U8 ( .A(n2), .B(\In<2> ), .C(n1), .Y(\Out<3> ) );
  NOR3X1 U9 ( .A(n2), .B(\In<2> ), .C(\In<0> ), .Y(\Out<2> ) );
  NOR3X1 U10 ( .A(n1), .B(\In<2> ), .C(\In<1> ), .Y(\Out<1> ) );
  NOR3X1 U11 ( .A(\In<0> ), .B(\In<2> ), .C(\In<1> ), .Y(\Out<0> ) );
  INVX1 U1 ( .A(\In<0> ), .Y(n1) );
  INVX1 U2 ( .A(\In<1> ), .Y(n2) );
  INVX1 U3 ( .A(\In<2> ), .Y(n3) );
endmodule


module mux8to1_16_1 ( .In({\In<127> , \In<126> , \In<125> , \In<124> , 
        \In<123> , \In<122> , \In<121> , \In<120> , \In<119> , \In<118> , 
        \In<117> , \In<116> , \In<115> , \In<114> , \In<113> , \In<112> , 
        \In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , 
        \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , 
        \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , 
        \In<78> , \In<77> , \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , 
        \In<71> , \In<70> , \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , 
        \In<64> , \In<63> , \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , 
        \In<57> , \In<56> , \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , 
        \In<50> , \In<49> , \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , 
        \In<43> , \In<42> , \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , 
        \In<36> , \In<35> , \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , 
        \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , 
        \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , 
        \In<0> }), .Sel({\Sel<2> , \Sel<1> , \Sel<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<127> , \In<126> , \In<125> , \In<124> , \In<123> , \In<122> ,
         \In<121> , \In<120> , \In<119> , \In<118> , \In<117> , \In<116> ,
         \In<115> , \In<114> , \In<113> , \In<112> , \In<111> , \In<110> ,
         \In<109> , \In<108> , \In<107> , \In<106> , \In<105> , \In<104> ,
         \In<103> , \In<102> , \In<101> , \In<100> , \In<99> , \In<98> ,
         \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , \In<92> , \In<91> ,
         \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , \In<85> , \In<84> ,
         \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , \In<78> , \In<77> ,
         \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , \In<71> , \In<70> ,
         \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , \In<64> , \In<63> ,
         \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , \In<57> , \In<56> ,
         \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , \In<50> , \In<49> ,
         \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> ,
         \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> ,
         \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , \In<29> , \In<28> ,
         \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , \In<22> , \In<21> ,
         \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , \In<15> , \In<14> ,
         \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , \In<8> , \In<7> ,
         \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , \In<0> ,
         \Sel<2> , \Sel<1> , \Sel<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \mux0_out<15> , \mux0_out<14> , \mux0_out<13> , \mux0_out<12> ,
         \mux0_out<11> , \mux0_out<10> , \mux0_out<9> , \mux0_out<8> ,
         \mux0_out<7> , \mux0_out<6> , \mux0_out<5> , \mux0_out<4> ,
         \mux0_out<3> , \mux0_out<2> , \mux0_out<1> , \mux0_out<0> ,
         \mux1_out<15> , \mux1_out<14> , \mux1_out<13> , \mux1_out<12> ,
         \mux1_out<11> , \mux1_out<10> , \mux1_out<9> , \mux1_out<8> ,
         \mux1_out<7> , \mux1_out<6> , \mux1_out<5> , \mux1_out<4> ,
         \mux1_out<3> , \mux1_out<2> , \mux1_out<1> , \mux1_out<0> , n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n35;

  AOI22X1 U18 ( .A(\mux0_out<9> ), .B(n18), .C(\mux1_out<9> ), .D(n35), .Y(n19) );
  AOI22X1 U19 ( .A(\mux0_out<8> ), .B(n18), .C(\mux1_out<8> ), .D(n35), .Y(n20) );
  AOI22X1 U20 ( .A(\mux0_out<7> ), .B(n18), .C(\mux1_out<7> ), .D(n35), .Y(n21) );
  AOI22X1 U21 ( .A(\mux0_out<6> ), .B(n18), .C(\mux1_out<6> ), .D(n35), .Y(n22) );
  AOI22X1 U22 ( .A(\mux0_out<5> ), .B(n18), .C(\mux1_out<5> ), .D(n35), .Y(n23) );
  AOI22X1 U23 ( .A(\mux0_out<4> ), .B(n18), .C(\mux1_out<4> ), .D(n35), .Y(n24) );
  AOI22X1 U24 ( .A(\mux0_out<3> ), .B(n18), .C(\mux1_out<3> ), .D(n35), .Y(n25) );
  AOI22X1 U25 ( .A(\mux0_out<2> ), .B(n18), .C(\mux1_out<2> ), .D(n35), .Y(n26) );
  AOI22X1 U26 ( .A(\mux0_out<1> ), .B(n18), .C(\mux1_out<1> ), .D(n35), .Y(n27) );
  AOI22X1 U27 ( .A(\mux0_out<15> ), .B(n18), .C(\mux1_out<15> ), .D(n35), .Y(
        n28) );
  AOI22X1 U28 ( .A(\mux0_out<14> ), .B(n18), .C(\mux1_out<14> ), .D(n35), .Y(
        n29) );
  AOI22X1 U29 ( .A(\mux0_out<13> ), .B(n18), .C(\mux1_out<13> ), .D(n35), .Y(
        n30) );
  AOI22X1 U30 ( .A(\mux0_out<12> ), .B(n18), .C(\mux1_out<12> ), .D(n17), .Y(
        n31) );
  AOI22X1 U31 ( .A(\mux0_out<11> ), .B(n18), .C(\mux1_out<11> ), .D(n17), .Y(
        n32) );
  AOI22X1 U32 ( .A(\mux0_out<10> ), .B(n18), .C(\mux1_out<10> ), .D(n35), .Y(
        n33) );
  AOI22X1 U33 ( .A(\mux0_out<0> ), .B(n18), .C(\mux1_out<0> ), .D(n17), .Y(n34) );
  mux4to1_16_3 mux0 ( .InA({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .InB({\In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> }), 
        .InC({\In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> , 
        \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> , 
        \In<34> , \In<33> , \In<32> }), .InD({\In<63> , \In<62> , \In<61> , 
        \In<60> , \In<59> , \In<58> , \In<57> , \In<56> , \In<55> , \In<54> , 
        \In<53> , \In<52> , \In<51> , \In<50> , \In<49> , \In<48> }), .S({
        \Sel<1> , \Sel<0> }), .Out({\mux0_out<15> , \mux0_out<14> , 
        \mux0_out<13> , \mux0_out<12> , \mux0_out<11> , \mux0_out<10> , 
        \mux0_out<9> , \mux0_out<8> , \mux0_out<7> , \mux0_out<6> , 
        \mux0_out<5> , \mux0_out<4> , \mux0_out<3> , \mux0_out<2> , 
        \mux0_out<1> , \mux0_out<0> }) );
  mux4to1_16_2 mux1 ( .InA({\In<79> , \In<78> , \In<77> , \In<76> , \In<75> , 
        \In<74> , \In<73> , \In<72> , \In<71> , \In<70> , \In<69> , \In<68> , 
        \In<67> , \In<66> , \In<65> , \In<64> }), .InB({\In<95> , \In<94> , 
        \In<93> , \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , 
        \In<86> , \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> }), 
        .InC({\In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> }), .InD({\In<127> , \In<126> , 
        \In<125> , \In<124> , \In<123> , \In<122> , \In<121> , \In<120> , 
        \In<119> , \In<118> , \In<117> , \In<116> , \In<115> , \In<114> , 
        \In<113> , \In<112> }), .S({\Sel<1> , \Sel<0> }), .Out({\mux1_out<15> , 
        \mux1_out<14> , \mux1_out<13> , \mux1_out<12> , \mux1_out<11> , 
        \mux1_out<10> , \mux1_out<9> , \mux1_out<8> , \mux1_out<7> , 
        \mux1_out<6> , \mux1_out<5> , \mux1_out<4> , \mux1_out<3> , 
        \mux1_out<2> , \mux1_out<1> , \mux1_out<0> }) );
  INVX1 U1 ( .A(\Sel<2> ), .Y(n18) );
  INVX1 U2 ( .A(n18), .Y(n35) );
  INVX1 U3 ( .A(n18), .Y(n17) );
  BUFX2 U4 ( .A(n34), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(\Out<0> ) );
  BUFX2 U6 ( .A(n33), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(\Out<10> ) );
  BUFX2 U8 ( .A(n32), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(\Out<11> ) );
  BUFX2 U10 ( .A(n31), .Y(n4) );
  INVX1 U11 ( .A(n4), .Y(\Out<12> ) );
  BUFX2 U12 ( .A(n30), .Y(n5) );
  INVX1 U13 ( .A(n5), .Y(\Out<13> ) );
  BUFX2 U14 ( .A(n29), .Y(n6) );
  INVX1 U15 ( .A(n6), .Y(\Out<14> ) );
  BUFX2 U16 ( .A(n28), .Y(n7) );
  INVX1 U17 ( .A(n7), .Y(\Out<15> ) );
  BUFX2 U34 ( .A(n27), .Y(n8) );
  INVX1 U35 ( .A(n8), .Y(\Out<1> ) );
  BUFX2 U36 ( .A(n26), .Y(n9) );
  INVX1 U37 ( .A(n9), .Y(\Out<2> ) );
  BUFX2 U38 ( .A(n25), .Y(n10) );
  INVX1 U39 ( .A(n10), .Y(\Out<3> ) );
  BUFX2 U40 ( .A(n24), .Y(n11) );
  INVX1 U41 ( .A(n11), .Y(\Out<4> ) );
  BUFX2 U42 ( .A(n23), .Y(n12) );
  INVX1 U43 ( .A(n12), .Y(\Out<5> ) );
  BUFX2 U44 ( .A(n22), .Y(n13) );
  INVX1 U45 ( .A(n13), .Y(\Out<6> ) );
  BUFX2 U46 ( .A(n21), .Y(n14) );
  INVX1 U47 ( .A(n14), .Y(\Out<7> ) );
  BUFX2 U48 ( .A(n20), .Y(n15) );
  INVX1 U49 ( .A(n15), .Y(\Out<8> ) );
  BUFX2 U50 ( .A(n19), .Y(n16) );
  INVX1 U51 ( .A(n16), .Y(\Out<9> ) );
endmodule


module mux8to1_16_0 ( .In({\In<127> , \In<126> , \In<125> , \In<124> , 
        \In<123> , \In<122> , \In<121> , \In<120> , \In<119> , \In<118> , 
        \In<117> , \In<116> , \In<115> , \In<114> , \In<113> , \In<112> , 
        \In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , 
        \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , 
        \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , 
        \In<78> , \In<77> , \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , 
        \In<71> , \In<70> , \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , 
        \In<64> , \In<63> , \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , 
        \In<57> , \In<56> , \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , 
        \In<50> , \In<49> , \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , 
        \In<43> , \In<42> , \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , 
        \In<36> , \In<35> , \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , 
        \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , 
        \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , 
        \In<0> }), .Sel({\Sel<2> , \Sel<1> , \Sel<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<127> , \In<126> , \In<125> , \In<124> , \In<123> , \In<122> ,
         \In<121> , \In<120> , \In<119> , \In<118> , \In<117> , \In<116> ,
         \In<115> , \In<114> , \In<113> , \In<112> , \In<111> , \In<110> ,
         \In<109> , \In<108> , \In<107> , \In<106> , \In<105> , \In<104> ,
         \In<103> , \In<102> , \In<101> , \In<100> , \In<99> , \In<98> ,
         \In<97> , \In<96> , \In<95> , \In<94> , \In<93> , \In<92> , \In<91> ,
         \In<90> , \In<89> , \In<88> , \In<87> , \In<86> , \In<85> , \In<84> ,
         \In<83> , \In<82> , \In<81> , \In<80> , \In<79> , \In<78> , \In<77> ,
         \In<76> , \In<75> , \In<74> , \In<73> , \In<72> , \In<71> , \In<70> ,
         \In<69> , \In<68> , \In<67> , \In<66> , \In<65> , \In<64> , \In<63> ,
         \In<62> , \In<61> , \In<60> , \In<59> , \In<58> , \In<57> , \In<56> ,
         \In<55> , \In<54> , \In<53> , \In<52> , \In<51> , \In<50> , \In<49> ,
         \In<48> , \In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> ,
         \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> ,
         \In<34> , \In<33> , \In<32> , \In<31> , \In<30> , \In<29> , \In<28> ,
         \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , \In<22> , \In<21> ,
         \In<20> , \In<19> , \In<18> , \In<17> , \In<16> , \In<15> , \In<14> ,
         \In<13> , \In<12> , \In<11> , \In<10> , \In<9> , \In<8> , \In<7> ,
         \In<6> , \In<5> , \In<4> , \In<3> , \In<2> , \In<1> , \In<0> ,
         \Sel<2> , \Sel<1> , \Sel<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \mux0_out<15> , \mux0_out<14> , \mux0_out<13> , \mux0_out<12> ,
         \mux0_out<11> , \mux0_out<10> , \mux0_out<9> , \mux0_out<8> ,
         \mux0_out<7> , \mux0_out<6> , \mux0_out<5> , \mux0_out<4> ,
         \mux0_out<3> , \mux0_out<2> , \mux0_out<1> , \mux0_out<0> ,
         \mux1_out<15> , \mux1_out<14> , \mux1_out<13> , \mux1_out<12> ,
         \mux1_out<11> , \mux1_out<10> , \mux1_out<9> , \mux1_out<8> ,
         \mux1_out<7> , \mux1_out<6> , \mux1_out<5> , \mux1_out<4> ,
         \mux1_out<3> , \mux1_out<2> , \mux1_out<1> , \mux1_out<0> , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n35, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67;

  AOI22X1 U18 ( .A(\mux0_out<9> ), .B(n18), .C(\mux1_out<9> ), .D(n35), .Y(n67) );
  AOI22X1 U19 ( .A(\mux0_out<8> ), .B(n18), .C(\mux1_out<8> ), .D(n35), .Y(n66) );
  AOI22X1 U20 ( .A(\mux0_out<7> ), .B(n18), .C(\mux1_out<7> ), .D(n35), .Y(n65) );
  AOI22X1 U21 ( .A(\mux0_out<6> ), .B(n18), .C(\mux1_out<6> ), .D(n35), .Y(n64) );
  AOI22X1 U22 ( .A(\mux0_out<5> ), .B(n18), .C(\mux1_out<5> ), .D(n35), .Y(n63) );
  AOI22X1 U23 ( .A(\mux0_out<4> ), .B(n18), .C(\mux1_out<4> ), .D(n35), .Y(n62) );
  AOI22X1 U24 ( .A(\mux0_out<3> ), .B(n18), .C(\mux1_out<3> ), .D(n35), .Y(n61) );
  AOI22X1 U25 ( .A(\mux0_out<2> ), .B(n18), .C(\mux1_out<2> ), .D(n35), .Y(n60) );
  AOI22X1 U26 ( .A(\mux0_out<1> ), .B(n18), .C(\mux1_out<1> ), .D(n35), .Y(n59) );
  AOI22X1 U27 ( .A(\mux0_out<15> ), .B(n18), .C(\mux1_out<15> ), .D(n35), .Y(
        n58) );
  AOI22X1 U28 ( .A(\mux0_out<14> ), .B(n18), .C(\mux1_out<14> ), .D(n35), .Y(
        n57) );
  AOI22X1 U29 ( .A(\mux0_out<13> ), .B(n18), .C(\mux1_out<13> ), .D(n35), .Y(
        n56) );
  AOI22X1 U30 ( .A(\mux0_out<12> ), .B(n18), .C(\mux1_out<12> ), .D(n17), .Y(
        n55) );
  AOI22X1 U31 ( .A(\mux0_out<11> ), .B(n18), .C(\mux1_out<11> ), .D(n17), .Y(
        n54) );
  AOI22X1 U32 ( .A(\mux0_out<10> ), .B(n18), .C(\mux1_out<10> ), .D(n35), .Y(
        n53) );
  AOI22X1 U33 ( .A(\mux0_out<0> ), .B(n18), .C(\mux1_out<0> ), .D(n17), .Y(n52) );
  mux4to1_16_1 mux0 ( .InA({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .InB({\In<31> , \In<30> , 
        \In<29> , \In<28> , \In<27> , \In<26> , \In<25> , \In<24> , \In<23> , 
        \In<22> , \In<21> , \In<20> , \In<19> , \In<18> , \In<17> , \In<16> }), 
        .InC({\In<47> , \In<46> , \In<45> , \In<44> , \In<43> , \In<42> , 
        \In<41> , \In<40> , \In<39> , \In<38> , \In<37> , \In<36> , \In<35> , 
        \In<34> , \In<33> , \In<32> }), .InD({\In<63> , \In<62> , \In<61> , 
        \In<60> , \In<59> , \In<58> , \In<57> , \In<56> , \In<55> , \In<54> , 
        \In<53> , \In<52> , \In<51> , \In<50> , \In<49> , \In<48> }), .S({
        \Sel<1> , \Sel<0> }), .Out({\mux0_out<15> , \mux0_out<14> , 
        \mux0_out<13> , \mux0_out<12> , \mux0_out<11> , \mux0_out<10> , 
        \mux0_out<9> , \mux0_out<8> , \mux0_out<7> , \mux0_out<6> , 
        \mux0_out<5> , \mux0_out<4> , \mux0_out<3> , \mux0_out<2> , 
        \mux0_out<1> , \mux0_out<0> }) );
  mux4to1_16_0 mux1 ( .InA({\In<79> , \In<78> , \In<77> , \In<76> , \In<75> , 
        \In<74> , \In<73> , \In<72> , \In<71> , \In<70> , \In<69> , \In<68> , 
        \In<67> , \In<66> , \In<65> , \In<64> }), .InB({\In<95> , \In<94> , 
        \In<93> , \In<92> , \In<91> , \In<90> , \In<89> , \In<88> , \In<87> , 
        \In<86> , \In<85> , \In<84> , \In<83> , \In<82> , \In<81> , \In<80> }), 
        .InC({\In<111> , \In<110> , \In<109> , \In<108> , \In<107> , \In<106> , 
        \In<105> , \In<104> , \In<103> , \In<102> , \In<101> , \In<100> , 
        \In<99> , \In<98> , \In<97> , \In<96> }), .InD({\In<127> , \In<126> , 
        \In<125> , \In<124> , \In<123> , \In<122> , \In<121> , \In<120> , 
        \In<119> , \In<118> , \In<117> , \In<116> , \In<115> , \In<114> , 
        \In<113> , \In<112> }), .S({\Sel<1> , \Sel<0> }), .Out({\mux1_out<15> , 
        \mux1_out<14> , \mux1_out<13> , \mux1_out<12> , \mux1_out<11> , 
        \mux1_out<10> , \mux1_out<9> , \mux1_out<8> , \mux1_out<7> , 
        \mux1_out<6> , \mux1_out<5> , \mux1_out<4> , \mux1_out<3> , 
        \mux1_out<2> , \mux1_out<1> , \mux1_out<0> }) );
  INVX1 U1 ( .A(\Sel<2> ), .Y(n18) );
  INVX1 U2 ( .A(n18), .Y(n35) );
  INVX1 U3 ( .A(n18), .Y(n17) );
  BUFX2 U4 ( .A(n52), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(\Out<0> ) );
  BUFX2 U6 ( .A(n53), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(\Out<10> ) );
  BUFX2 U8 ( .A(n54), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(\Out<11> ) );
  BUFX2 U10 ( .A(n55), .Y(n4) );
  INVX1 U11 ( .A(n4), .Y(\Out<12> ) );
  BUFX2 U12 ( .A(n56), .Y(n5) );
  INVX1 U13 ( .A(n5), .Y(\Out<13> ) );
  BUFX2 U14 ( .A(n57), .Y(n6) );
  INVX1 U15 ( .A(n6), .Y(\Out<14> ) );
  BUFX2 U16 ( .A(n58), .Y(n7) );
  INVX1 U17 ( .A(n7), .Y(\Out<15> ) );
  BUFX2 U34 ( .A(n59), .Y(n8) );
  INVX1 U35 ( .A(n8), .Y(\Out<1> ) );
  BUFX2 U36 ( .A(n60), .Y(n9) );
  INVX1 U37 ( .A(n9), .Y(\Out<2> ) );
  BUFX2 U38 ( .A(n61), .Y(n10) );
  INVX1 U39 ( .A(n10), .Y(\Out<3> ) );
  BUFX2 U40 ( .A(n62), .Y(n11) );
  INVX1 U41 ( .A(n11), .Y(\Out<4> ) );
  BUFX2 U42 ( .A(n63), .Y(n12) );
  INVX1 U43 ( .A(n12), .Y(\Out<5> ) );
  BUFX2 U44 ( .A(n64), .Y(n13) );
  INVX1 U45 ( .A(n13), .Y(\Out<6> ) );
  BUFX2 U46 ( .A(n65), .Y(n14) );
  INVX1 U47 ( .A(n14), .Y(\Out<7> ) );
  BUFX2 U48 ( .A(n66), .Y(n15) );
  INVX1 U49 ( .A(n15), .Y(\Out<8> ) );
  BUFX2 U50 ( .A(n67), .Y(n16) );
  INVX1 U51 ( .A(n16), .Y(\Out<9> ) );
endmodule


module demux1to8_16 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<2> , \S<1> , \S<0> }), 
    .Out0({\Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , 
        \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , 
        \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({
        \Out1<15> , \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , 
        \Out1<9> , \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , 
        \Out1<3> , \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , 
        \Out2<14> , \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , 
        \Out2<8> , \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , 
        \Out2<2> , \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , 
        \Out3<13> , \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , 
        \Out3<7> , \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , 
        \Out3<1> , \Out3<0> }), .Out4({\Out4<15> , \Out4<14> , \Out4<13> , 
        \Out4<12> , \Out4<11> , \Out4<10> , \Out4<9> , \Out4<8> , \Out4<7> , 
        \Out4<6> , \Out4<5> , \Out4<4> , \Out4<3> , \Out4<2> , \Out4<1> , 
        \Out4<0> }), .Out5({\Out5<15> , \Out5<14> , \Out5<13> , \Out5<12> , 
        \Out5<11> , \Out5<10> , \Out5<9> , \Out5<8> , \Out5<7> , \Out5<6> , 
        \Out5<5> , \Out5<4> , \Out5<3> , \Out5<2> , \Out5<1> , \Out5<0> }), 
    .Out6({\Out6<15> , \Out6<14> , \Out6<13> , \Out6<12> , \Out6<11> , 
        \Out6<10> , \Out6<9> , \Out6<8> , \Out6<7> , \Out6<6> , \Out6<5> , 
        \Out6<4> , \Out6<3> , \Out6<2> , \Out6<1> , \Out6<0> }), .Out7({
        \Out7<15> , \Out7<14> , \Out7<13> , \Out7<12> , \Out7<11> , \Out7<10> , 
        \Out7<9> , \Out7<8> , \Out7<7> , \Out7<6> , \Out7<5> , \Out7<4> , 
        \Out7<3> , \Out7<2> , \Out7<1> , \Out7<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<2> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> , \Out4<15> ,
         \Out4<14> , \Out4<13> , \Out4<12> , \Out4<11> , \Out4<10> , \Out4<9> ,
         \Out4<8> , \Out4<7> , \Out4<6> , \Out4<5> , \Out4<4> , \Out4<3> ,
         \Out4<2> , \Out4<1> , \Out4<0> , \Out5<15> , \Out5<14> , \Out5<13> ,
         \Out5<12> , \Out5<11> , \Out5<10> , \Out5<9> , \Out5<8> , \Out5<7> ,
         \Out5<6> , \Out5<5> , \Out5<4> , \Out5<3> , \Out5<2> , \Out5<1> ,
         \Out5<0> , \Out6<15> , \Out6<14> , \Out6<13> , \Out6<12> , \Out6<11> ,
         \Out6<10> , \Out6<9> , \Out6<8> , \Out6<7> , \Out6<6> , \Out6<5> ,
         \Out6<4> , \Out6<3> , \Out6<2> , \Out6<1> , \Out6<0> , \Out7<15> ,
         \Out7<14> , \Out7<13> , \Out7<12> , \Out7<11> , \Out7<10> , \Out7<9> ,
         \Out7<8> , \Out7<7> , \Out7<6> , \Out7<5> , \Out7<4> , \Out7<3> ,
         \Out7<2> , \Out7<1> , \Out7<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  demux1to8_0 \demux[0]  ( .In(\In<0> ), .S({n8, n3, \S<0> }), .Out0(\Out0<0> ), .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ), .Out4(\Out4<0> ), 
        .Out5(\Out5<0> ), .Out6(\Out6<0> ), .Out7(\Out7<0> ) );
  demux1to8_1 \demux[1]  ( .In(\In<1> ), .S({n9, n6, n4}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ), .Out4(\Out4<1> ), 
        .Out5(\Out5<1> ), .Out6(\Out6<1> ), .Out7(\Out7<1> ) );
  demux1to8_2 \demux[2]  ( .In(\In<2> ), .S({n9, n6, n4}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ), .Out4(\Out4<2> ), 
        .Out5(\Out5<2> ), .Out6(\Out6<2> ), .Out7(\Out7<2> ) );
  demux1to8_3 \demux[3]  ( .In(\In<3> ), .S({n9, n6, n4}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ), .Out4(\Out4<3> ), 
        .Out5(\Out5<3> ), .Out6(\Out6<3> ), .Out7(\Out7<3> ) );
  demux1to8_4 \demux[4]  ( .In(\In<4> ), .S({n9, n6, n4}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ), .Out4(\Out4<4> ), 
        .Out5(\Out5<4> ), .Out6(\Out6<4> ), .Out7(\Out7<4> ) );
  demux1to8_5 \demux[5]  ( .In(\In<5> ), .S({n8, n1, \S<0> }), .Out0(\Out0<5> ), .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ), .Out4(\Out4<5> ), 
        .Out5(\Out5<5> ), .Out6(\Out6<5> ), .Out7(\Out7<5> ) );
  demux1to8_6 \demux[6]  ( .In(\In<6> ), .S({n8, n2, \S<0> }), .Out0(\Out0<6> ), .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ), .Out4(\Out4<6> ), 
        .Out5(\Out5<6> ), .Out6(\Out6<6> ), .Out7(\Out7<6> ) );
  demux1to8_7 \demux[7]  ( .In(\In<7> ), .S({n8, n3, \S<0> }), .Out0(\Out0<7> ), .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ), .Out4(\Out4<7> ), 
        .Out5(\Out5<7> ), .Out6(\Out6<7> ), .Out7(\Out7<7> ) );
  demux1to8_8 \demux[8]  ( .In(\In<8> ), .S({n8, n1, \S<0> }), .Out0(\Out0<8> ), .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ), .Out4(\Out4<8> ), 
        .Out5(\Out5<8> ), .Out6(\Out6<8> ), .Out7(\Out7<8> ) );
  demux1to8_9 \demux[9]  ( .In(\In<9> ), .S({n8, n2, \S<0> }), .Out0(\Out0<9> ), .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ), .Out4(\Out4<9> ), 
        .Out5(\Out5<9> ), .Out6(\Out6<9> ), .Out7(\Out7<9> ) );
  demux1to8_10 \demux[10]  ( .In(\In<10> ), .S({n8, n3, \S<0> }), .Out0(
        \Out0<10> ), .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ), 
        .Out4(\Out4<10> ), .Out5(\Out5<10> ), .Out6(\Out6<10> ), .Out7(
        \Out7<10> ) );
  demux1to8_11 \demux[11]  ( .In(\In<11> ), .S({n8, n1, \S<0> }), .Out0(
        \Out0<11> ), .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ), 
        .Out4(\Out4<11> ), .Out5(\Out5<11> ), .Out6(\Out6<11> ), .Out7(
        \Out7<11> ) );
  demux1to8_12 \demux[12]  ( .In(\In<12> ), .S({n8, n2, \S<0> }), .Out0(
        \Out0<12> ), .Out1(\Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ), 
        .Out4(\Out4<12> ), .Out5(\Out5<12> ), .Out6(\Out6<12> ), .Out7(
        \Out7<12> ) );
  demux1to8_13 \demux[13]  ( .In(\In<13> ), .S({n8, n3, \S<0> }), .Out0(
        \Out0<13> ), .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ), 
        .Out4(\Out4<13> ), .Out5(\Out5<13> ), .Out6(\Out6<13> ), .Out7(
        \Out7<13> ) );
  demux1to8_14 \demux[14]  ( .In(\In<14> ), .S({n8, n1, \S<0> }), .Out0(
        \Out0<14> ), .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ), 
        .Out4(\Out4<14> ), .Out5(\Out5<14> ), .Out6(\Out6<14> ), .Out7(
        \Out7<14> ) );
  demux1to8_15 \demux[15]  ( .In(\In<15> ), .S({n8, n2, \S<0> }), .Out0(
        \Out0<15> ), .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ), 
        .Out4(\Out4<15> ), .Out5(\Out5<15> ), .Out6(\Out6<15> ), .Out7(
        \Out7<15> ) );
  INVX1 U1 ( .A(n7), .Y(n6) );
  INVX1 U2 ( .A(n7), .Y(n3) );
  INVX1 U3 ( .A(n7), .Y(n1) );
  INVX1 U4 ( .A(n7), .Y(n2) );
  INVX1 U5 ( .A(n5), .Y(n4) );
  INVX1 U6 ( .A(\S<2> ), .Y(n10) );
  INVX1 U7 ( .A(n10), .Y(n9) );
  INVX1 U8 ( .A(n10), .Y(n8) );
  INVX1 U9 ( .A(\S<0> ), .Y(n5) );
  INVX1 U10 ( .A(\S<1> ), .Y(n7) );
endmodule


module demux1to2_17 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_18 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2, n3;

  INVX1 U1 ( .A(S), .Y(n3) );
  INVX1 U2 ( .A(In), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U5 ( .A(n2), .B(n3), .Y(Out0) );
endmodule


module demux1to2_19 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_20 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_21 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_22 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X1 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_23 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_24 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_25 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_26 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_27 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_28 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_29 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_30 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_31 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_32 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_15 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  INVX1 U1 ( .A(S), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U3 ( .A(In), .B(n1), .Y(Out0) );
endmodule


module demux1to2_14 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(S), .Y(n2) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_13 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(In), .B(S), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_12 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  INVX1 U1 ( .A(S), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U3 ( .A(S), .B(In), .Y(Out1) );
  AND2X2 U4 ( .A(n1), .B(n2), .Y(Out0) );
endmodule


module demux1to2_11 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_10 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_9 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_8 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_7 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  INVX1 U1 ( .A(n1), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_6 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  BUFX2 U1 ( .A(In), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U4 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_5 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  AND2X2 U1 ( .A(In), .B(S), .Y(Out1) );
  INVX1 U2 ( .A(In), .Y(n1) );
endmodule


module demux1to2_4 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1, n2;

  NOR2X1 U3 ( .A(S), .B(n2), .Y(Out0) );
  INVX1 U1 ( .A(n1), .Y(n2) );
  BUFX2 U2 ( .A(In), .Y(n1) );
  AND2X2 U4 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_3 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_2 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X1 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to2_1 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(S), .B(In), .Y(Out1) );
endmodule


module demux1to2_0 ( In, S, Out0, Out1 );
  input In, S;
  output Out0, Out1;
  wire   n1;

  NOR2X1 U3 ( .A(S), .B(n1), .Y(Out0) );
  INVX1 U1 ( .A(In), .Y(n1) );
  AND2X2 U2 ( .A(In), .B(S), .Y(Out1) );
endmodule


module demux1to4_16_1 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<1> , \S<0> }), .Out0({
        \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , 
        \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , 
        \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , 
        \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , 
        \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , 
        \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , \Out2<14> , 
        \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , 
        \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , 
        \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , \Out3<13> , 
        \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , 
        \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , 
        \Out3<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> ;
  wire   n11, n12, n3, n4, n5, n6, n7, n8, n9, n10;

  demux1to4_17 \demux[0]  ( .In(\In<0> ), .S({n5, n3}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ) );
  demux1to4_18 \demux[1]  ( .In(\In<1> ), .S({n7, n8}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ) );
  demux1to4_19 \demux[2]  ( .In(\In<2> ), .S({n7, n4}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ) );
  demux1to4_20 \demux[3]  ( .In(\In<3> ), .S({n5, n3}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ) );
  demux1to4_21 \demux[4]  ( .In(\In<4> ), .S({n6, n4}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ) );
  demux1to4_22 \demux[5]  ( .In(\In<5> ), .S({n5, n3}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ) );
  demux1to4_23 \demux[6]  ( .In(\In<6> ), .S({n5, n3}), .Out0(\Out0<6> ), 
        .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ) );
  demux1to4_24 \demux[7]  ( .In(\In<7> ), .S({n7, n8}), .Out0(n12), .Out1(
        \Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ) );
  demux1to4_25 \demux[8]  ( .In(\In<8> ), .S({n7, n3}), .Out0(\Out0<8> ), 
        .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ) );
  demux1to4_26 \demux[9]  ( .In(\In<9> ), .S({n6, n4}), .Out0(\Out0<9> ), 
        .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ) );
  demux1to4_27 \demux[10]  ( .In(\In<10> ), .S({n7, n3}), .Out0(n11), .Out1(
        \Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ) );
  demux1to4_28 \demux[11]  ( .In(\In<11> ), .S({n6, n4}), .Out0(\Out0<11> ), 
        .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ) );
  demux1to4_29 \demux[12]  ( .In(\In<12> ), .S({n6, n4}), .Out0(\Out0<12> ), 
        .Out1(\Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ) );
  demux1to4_30 \demux[13]  ( .In(\In<13> ), .S({n6, n4}), .Out0(\Out0<13> ), 
        .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ) );
  demux1to4_31 \demux[14]  ( .In(\In<14> ), .S({n7, n8}), .Out0(\Out0<14> ), 
        .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ) );
  demux1to4_32 \demux[15]  ( .In(\In<15> ), .S({n6, n4}), .Out0(\Out0<15> ), 
        .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ) );
  INVX2 U1 ( .A(n9), .Y(n8) );
  BUFX4 U2 ( .A(n11), .Y(\Out0<10> ) );
  BUFX2 U3 ( .A(n12), .Y(\Out0<7> ) );
  INVX4 U4 ( .A(\S<0> ), .Y(n9) );
  INVX4 U5 ( .A(n10), .Y(n6) );
  INVX8 U6 ( .A(n9), .Y(n3) );
  INVX8 U7 ( .A(n9), .Y(n4) );
  INVX8 U8 ( .A(n10), .Y(n5) );
  INVX8 U9 ( .A(n10), .Y(n7) );
  INVX8 U10 ( .A(\S<1> ), .Y(n10) );
endmodule


module demux1to4_16_0 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .S({\S<1> , \S<0> }), .Out0({
        \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , 
        \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , 
        \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , 
        \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , 
        \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , 
        \Out1<2> , \Out1<1> , \Out1<0> }), .Out2({\Out2<15> , \Out2<14> , 
        \Out2<13> , \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , 
        \Out2<7> , \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , 
        \Out2<1> , \Out2<0> }), .Out3({\Out3<15> , \Out3<14> , \Out3<13> , 
        \Out3<12> , \Out3<11> , \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , 
        \Out3<6> , \Out3<5> , \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , 
        \Out3<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \S<1> , \S<0> ;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> , \Out2<15> , \Out2<14> , \Out2<13> ,
         \Out2<12> , \Out2<11> , \Out2<10> , \Out2<9> , \Out2<8> , \Out2<7> ,
         \Out2<6> , \Out2<5> , \Out2<4> , \Out2<3> , \Out2<2> , \Out2<1> ,
         \Out2<0> , \Out3<15> , \Out3<14> , \Out3<13> , \Out3<12> , \Out3<11> ,
         \Out3<10> , \Out3<9> , \Out3<8> , \Out3<7> , \Out3<6> , \Out3<5> ,
         \Out3<4> , \Out3<3> , \Out3<2> , \Out3<1> , \Out3<0> ;
  wire   n9, n2, n3, n4, n5, n6, n7, n8;

  demux1to4_15 \demux[0]  ( .In(\In<0> ), .S({n7, n3}), .Out0(\Out0<0> ), 
        .Out1(\Out1<0> ), .Out2(\Out2<0> ), .Out3(\Out3<0> ) );
  demux1to4_14 \demux[1]  ( .In(\In<1> ), .S({n7, n3}), .Out0(\Out0<1> ), 
        .Out1(\Out1<1> ), .Out2(\Out2<1> ), .Out3(\Out3<1> ) );
  demux1to4_13 \demux[2]  ( .In(\In<2> ), .S({n7, n4}), .Out0(\Out0<2> ), 
        .Out1(\Out1<2> ), .Out2(\Out2<2> ), .Out3(\Out3<2> ) );
  demux1to4_12 \demux[3]  ( .In(\In<3> ), .S({n7, n3}), .Out0(\Out0<3> ), 
        .Out1(\Out1<3> ), .Out2(\Out2<3> ), .Out3(\Out3<3> ) );
  demux1to4_11 \demux[4]  ( .In(\In<4> ), .S({n7, n4}), .Out0(\Out0<4> ), 
        .Out1(\Out1<4> ), .Out2(\Out2<4> ), .Out3(\Out3<4> ) );
  demux1to4_10 \demux[5]  ( .In(\In<5> ), .S({n7, n3}), .Out0(\Out0<5> ), 
        .Out1(\Out1<5> ), .Out2(\Out2<5> ), .Out3(\Out3<5> ) );
  demux1to4_9 \demux[6]  ( .In(\In<6> ), .S({n7, n4}), .Out0(\Out0<6> ), 
        .Out1(\Out1<6> ), .Out2(\Out2<6> ), .Out3(\Out3<6> ) );
  demux1to4_8 \demux[7]  ( .In(\In<7> ), .S({n7, n3}), .Out0(\Out0<7> ), 
        .Out1(\Out1<7> ), .Out2(\Out2<7> ), .Out3(\Out3<7> ) );
  demux1to4_7 \demux[8]  ( .In(\In<8> ), .S({n7, n4}), .Out0(\Out0<8> ), 
        .Out1(\Out1<8> ), .Out2(\Out2<8> ), .Out3(\Out3<8> ) );
  demux1to4_6 \demux[9]  ( .In(\In<9> ), .S({n7, n5}), .Out0(\Out0<9> ), 
        .Out1(\Out1<9> ), .Out2(\Out2<9> ), .Out3(\Out3<9> ) );
  demux1to4_5 \demux[10]  ( .In(\In<10> ), .S({n7, n3}), .Out0(\Out0<10> ), 
        .Out1(\Out1<10> ), .Out2(\Out2<10> ), .Out3(\Out3<10> ) );
  demux1to4_4 \demux[11]  ( .In(\In<11> ), .S({n7, n3}), .Out0(\Out0<11> ), 
        .Out1(\Out1<11> ), .Out2(\Out2<11> ), .Out3(\Out3<11> ) );
  demux1to4_3 \demux[12]  ( .In(\In<12> ), .S({n7, n4}), .Out0(n9), .Out1(
        \Out1<12> ), .Out2(\Out2<12> ), .Out3(\Out3<12> ) );
  demux1to4_2 \demux[13]  ( .In(\In<13> ), .S({n7, n4}), .Out0(\Out0<13> ), 
        .Out1(\Out1<13> ), .Out2(\Out2<13> ), .Out3(\Out3<13> ) );
  demux1to4_1 \demux[14]  ( .In(\In<14> ), .S({n7, n3}), .Out0(\Out0<14> ), 
        .Out1(\Out1<14> ), .Out2(\Out2<14> ), .Out3(\Out3<14> ) );
  demux1to4_0 \demux[15]  ( .In(\In<15> ), .S({n7, n3}), .Out0(\Out0<15> ), 
        .Out1(\Out1<15> ), .Out2(\Out2<15> ), .Out3(\Out3<15> ) );
  INVX2 U1 ( .A(n5), .Y(n2) );
  BUFX2 U2 ( .A(n9), .Y(\Out0<12> ) );
  INVX1 U3 ( .A(\S<0> ), .Y(n6) );
  INVX1 U4 ( .A(n6), .Y(n5) );
  INVX1 U5 ( .A(\S<1> ), .Y(n8) );
  INVX8 U6 ( .A(n2), .Y(n3) );
  INVX8 U7 ( .A(n2), .Y(n4) );
  INVX8 U8 ( .A(n8), .Y(n7) );
endmodule


module cla16_0 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n1,
         n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22;

  cla4_3 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_2 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n2), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_1 ca2 ( .A({\A<11> , \A<10> , \A<9> , n15}), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n22), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_0 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n8), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  INVX1 U1 ( .A(n7), .Y(n8) );
  INVX2 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(\G<3> ), .Y(n21) );
  AND2X2 U4 ( .A(n19), .B(n20), .Y(n1) );
  AND2X2 U5 ( .A(n21), .B(n12), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(Cout) );
  BUFX2 U7 ( .A(n18), .Y(n5) );
  BUFX2 U8 ( .A(n17), .Y(n6) );
  AND2X2 U9 ( .A(n5), .B(n6), .Y(n7) );
  INVX1 U10 ( .A(n7), .Y(n9) );
  BUFX2 U11 ( .A(\G<0> ), .Y(n10) );
  AND2X2 U12 ( .A(\P<3> ), .B(n9), .Y(n11) );
  INVX1 U13 ( .A(n11), .Y(n12) );
  AOI21X1 U14 ( .A(Cin), .B(\P<0> ), .C(n10), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(n16) );
  AOI21X1 U16 ( .A(\P<1> ), .B(n16), .C(\G<1> ), .Y(n14) );
  INVX1 U17 ( .A(n14), .Y(n22) );
  BUFX4 U18 ( .A(\A<8> ), .Y(n15) );
  INVX1 U19 ( .A(n10), .Y(n20) );
  AOI21X1 U20 ( .A(\G<1> ), .B(\P<2> ), .C(\G<2> ), .Y(n18) );
  NAND2X1 U21 ( .A(Cin), .B(\P<0> ), .Y(n19) );
  NAND3X1 U22 ( .A(\P<1> ), .B(\P<2> ), .C(n16), .Y(n17) );
endmodule


module mux4to1_16_4 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n150, n151, n1, n2, n3, n5, n7, n9, n10, n12, n13, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n97, n100, n101, n103, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146;

  INVX1 U1 ( .A(\InC<11> ), .Y(n133) );
  INVX1 U2 ( .A(\InD<10> ), .Y(n129) );
  AND2X1 U3 ( .A(\InA<2> ), .B(n112), .Y(n19) );
  OR2X1 U4 ( .A(\InA<11> ), .B(n134), .Y(n25) );
  INVX1 U5 ( .A(\InC<13> ), .Y(n139) );
  INVX1 U6 ( .A(n1), .Y(\Out<12> ) );
  AND2X1 U7 ( .A(\InA<7> ), .B(n112), .Y(n21) );
  AND2X1 U8 ( .A(\InA<5> ), .B(n112), .Y(n23) );
  OAI21X1 U9 ( .A(n137), .B(\InA<12> ), .C(n84), .Y(n1) );
  INVX1 U10 ( .A(\InA<14> ), .Y(n141) );
  AND2X2 U11 ( .A(n115), .B(n116), .Y(n2) );
  AND2X1 U12 ( .A(\InA<8> ), .B(n112), .Y(n15) );
  AND2X2 U13 ( .A(n70), .B(n9), .Y(n3) );
  INVX1 U14 ( .A(n3), .Y(\Out<1> ) );
  AND2X2 U15 ( .A(n35), .B(n22), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(\Out<7> ) );
  AND2X2 U17 ( .A(n36), .B(n20), .Y(n7) );
  INVX1 U18 ( .A(n7), .Y(\Out<2> ) );
  AND2X2 U19 ( .A(n67), .B(n18), .Y(n9) );
  AND2X2 U20 ( .A(n24), .B(n37), .Y(n10) );
  INVX1 U21 ( .A(n10), .Y(\Out<5> ) );
  AND2X1 U22 ( .A(\InA<4> ), .B(n112), .Y(n12) );
  OR2X2 U23 ( .A(n26), .B(n81), .Y(n13) );
  INVX1 U24 ( .A(n13), .Y(\Out<11> ) );
  INVX1 U25 ( .A(n15), .Y(n16) );
  AND2X1 U26 ( .A(\InA<1> ), .B(n112), .Y(n17) );
  INVX1 U27 ( .A(n17), .Y(n18) );
  INVX1 U28 ( .A(n19), .Y(n20) );
  INVX1 U29 ( .A(n21), .Y(n22) );
  INVX1 U30 ( .A(n23), .Y(n24) );
  INVX1 U31 ( .A(n25), .Y(n26) );
  AND2X1 U32 ( .A(\InA<3> ), .B(n112), .Y(n27) );
  INVX1 U33 ( .A(n27), .Y(n28) );
  AND2X1 U34 ( .A(\InA<6> ), .B(n112), .Y(n29) );
  INVX1 U35 ( .A(n29), .Y(n30) );
  AND2X1 U36 ( .A(n114), .B(n116), .Y(n31) );
  AND2X1 U37 ( .A(n114), .B(n117), .Y(n32) );
  OR2X1 U38 ( .A(n100), .B(n34), .Y(\Out<0> ) );
  OR2X1 U39 ( .A(n43), .B(n42), .Y(n34) );
  AND2X1 U40 ( .A(n79), .B(n64), .Y(n35) );
  AND2X1 U41 ( .A(n72), .B(n61), .Y(n36) );
  AND2X1 U42 ( .A(n77), .B(n63), .Y(n37) );
  AND2X2 U43 ( .A(n75), .B(n40), .Y(n38) );
  INVX1 U44 ( .A(n38), .Y(\Out<4> ) );
  AND2X1 U45 ( .A(n74), .B(n62), .Y(n40) );
  AND2X1 U46 ( .A(n68), .B(n66), .Y(n41) );
  AND2X1 U47 ( .A(\InA<0> ), .B(n112), .Y(n42) );
  AND2X1 U48 ( .A(\InB<0> ), .B(n32), .Y(n43) );
  AND2X1 U49 ( .A(\InD<9> ), .B(n31), .Y(n44) );
  INVX1 U50 ( .A(n44), .Y(n45) );
  AND2X1 U51 ( .A(\InD<14> ), .B(n31), .Y(n46) );
  INVX1 U52 ( .A(n46), .Y(n47) );
  AND2X1 U53 ( .A(\InD<15> ), .B(n31), .Y(n48) );
  INVX1 U54 ( .A(n48), .Y(n49) );
  AND2X1 U55 ( .A(\InB<9> ), .B(n32), .Y(n50) );
  INVX1 U56 ( .A(n50), .Y(n51) );
  AND2X1 U57 ( .A(\InB<14> ), .B(n32), .Y(n52) );
  INVX1 U58 ( .A(n52), .Y(n53) );
  AND2X1 U59 ( .A(\InB<15> ), .B(n32), .Y(n54) );
  INVX1 U60 ( .A(n54), .Y(n55) );
  BUFX2 U61 ( .A(n132), .Y(n56) );
  BUFX2 U62 ( .A(n135), .Y(n57) );
  BUFX2 U63 ( .A(n138), .Y(n58) );
  AND2X1 U64 ( .A(\InB<10> ), .B(n32), .Y(n59) );
  INVX1 U65 ( .A(n59), .Y(n60) );
  BUFX2 U66 ( .A(n120), .Y(n61) );
  BUFX2 U67 ( .A(n122), .Y(n62) );
  BUFX2 U68 ( .A(n123), .Y(n63) );
  BUFX2 U69 ( .A(n125), .Y(n64) );
  AND2X1 U70 ( .A(\InC<8> ), .B(n2), .Y(n65) );
  INVX1 U71 ( .A(n65), .Y(n66) );
  BUFX2 U72 ( .A(n119), .Y(n67) );
  BUFX2 U73 ( .A(n126), .Y(n68) );
  AND2X1 U74 ( .A(\InB<1> ), .B(n32), .Y(n69) );
  INVX1 U75 ( .A(n69), .Y(n70) );
  AND2X1 U76 ( .A(\InC<2> ), .B(n2), .Y(n71) );
  INVX1 U77 ( .A(n71), .Y(n72) );
  AND2X1 U78 ( .A(\InC<4> ), .B(n2), .Y(n73) );
  INVX1 U79 ( .A(n73), .Y(n74) );
  INVX1 U80 ( .A(n12), .Y(n75) );
  AND2X1 U81 ( .A(\InC<5> ), .B(n2), .Y(n76) );
  INVX1 U82 ( .A(n76), .Y(n77) );
  AND2X1 U83 ( .A(\InC<7> ), .B(n2), .Y(n78) );
  INVX1 U84 ( .A(n78), .Y(n79) );
  OR2X1 U85 ( .A(n134), .B(n112), .Y(n80) );
  INVX1 U86 ( .A(n80), .Y(n81) );
  AND2X2 U87 ( .A(n45), .B(n51), .Y(n82) );
  INVX1 U88 ( .A(n82), .Y(n83) );
  OR2X1 U89 ( .A(n137), .B(n112), .Y(n84) );
  AND2X2 U90 ( .A(n47), .B(n53), .Y(n85) );
  INVX1 U91 ( .A(n85), .Y(n86) );
  AND2X2 U92 ( .A(n49), .B(n55), .Y(n87) );
  INVX1 U93 ( .A(n87), .Y(n88) );
  BUFX2 U94 ( .A(n121), .Y(n89) );
  BUFX2 U95 ( .A(n124), .Y(n90) );
  AND2X2 U96 ( .A(\InB<3> ), .B(n32), .Y(n91) );
  INVX1 U97 ( .A(n91), .Y(n92) );
  AND2X1 U98 ( .A(\InB<6> ), .B(n32), .Y(n93) );
  INVX1 U99 ( .A(n93), .Y(n94) );
  INVX1 U100 ( .A(n146), .Y(n95) );
  INVX1 U101 ( .A(n95), .Y(\Out<9> ) );
  AND2X2 U102 ( .A(n16), .B(n41), .Y(n97) );
  INVX1 U103 ( .A(n97), .Y(\Out<8> ) );
  INVX1 U104 ( .A(n118), .Y(n100) );
  INVX1 U105 ( .A(n151), .Y(n101) );
  INVX1 U106 ( .A(n101), .Y(\Out<3> ) );
  INVX1 U107 ( .A(n150), .Y(n103) );
  INVX1 U108 ( .A(n103), .Y(\Out<6> ) );
  BUFX2 U109 ( .A(n144), .Y(n105) );
  BUFX2 U110 ( .A(n128), .Y(n106) );
  BUFX2 U111 ( .A(n142), .Y(n107) );
  INVX1 U112 ( .A(n31), .Y(n108) );
  INVX1 U113 ( .A(n115), .Y(n114) );
  INVX1 U114 ( .A(\S<0> ), .Y(n115) );
  INVX1 U115 ( .A(n2), .Y(n109) );
  INVX1 U116 ( .A(n117), .Y(n116) );
  AOI21X1 U117 ( .A(\InA<10> ), .B(n112), .C(n110), .Y(n111) );
  INVX1 U118 ( .A(n131), .Y(n110) );
  INVX1 U119 ( .A(n111), .Y(\Out<10> ) );
  AOI21X1 U120 ( .A(n112), .B(\InA<13> ), .C(n140), .Y(n113) );
  INVX1 U121 ( .A(n145), .Y(n112) );
  INVX1 U122 ( .A(n113), .Y(\Out<13> ) );
  INVX1 U123 ( .A(\S<1> ), .Y(n117) );
  INVX1 U124 ( .A(\InA<9> ), .Y(n127) );
  INVX1 U125 ( .A(\InA<15> ), .Y(n143) );
  AOI22X1 U126 ( .A(\InD<0> ), .B(n31), .C(\InC<0> ), .D(n2), .Y(n118) );
  OR2X2 U127 ( .A(n116), .B(n114), .Y(n145) );
  AOI22X1 U128 ( .A(\InD<1> ), .B(n31), .C(\InC<1> ), .D(n2), .Y(n119) );
  AOI22X1 U129 ( .A(\InD<2> ), .B(n31), .C(\InB<2> ), .D(n32), .Y(n120) );
  AOI22X1 U130 ( .A(\InD<3> ), .B(n31), .C(\InC<3> ), .D(n2), .Y(n121) );
  NAND3X1 U131 ( .A(n28), .B(n89), .C(n92), .Y(n151) );
  AOI22X1 U132 ( .A(\InD<4> ), .B(n31), .C(\InB<4> ), .D(n32), .Y(n122) );
  AOI22X1 U133 ( .A(\InB<5> ), .B(n32), .C(\InD<5> ), .D(n31), .Y(n123) );
  AOI22X1 U134 ( .A(\InD<6> ), .B(n31), .C(\InC<6> ), .D(n2), .Y(n124) );
  NAND3X1 U135 ( .A(n30), .B(n90), .C(n94), .Y(n150) );
  AOI22X1 U136 ( .A(\InD<7> ), .B(n31), .C(\InB<7> ), .D(n32), .Y(n125) );
  AOI22X1 U137 ( .A(\InD<8> ), .B(n31), .C(\InB<8> ), .D(n32), .Y(n126) );
  AOI21X1 U138 ( .A(\InC<9> ), .B(n2), .C(n83), .Y(n128) );
  AOI22X1 U139 ( .A(n145), .B(n106), .C(n127), .D(n106), .Y(n146) );
  OAI21X1 U140 ( .A(n108), .B(n129), .C(n60), .Y(n130) );
  AOI21X1 U141 ( .A(\InC<10> ), .B(n2), .C(n130), .Y(n131) );
  AOI22X1 U142 ( .A(\InD<11> ), .B(n31), .C(\InB<11> ), .D(n32), .Y(n132) );
  OAI21X1 U143 ( .A(n109), .B(n133), .C(n56), .Y(n134) );
  INVX2 U144 ( .A(\InC<12> ), .Y(n136) );
  AOI22X1 U145 ( .A(\InD<12> ), .B(n31), .C(\InB<12> ), .D(n32), .Y(n135) );
  OAI21X1 U146 ( .A(n109), .B(n136), .C(n57), .Y(n137) );
  AOI22X1 U147 ( .A(\InD<13> ), .B(n31), .C(\InB<13> ), .D(n32), .Y(n138) );
  OAI21X1 U148 ( .A(n109), .B(n139), .C(n58), .Y(n140) );
  AOI21X1 U149 ( .A(\InC<14> ), .B(n2), .C(n86), .Y(n142) );
  AOI22X1 U150 ( .A(n145), .B(n107), .C(n107), .D(n141), .Y(\Out<14> ) );
  AOI21X1 U151 ( .A(\InC<15> ), .B(n2), .C(n88), .Y(n144) );
  AOI22X1 U152 ( .A(n145), .B(n105), .C(n105), .D(n143), .Y(\Out<15> ) );
endmodule


module lshifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), Rot_sel, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , Rot_sel;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n127, n129, n131, n133, n135, n137, n139, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277;

  INVX4 U2 ( .A(n173), .Y(n174) );
  INVX1 U3 ( .A(\In<13> ), .Y(n213) );
  INVX1 U4 ( .A(\In<14> ), .Y(n225) );
  INVX1 U5 ( .A(\In<10> ), .Y(n217) );
  INVX1 U6 ( .A(\In<1> ), .Y(n204) );
  INVX1 U7 ( .A(\Cnt<0> ), .Y(n202) );
  INVX1 U8 ( .A(\Cnt<2> ), .Y(n207) );
  INVX1 U9 ( .A(\Cnt<3> ), .Y(n201) );
  INVX1 U10 ( .A(\In<12> ), .Y(n244) );
  INVX1 U11 ( .A(\In<11> ), .Y(n229) );
  AND2X1 U12 ( .A(n85), .B(n95), .Y(n135) );
  INVX1 U13 ( .A(\In<0> ), .Y(n211) );
  INVX4 U14 ( .A(n32), .Y(n33) );
  AND2X2 U15 ( .A(\In<9> ), .B(n32), .Y(n59) );
  AND2X2 U16 ( .A(n202), .B(\Cnt<1> ), .Y(n171) );
  OR2X2 U17 ( .A(n8), .B(n2), .Y(n1) );
  OR2X2 U18 ( .A(n179), .B(n61), .Y(n2) );
  OR2X2 U19 ( .A(n6), .B(n4), .Y(n3) );
  OR2X2 U20 ( .A(n192), .B(n59), .Y(n4) );
  AND2X2 U21 ( .A(n63), .B(n12), .Y(n5) );
  AND2X2 U22 ( .A(\In<10> ), .B(n254), .Y(n6) );
  AND2X2 U23 ( .A(\Cnt<0> ), .B(n212), .Y(n7) );
  AND2X2 U24 ( .A(\In<6> ), .B(n254), .Y(n8) );
  AND2X2 U25 ( .A(\In<14> ), .B(n254), .Y(n9) );
  INVX1 U26 ( .A(n9), .Y(n10) );
  AND2X2 U27 ( .A(\In<0> ), .B(n7), .Y(n11) );
  INVX1 U28 ( .A(n11), .Y(n12) );
  BUFX2 U29 ( .A(n216), .Y(n13) );
  BUFX2 U30 ( .A(n263), .Y(n14) );
  BUFX2 U31 ( .A(n265), .Y(n15) );
  BUFX2 U32 ( .A(n277), .Y(n16) );
  BUFX2 U33 ( .A(n262), .Y(n17) );
  BUFX2 U34 ( .A(n264), .Y(n18) );
  BUFX2 U35 ( .A(n270), .Y(n19) );
  BUFX2 U36 ( .A(n218), .Y(n20) );
  BUFX2 U37 ( .A(n223), .Y(n21) );
  BUFX2 U38 ( .A(n236), .Y(n22) );
  AND2X2 U39 ( .A(Rot_sel), .B(n214), .Y(n23) );
  INVX1 U40 ( .A(n23), .Y(n24) );
  AND2X2 U41 ( .A(Rot_sel), .B(n226), .Y(n25) );
  INVX1 U42 ( .A(n25), .Y(n26) );
  BUFX2 U43 ( .A(n239), .Y(n27) );
  AND2X2 U44 ( .A(\In<15> ), .B(n254), .Y(n28) );
  INVX1 U45 ( .A(n28), .Y(n29) );
  AND2X2 U46 ( .A(n166), .B(n185), .Y(n30) );
  INVX1 U47 ( .A(n30), .Y(n31) );
  AND2X2 U48 ( .A(\Cnt<0> ), .B(\Cnt<1> ), .Y(n32) );
  AND2X2 U49 ( .A(\Cnt<3> ), .B(\Cnt<2> ), .Y(n34) );
  INVX1 U50 ( .A(n215), .Y(n35) );
  INVX1 U51 ( .A(n35), .Y(n36) );
  OR2X1 U52 ( .A(n33), .B(n204), .Y(n37) );
  INVX1 U53 ( .A(n37), .Y(n38) );
  OR2X1 U54 ( .A(n33), .B(n217), .Y(n39) );
  INVX1 U55 ( .A(n39), .Y(n40) );
  OR2X1 U56 ( .A(n33), .B(n240), .Y(n41) );
  INVX1 U57 ( .A(n41), .Y(n42) );
  OR2X1 U58 ( .A(n33), .B(n222), .Y(n43) );
  INVX1 U59 ( .A(n43), .Y(n44) );
  OR2X1 U60 ( .A(n33), .B(n229), .Y(n45) );
  INVX1 U61 ( .A(n45), .Y(n46) );
  OR2X1 U62 ( .A(n33), .B(n232), .Y(n47) );
  INVX1 U63 ( .A(n47), .Y(n48) );
  OR2X1 U64 ( .A(n33), .B(n235), .Y(n49) );
  INVX1 U65 ( .A(n49), .Y(n50) );
  OR2X1 U66 ( .A(n33), .B(n244), .Y(n51) );
  INVX1 U67 ( .A(n51), .Y(n52) );
  OR2X1 U68 ( .A(n33), .B(n247), .Y(n53) );
  INVX1 U69 ( .A(n53), .Y(n54) );
  OR2X1 U70 ( .A(n33), .B(n250), .Y(n55) );
  INVX1 U71 ( .A(n55), .Y(n56) );
  OR2X1 U72 ( .A(n33), .B(n211), .Y(n57) );
  INVX1 U73 ( .A(n57), .Y(n58) );
  AND2X2 U74 ( .A(Rot_sel), .B(n168), .Y(n60) );
  AND2X1 U75 ( .A(\In<5> ), .B(n208), .Y(n61) );
  INVX1 U76 ( .A(n33), .Y(n208) );
  AND2X2 U77 ( .A(\In<1> ), .B(n253), .Y(n62) );
  INVX1 U78 ( .A(n62), .Y(n63) );
  AND2X2 U79 ( .A(n167), .B(n1), .Y(n64) );
  INVX1 U80 ( .A(n64), .Y(n65) );
  BUFX2 U81 ( .A(n206), .Y(n66) );
  INVX1 U82 ( .A(n219), .Y(n67) );
  INVX1 U83 ( .A(n67), .Y(n68) );
  BUFX2 U84 ( .A(n221), .Y(n69) );
  INVX1 U85 ( .A(n228), .Y(n70) );
  INVX1 U86 ( .A(n70), .Y(n71) );
  INVX1 U87 ( .A(n224), .Y(n72) );
  INVX1 U88 ( .A(n72), .Y(n73) );
  BUFX2 U89 ( .A(n231), .Y(n74) );
  BUFX2 U90 ( .A(n234), .Y(n75) );
  BUFX2 U91 ( .A(n243), .Y(n76) );
  INVX1 U92 ( .A(n237), .Y(n77) );
  INVX1 U93 ( .A(n77), .Y(n78) );
  BUFX2 U94 ( .A(n246), .Y(n79) );
  BUFX2 U95 ( .A(n249), .Y(n80) );
  INVX1 U96 ( .A(n258), .Y(n81) );
  INVX1 U97 ( .A(n81), .Y(n82) );
  BUFX2 U98 ( .A(n252), .Y(n83) );
  BUFX2 U99 ( .A(n256), .Y(n84) );
  BUFX2 U100 ( .A(n269), .Y(n85) );
  INVX1 U101 ( .A(n271), .Y(n86) );
  INVX1 U102 ( .A(n86), .Y(n87) );
  AND2X2 U103 ( .A(n212), .B(n238), .Y(n88) );
  INVX1 U104 ( .A(n88), .Y(n89) );
  BUFX2 U105 ( .A(n227), .Y(n90) );
  BUFX2 U106 ( .A(n242), .Y(n91) );
  INVX1 U107 ( .A(n257), .Y(n92) );
  INVX1 U108 ( .A(n92), .Y(n93) );
  INVX1 U109 ( .A(n268), .Y(n94) );
  INVX1 U110 ( .A(n94), .Y(n95) );
  INVX1 U111 ( .A(n276), .Y(n96) );
  INVX1 U112 ( .A(n96), .Y(n97) );
  INVX1 U113 ( .A(n205), .Y(n98) );
  INVX1 U114 ( .A(n98), .Y(n99) );
  INVX1 U115 ( .A(n220), .Y(n100) );
  INVX1 U116 ( .A(n100), .Y(n101) );
  INVX1 U117 ( .A(n230), .Y(n102) );
  INVX1 U118 ( .A(n102), .Y(n103) );
  INVX1 U119 ( .A(n233), .Y(n104) );
  INVX1 U120 ( .A(n104), .Y(n105) );
  INVX1 U121 ( .A(n245), .Y(n106) );
  INVX1 U122 ( .A(n106), .Y(n107) );
  BUFX2 U123 ( .A(n248), .Y(n108) );
  BUFX2 U124 ( .A(n251), .Y(n109) );
  INVX1 U125 ( .A(n255), .Y(n110) );
  INVX1 U126 ( .A(n110), .Y(n111) );
  AND2X2 U127 ( .A(n167), .B(n181), .Y(n112) );
  INVX1 U128 ( .A(n112), .Y(n113) );
  AND2X2 U129 ( .A(n167), .B(n183), .Y(n114) );
  INVX1 U130 ( .A(n114), .Y(n115) );
  AND2X1 U131 ( .A(n168), .B(n174), .Y(n116) );
  INVX1 U132 ( .A(n116), .Y(n117) );
  AND2X1 U133 ( .A(n168), .B(n273), .Y(n118) );
  INVX1 U134 ( .A(n118), .Y(n119) );
  AND2X1 U135 ( .A(n34), .B(n174), .Y(n120) );
  INVX1 U136 ( .A(n120), .Y(n121) );
  AND2X1 U137 ( .A(n34), .B(n273), .Y(n122) );
  INVX1 U138 ( .A(n122), .Y(n123) );
  AND2X1 U139 ( .A(Rot_sel), .B(n166), .Y(n124) );
  AND2X2 U140 ( .A(n13), .B(n36), .Y(n125) );
  INVX1 U141 ( .A(n125), .Y(\Out<0> ) );
  AND2X2 U142 ( .A(n71), .B(n90), .Y(n127) );
  INVX1 U143 ( .A(n127), .Y(\Out<1> ) );
  AND2X2 U144 ( .A(n82), .B(n93), .Y(n129) );
  INVX1 U145 ( .A(n129), .Y(\Out<3> ) );
  AND2X2 U146 ( .A(n14), .B(n17), .Y(n131) );
  INVX1 U147 ( .A(n131), .Y(\Out<7> ) );
  AND2X2 U148 ( .A(n15), .B(n18), .Y(n133) );
  INVX1 U149 ( .A(n133), .Y(\Out<8> ) );
  INVX1 U150 ( .A(n135), .Y(\Out<11> ) );
  AND2X2 U151 ( .A(n87), .B(n19), .Y(n137) );
  INVX1 U152 ( .A(n137), .Y(\Out<12> ) );
  AND2X2 U153 ( .A(n16), .B(n97), .Y(n139) );
  INVX1 U154 ( .A(n139), .Y(\Out<15> ) );
  AND2X2 U155 ( .A(\In<15> ), .B(Rot_sel), .Y(n141) );
  INVX1 U156 ( .A(n141), .Y(n142) );
  AND2X2 U157 ( .A(n166), .B(n174), .Y(n143) );
  INVX1 U158 ( .A(n143), .Y(n144) );
  AND2X1 U159 ( .A(n166), .B(n273), .Y(n145) );
  INVX1 U160 ( .A(n145), .Y(n146) );
  AND2X1 U161 ( .A(n167), .B(n176), .Y(n147) );
  INVX1 U162 ( .A(n147), .Y(n148) );
  AND2X1 U163 ( .A(n167), .B(n178), .Y(n149) );
  INVX1 U164 ( .A(n149), .Y(n150) );
  AND2X2 U165 ( .A(n168), .B(n187), .Y(n151) );
  INVX1 U166 ( .A(n151), .Y(n152) );
  AND2X1 U167 ( .A(n168), .B(n189), .Y(n153) );
  INVX1 U168 ( .A(n153), .Y(n154) );
  INVX1 U169 ( .A(n259), .Y(n155) );
  INVX1 U170 ( .A(n155), .Y(n156) );
  INVX1 U171 ( .A(n260), .Y(n157) );
  INVX1 U172 ( .A(n157), .Y(n158) );
  INVX1 U173 ( .A(n261), .Y(n159) );
  INVX1 U174 ( .A(n159), .Y(n160) );
  BUFX2 U175 ( .A(n266), .Y(n161) );
  BUFX2 U176 ( .A(n267), .Y(n162) );
  INVX1 U177 ( .A(n272), .Y(n163) );
  INVX1 U178 ( .A(n163), .Y(n164) );
  BUFX2 U179 ( .A(n274), .Y(n165) );
  AND2X1 U180 ( .A(n201), .B(\Cnt<2> ), .Y(n166) );
  AND2X1 U181 ( .A(Rot_sel), .B(n34), .Y(n167) );
  AND2X1 U182 ( .A(\Cnt<3> ), .B(n207), .Y(n168) );
  AND2X2 U183 ( .A(n76), .B(n91), .Y(n169) );
  INVX1 U184 ( .A(n169), .Y(\Out<2> ) );
  INVX1 U185 ( .A(n171), .Y(n172) );
  AND2X2 U186 ( .A(n5), .B(n26), .Y(n173) );
  AND2X2 U187 ( .A(n68), .B(n20), .Y(n175) );
  INVX1 U188 ( .A(n175), .Y(n176) );
  AND2X2 U189 ( .A(n74), .B(n103), .Y(n177) );
  INVX1 U190 ( .A(n177), .Y(n178) );
  INVX1 U191 ( .A(n209), .Y(n179) );
  AND2X2 U192 ( .A(n73), .B(n21), .Y(n180) );
  INVX1 U193 ( .A(n180), .Y(n181) );
  AND2X2 U194 ( .A(n78), .B(n22), .Y(n182) );
  INVX1 U195 ( .A(n182), .Y(n183) );
  AND2X2 U196 ( .A(n89), .B(n24), .Y(n184) );
  INVX1 U197 ( .A(n184), .Y(n185) );
  AND2X2 U198 ( .A(n69), .B(n101), .Y(n186) );
  INVX1 U199 ( .A(n186), .Y(n187) );
  AND2X2 U200 ( .A(n75), .B(n105), .Y(n188) );
  INVX1 U201 ( .A(n188), .Y(n189) );
  AND2X2 U202 ( .A(n79), .B(n107), .Y(n190) );
  INVX1 U203 ( .A(n190), .Y(n191) );
  INVX1 U204 ( .A(n203), .Y(n192) );
  AND2X2 U205 ( .A(n83), .B(n109), .Y(n193) );
  INVX1 U206 ( .A(n193), .Y(n194) );
  AND2X2 U207 ( .A(n66), .B(n99), .Y(n195) );
  INVX1 U208 ( .A(n195), .Y(n196) );
  AND2X2 U209 ( .A(n80), .B(n108), .Y(n197) );
  INVX1 U210 ( .A(n197), .Y(n198) );
  AND2X2 U211 ( .A(n84), .B(n111), .Y(n199) );
  INVX1 U212 ( .A(n199), .Y(n200) );
  INVX1 U213 ( .A(\Cnt<1> ), .Y(n212) );
  INVX4 U214 ( .A(n172), .Y(n254) );
  INVX8 U215 ( .A(n241), .Y(n253) );
  INVX8 U216 ( .A(n210), .Y(n275) );
  OR2X2 U217 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n241) );
  AOI22X1 U218 ( .A(\In<11> ), .B(n7), .C(\In<12> ), .D(n253), .Y(n203) );
  AOI22X1 U219 ( .A(\In<4> ), .B(n253), .C(\In<3> ), .D(n7), .Y(n206) );
  AOI21X1 U220 ( .A(\In<2> ), .B(n254), .C(n38), .Y(n205) );
  AOI22X1 U221 ( .A(n124), .B(n3), .C(n167), .D(n196), .Y(n216) );
  AOI22X1 U222 ( .A(\In<7> ), .B(n7), .C(\In<8> ), .D(n253), .Y(n209) );
  OR2X2 U223 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n210) );
  MUX2X1 U224 ( .B(n211), .A(n142), .S(\Cnt<0> ), .Y(n238) );
  OAI21X1 U225 ( .A(n33), .B(n213), .C(n10), .Y(n214) );
  AOI22X1 U226 ( .A(n60), .B(n1), .C(n275), .D(n185), .Y(n215) );
  AOI22X1 U227 ( .A(\In<13> ), .B(n253), .C(\In<12> ), .D(n7), .Y(n219) );
  AOI21X1 U228 ( .A(\In<11> ), .B(n254), .C(n40), .Y(n218) );
  AOI22X1 U229 ( .A(\In<5> ), .B(n253), .C(\In<4> ), .D(n7), .Y(n221) );
  INVX2 U230 ( .A(\In<2> ), .Y(n240) );
  AOI21X1 U231 ( .A(\In<3> ), .B(n254), .C(n42), .Y(n220) );
  AOI22X1 U232 ( .A(n124), .B(n176), .C(n167), .D(n187), .Y(n228) );
  AOI22X1 U233 ( .A(\In<9> ), .B(n253), .C(\In<8> ), .D(n7), .Y(n224) );
  INVX2 U234 ( .A(\In<6> ), .Y(n222) );
  AOI21X1 U235 ( .A(\In<7> ), .B(n254), .C(n44), .Y(n223) );
  OAI21X1 U236 ( .A(n33), .B(n225), .C(n29), .Y(n226) );
  AOI22X1 U237 ( .A(n60), .B(n181), .C(n275), .D(n174), .Y(n227) );
  AOI22X1 U238 ( .A(\In<14> ), .B(n253), .C(\In<13> ), .D(n7), .Y(n231) );
  AOI21X1 U239 ( .A(\In<12> ), .B(n254), .C(n46), .Y(n230) );
  AOI22X1 U240 ( .A(\In<6> ), .B(n253), .C(\In<5> ), .D(n7), .Y(n234) );
  INVX2 U241 ( .A(\In<3> ), .Y(n232) );
  AOI21X1 U242 ( .A(\In<4> ), .B(n254), .C(n48), .Y(n233) );
  AOI22X1 U243 ( .A(n124), .B(n178), .C(n167), .D(n189), .Y(n243) );
  AOI22X1 U244 ( .A(\In<10> ), .B(n253), .C(\In<9> ), .D(n7), .Y(n237) );
  INVX2 U245 ( .A(\In<7> ), .Y(n235) );
  AOI21X1 U246 ( .A(\In<8> ), .B(n254), .C(n50), .Y(n236) );
  AOI22X1 U247 ( .A(\In<1> ), .B(n7), .C(\Cnt<1> ), .D(n238), .Y(n239) );
  OAI21X1 U248 ( .A(n241), .B(n240), .C(n27), .Y(n273) );
  AOI22X1 U249 ( .A(n60), .B(n183), .C(n275), .D(n273), .Y(n242) );
  AOI22X1 U250 ( .A(\In<15> ), .B(n253), .C(\In<14> ), .D(n7), .Y(n246) );
  AOI21X1 U251 ( .A(\In<13> ), .B(n254), .C(n52), .Y(n245) );
  AOI22X1 U252 ( .A(\In<7> ), .B(n253), .C(\In<6> ), .D(n7), .Y(n249) );
  INVX2 U253 ( .A(\In<4> ), .Y(n247) );
  AOI21X1 U254 ( .A(\In<5> ), .B(n254), .C(n54), .Y(n248) );
  AOI22X1 U255 ( .A(n124), .B(n191), .C(n167), .D(n198), .Y(n258) );
  AOI22X1 U256 ( .A(\In<11> ), .B(n253), .C(\In<10> ), .D(n7), .Y(n252) );
  INVX2 U257 ( .A(\In<8> ), .Y(n250) );
  AOI21X1 U258 ( .A(\In<9> ), .B(n254), .C(n56), .Y(n251) );
  AOI22X1 U259 ( .A(\In<3> ), .B(n253), .C(\In<2> ), .D(n7), .Y(n256) );
  AOI21X1 U260 ( .A(\In<1> ), .B(n254), .C(n58), .Y(n255) );
  AOI22X1 U261 ( .A(n60), .B(n194), .C(n275), .D(n200), .Y(n257) );
  AOI22X1 U262 ( .A(n3), .B(n60), .C(n196), .D(n275), .Y(n259) );
  NAND3X1 U263 ( .A(n65), .B(n31), .C(n156), .Y(\Out<4> ) );
  AOI22X1 U264 ( .A(n60), .B(n176), .C(n275), .D(n187), .Y(n260) );
  NAND3X1 U265 ( .A(n113), .B(n144), .C(n158), .Y(\Out<5> ) );
  AOI22X1 U266 ( .A(n60), .B(n178), .C(n275), .D(n189), .Y(n261) );
  NAND3X1 U267 ( .A(n115), .B(n146), .C(n160), .Y(\Out<6> ) );
  AOI22X1 U268 ( .A(n166), .B(n200), .C(n167), .D(n194), .Y(n263) );
  AOI22X1 U269 ( .A(n60), .B(n191), .C(n275), .D(n198), .Y(n262) );
  AOI22X1 U270 ( .A(n167), .B(n3), .C(n185), .D(n168), .Y(n265) );
  AOI22X1 U271 ( .A(n275), .B(n1), .C(n196), .D(n166), .Y(n264) );
  AOI22X1 U272 ( .A(n275), .B(n181), .C(n166), .D(n187), .Y(n266) );
  NAND3X1 U273 ( .A(n117), .B(n148), .C(n161), .Y(\Out<9> ) );
  AOI22X1 U274 ( .A(n275), .B(n183), .C(n166), .D(n189), .Y(n267) );
  NAND3X1 U275 ( .A(n119), .B(n150), .C(n162), .Y(\Out<10> ) );
  AOI22X1 U276 ( .A(n167), .B(n191), .C(n168), .D(n200), .Y(n269) );
  AOI22X1 U277 ( .A(n275), .B(n194), .C(n166), .D(n198), .Y(n268) );
  AOI22X1 U278 ( .A(n196), .B(n168), .C(n34), .D(n185), .Y(n271) );
  AOI22X1 U279 ( .A(n3), .B(n275), .C(n166), .D(n1), .Y(n270) );
  AOI22X1 U280 ( .A(n275), .B(n176), .C(n166), .D(n181), .Y(n272) );
  NAND3X1 U281 ( .A(n121), .B(n152), .C(n164), .Y(\Out<13> ) );
  AOI22X1 U282 ( .A(n275), .B(n178), .C(n166), .D(n183), .Y(n274) );
  NAND3X1 U283 ( .A(n123), .B(n154), .C(n165), .Y(\Out<14> ) );
  AOI22X1 U284 ( .A(n168), .B(n198), .C(n34), .D(n200), .Y(n277) );
  AOI22X1 U285 ( .A(n275), .B(n191), .C(n166), .D(n194), .Y(n276) );
endmodule


module rshifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), Rot_sel, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> })
 );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , Rot_sel;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n140, n142, n144, n146, n147, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281;

  INVX1 U2 ( .A(\In<7> ), .Y(n212) );
  INVX1 U3 ( .A(\In<3> ), .Y(n216) );
  INVX1 U4 ( .A(\In<4> ), .Y(n230) );
  INVX1 U5 ( .A(\Cnt<0> ), .Y(n204) );
  INVX1 U6 ( .A(\In<6> ), .Y(n258) );
  INVX1 U7 ( .A(\In<8> ), .Y(n227) );
  INVX1 U8 ( .A(\Cnt<2> ), .Y(n203) );
  INVX1 U9 ( .A(\Cnt<3> ), .Y(n211) );
  INVX1 U10 ( .A(\In<15> ), .Y(n208) );
  INVX1 U11 ( .A(\In<9> ), .Y(n240) );
  INVX1 U12 ( .A(\In<12> ), .Y(n224) );
  INVX1 U13 ( .A(n248), .Y(n222) );
  INVX1 U14 ( .A(Rot_sel), .Y(n202) );
  AND2X1 U15 ( .A(n29), .B(n85), .Y(n138) );
  INVX4 U16 ( .A(n169), .Y(n170) );
  INVX1 U17 ( .A(n175), .Y(n1) );
  AND2X2 U18 ( .A(n181), .B(n174), .Y(n135) );
  AND2X2 U19 ( .A(n280), .B(n181), .Y(n129) );
  AND2X2 U20 ( .A(n171), .B(n181), .Y(n61) );
  OR2X2 U21 ( .A(n170), .B(n230), .Y(n113) );
  OR2X2 U22 ( .A(n170), .B(n216), .Y(n107) );
  OR2X2 U23 ( .A(n170), .B(n224), .Y(n109) );
  OR2X2 U24 ( .A(n170), .B(n227), .Y(n111) );
  OR2X2 U25 ( .A(n170), .B(n243), .Y(n119) );
  OR2X2 U26 ( .A(n170), .B(n240), .Y(n117) );
  OR2X2 U27 ( .A(n170), .B(n237), .Y(n115) );
  OR2X2 U28 ( .A(n170), .B(n247), .Y(n121) );
  INVX1 U29 ( .A(n170), .Y(n205) );
  OR2X2 U30 ( .A(n170), .B(n251), .Y(n123) );
  AND2X2 U31 ( .A(n204), .B(\Cnt<1> ), .Y(n175) );
  AND2X2 U32 ( .A(\Cnt<0> ), .B(\Cnt<1> ), .Y(n169) );
  OR2X2 U33 ( .A(n60), .B(n3), .Y(\Out<3> ) );
  OR2X2 U34 ( .A(n137), .B(n61), .Y(n3) );
  OR2X2 U35 ( .A(n52), .B(n5), .Y(n4) );
  OR2X2 U36 ( .A(n53), .B(n11), .Y(n5) );
  OR2X2 U37 ( .A(n56), .B(n7), .Y(n6) );
  OR2X2 U38 ( .A(n57), .B(n14), .Y(n7) );
  OR2X2 U39 ( .A(n41), .B(n9), .Y(n8) );
  OR2X2 U40 ( .A(n182), .B(n10), .Y(n9) );
  AND2X2 U41 ( .A(\In<11> ), .B(n205), .Y(n10) );
  AND2X2 U42 ( .A(\Cnt<1> ), .B(n222), .Y(n11) );
  AND2X2 U43 ( .A(n40), .B(n4), .Y(n12) );
  INVX1 U44 ( .A(n12), .Y(n13) );
  AND2X2 U45 ( .A(n201), .B(n235), .Y(n14) );
  AND2X2 U46 ( .A(n40), .B(n6), .Y(n15) );
  INVX1 U47 ( .A(n15), .Y(n16) );
  OR2X2 U48 ( .A(n170), .B(n254), .Y(n17) );
  INVX1 U49 ( .A(n17), .Y(n18) );
  OR2X2 U50 ( .A(n170), .B(n258), .Y(n19) );
  INVX1 U51 ( .A(n19), .Y(n20) );
  AND2X1 U52 ( .A(n184), .B(n174), .Y(n21) );
  INVX1 U53 ( .A(n21), .Y(n22) );
  AND2X2 U54 ( .A(n102), .B(n100), .Y(n23) );
  INVX1 U55 ( .A(n23), .Y(\Out<5> ) );
  AND2X2 U56 ( .A(n173), .B(n6), .Y(n25) );
  INVX1 U57 ( .A(n25), .Y(n26) );
  AND2X2 U58 ( .A(n280), .B(n6), .Y(n27) );
  INVX1 U59 ( .A(n27), .Y(n28) );
  BUFX2 U60 ( .A(n220), .Y(n29) );
  BUFX2 U61 ( .A(n266), .Y(n30) );
  BUFX2 U62 ( .A(n270), .Y(n31) );
  BUFX2 U63 ( .A(n275), .Y(n32) );
  BUFX2 U64 ( .A(n225), .Y(n33) );
  BUFX2 U65 ( .A(n228), .Y(n34) );
  BUFX2 U66 ( .A(n238), .Y(n35) );
  BUFX2 U67 ( .A(n252), .Y(n36) );
  BUFX2 U68 ( .A(n255), .Y(n37) );
  BUFX2 U69 ( .A(n250), .Y(n38) );
  BUFX2 U70 ( .A(n263), .Y(n39) );
  AND2X1 U71 ( .A(\Cnt<3> ), .B(\Cnt<2> ), .Y(n40) );
  AND2X2 U72 ( .A(\In<10> ), .B(n259), .Y(n41) );
  AND2X1 U73 ( .A(n8), .B(n173), .Y(n42) );
  INVX1 U74 ( .A(n42), .Y(n43) );
  INVX1 U75 ( .A(n268), .Y(n44) );
  INVX1 U76 ( .A(n44), .Y(n45) );
  INVX1 U77 ( .A(n241), .Y(n46) );
  INVX1 U78 ( .A(n46), .Y(n47) );
  INVX1 U79 ( .A(n233), .Y(n48) );
  INVX1 U80 ( .A(n48), .Y(n49) );
  INVX1 U81 ( .A(n246), .Y(n50) );
  INVX1 U82 ( .A(n50), .Y(n51) );
  AND2X2 U83 ( .A(\In<14> ), .B(n172), .Y(n52) );
  AND2X1 U84 ( .A(\In<13> ), .B(n223), .Y(n53) );
  INVX1 U85 ( .A(n236), .Y(n223) );
  AND2X1 U86 ( .A(n171), .B(n177), .Y(n54) );
  INVX1 U87 ( .A(n54), .Y(n55) );
  AND2X1 U88 ( .A(\In<15> ), .B(n172), .Y(n56) );
  AND2X1 U89 ( .A(\In<14> ), .B(n223), .Y(n57) );
  AND2X1 U90 ( .A(n171), .B(n179), .Y(n58) );
  INVX1 U91 ( .A(n58), .Y(n59) );
  AND2X1 U92 ( .A(n40), .B(n279), .Y(n60) );
  AND2X2 U93 ( .A(n201), .B(n171), .Y(n62) );
  BUFX2 U94 ( .A(n210), .Y(n63) );
  BUFX2 U95 ( .A(n214), .Y(n64) );
  BUFX2 U96 ( .A(n218), .Y(n65) );
  BUFX2 U97 ( .A(n226), .Y(n66) );
  BUFX2 U98 ( .A(n229), .Y(n67) );
  BUFX2 U99 ( .A(n232), .Y(n68) );
  BUFX2 U100 ( .A(n239), .Y(n69) );
  BUFX2 U101 ( .A(n242), .Y(n70) );
  BUFX2 U102 ( .A(n245), .Y(n71) );
  BUFX2 U103 ( .A(n253), .Y(n72) );
  INVX1 U104 ( .A(n256), .Y(n73) );
  INVX1 U105 ( .A(n73), .Y(n74) );
  BUFX2 U106 ( .A(n261), .Y(n75) );
  INVX1 U107 ( .A(n267), .Y(n76) );
  INVX1 U108 ( .A(n76), .Y(n77) );
  INVX1 U109 ( .A(n269), .Y(n78) );
  INVX1 U110 ( .A(n78), .Y(n79) );
  INVX1 U111 ( .A(n271), .Y(n80) );
  INVX1 U112 ( .A(n80), .Y(n81) );
  INVX1 U113 ( .A(n276), .Y(n82) );
  INVX1 U114 ( .A(n82), .Y(n83) );
  INVX1 U115 ( .A(n219), .Y(n84) );
  INVX1 U116 ( .A(n84), .Y(n85) );
  INVX1 U117 ( .A(n209), .Y(n86) );
  INVX1 U118 ( .A(n86), .Y(n87) );
  INVX1 U119 ( .A(n213), .Y(n88) );
  INVX1 U120 ( .A(n88), .Y(n89) );
  INVX1 U121 ( .A(n217), .Y(n90) );
  INVX1 U122 ( .A(n90), .Y(n91) );
  INVX1 U123 ( .A(n231), .Y(n92) );
  INVX1 U124 ( .A(n92), .Y(n93) );
  INVX1 U125 ( .A(n244), .Y(n94) );
  INVX1 U126 ( .A(n94), .Y(n95) );
  INVX1 U127 ( .A(n260), .Y(n96) );
  INVX1 U128 ( .A(n96), .Y(n97) );
  AND2X2 U129 ( .A(\In<0> ), .B(n175), .Y(n98) );
  INVX1 U130 ( .A(n98), .Y(n99) );
  BUFX2 U131 ( .A(n264), .Y(n100) );
  INVX1 U132 ( .A(n265), .Y(n101) );
  INVX1 U133 ( .A(n101), .Y(n102) );
  OR2X2 U134 ( .A(n170), .B(n208), .Y(n103) );
  INVX1 U135 ( .A(n103), .Y(n104) );
  OR2X2 U136 ( .A(n170), .B(n212), .Y(n105) );
  INVX1 U137 ( .A(n105), .Y(n106) );
  INVX1 U138 ( .A(n107), .Y(n108) );
  INVX1 U139 ( .A(n109), .Y(n110) );
  INVX1 U140 ( .A(n111), .Y(n112) );
  INVX1 U141 ( .A(n113), .Y(n114) );
  INVX1 U142 ( .A(n115), .Y(n116) );
  INVX1 U143 ( .A(n117), .Y(n118) );
  INVX1 U144 ( .A(n119), .Y(n120) );
  INVX1 U145 ( .A(n121), .Y(n122) );
  INVX1 U146 ( .A(n123), .Y(n124) );
  AND2X2 U147 ( .A(n280), .B(n177), .Y(n125) );
  INVX1 U148 ( .A(n125), .Y(n126) );
  AND2X1 U149 ( .A(n280), .B(n179), .Y(n127) );
  INVX1 U150 ( .A(n127), .Y(n128) );
  INVX1 U151 ( .A(n129), .Y(n130) );
  AND2X1 U152 ( .A(n177), .B(n174), .Y(n131) );
  INVX1 U153 ( .A(n131), .Y(n132) );
  AND2X1 U154 ( .A(n179), .B(n174), .Y(n133) );
  INVX1 U155 ( .A(n133), .Y(n134) );
  INVX1 U156 ( .A(n135), .Y(n136) );
  INVX1 U157 ( .A(n262), .Y(n137) );
  INVX1 U158 ( .A(n138), .Y(\Out<0> ) );
  AND2X2 U159 ( .A(n77), .B(n30), .Y(n140) );
  INVX1 U160 ( .A(n140), .Y(\Out<6> ) );
  AND2X2 U161 ( .A(n79), .B(n45), .Y(n142) );
  INVX1 U162 ( .A(n142), .Y(\Out<7> ) );
  AND2X2 U163 ( .A(n81), .B(n31), .Y(n144) );
  INVX1 U164 ( .A(n144), .Y(\Out<8> ) );
  AND2X1 U165 ( .A(n201), .B(n173), .Y(n146) );
  AND2X2 U166 ( .A(n83), .B(n32), .Y(n147) );
  INVX1 U167 ( .A(n147), .Y(\Out<12> ) );
  AND2X2 U168 ( .A(n173), .B(n4), .Y(n149) );
  INVX1 U169 ( .A(n149), .Y(n150) );
  AND2X1 U170 ( .A(n173), .B(n279), .Y(n151) );
  INVX1 U171 ( .A(n151), .Y(n152) );
  AND2X1 U172 ( .A(n280), .B(n4), .Y(n153) );
  INVX1 U173 ( .A(n153), .Y(n154) );
  AND2X1 U174 ( .A(n280), .B(n279), .Y(n155) );
  INVX1 U175 ( .A(n155), .Y(n156) );
  INVX1 U176 ( .A(n272), .Y(n157) );
  INVX1 U177 ( .A(n157), .Y(n158) );
  INVX1 U178 ( .A(n273), .Y(n159) );
  INVX1 U179 ( .A(n159), .Y(n160) );
  INVX1 U180 ( .A(n274), .Y(n161) );
  INVX1 U181 ( .A(n161), .Y(n162) );
  INVX1 U182 ( .A(n277), .Y(n163) );
  INVX1 U183 ( .A(n163), .Y(n164) );
  INVX1 U184 ( .A(n278), .Y(n165) );
  INVX1 U185 ( .A(n165), .Y(n166) );
  INVX1 U186 ( .A(n281), .Y(n167) );
  INVX1 U187 ( .A(n167), .Y(n168) );
  AND2X1 U188 ( .A(\Cnt<3> ), .B(n203), .Y(n171) );
  AND2X2 U189 ( .A(\Cnt<0> ), .B(n206), .Y(n172) );
  AND2X1 U190 ( .A(n211), .B(\Cnt<2> ), .Y(n173) );
  AND2X1 U191 ( .A(n201), .B(n40), .Y(n174) );
  AND2X2 U192 ( .A(n66), .B(n33), .Y(n176) );
  INVX1 U193 ( .A(n176), .Y(n177) );
  AND2X2 U194 ( .A(n69), .B(n35), .Y(n178) );
  INVX1 U195 ( .A(n178), .Y(n179) );
  AND2X2 U196 ( .A(n72), .B(n36), .Y(n180) );
  INVX1 U197 ( .A(n180), .Y(n181) );
  INVX1 U198 ( .A(n207), .Y(n182) );
  AND2X2 U199 ( .A(n65), .B(n91), .Y(n183) );
  INVX1 U200 ( .A(n183), .Y(n184) );
  AND2X2 U201 ( .A(n64), .B(n89), .Y(n185) );
  INVX1 U202 ( .A(n185), .Y(n186) );
  AND2X2 U203 ( .A(n67), .B(n34), .Y(n187) );
  INVX1 U204 ( .A(n187), .Y(n188) );
  AND2X2 U205 ( .A(n70), .B(n47), .Y(n189) );
  INVX1 U206 ( .A(n189), .Y(n190) );
  AND2X2 U207 ( .A(n74), .B(n37), .Y(n191) );
  INVX1 U208 ( .A(n191), .Y(n192) );
  AND2X2 U209 ( .A(n63), .B(n87), .Y(n193) );
  INVX1 U210 ( .A(n193), .Y(n194) );
  AND2X2 U211 ( .A(n68), .B(n93), .Y(n195) );
  INVX1 U212 ( .A(n195), .Y(n196) );
  AND2X2 U213 ( .A(n71), .B(n95), .Y(n197) );
  INVX1 U214 ( .A(n197), .Y(n198) );
  AND2X2 U215 ( .A(n75), .B(n97), .Y(n199) );
  INVX1 U216 ( .A(n199), .Y(n200) );
  INVX1 U217 ( .A(\Cnt<1> ), .Y(n206) );
  INVX4 U218 ( .A(n1), .Y(n259) );
  INVX8 U219 ( .A(n236), .Y(n257) );
  INVX8 U220 ( .A(n215), .Y(n280) );
  INVX8 U221 ( .A(n202), .Y(n201) );
  OR2X2 U222 ( .A(\Cnt<1> ), .B(\Cnt<0> ), .Y(n236) );
  AOI22X1 U223 ( .A(\In<9> ), .B(n172), .C(\In<8> ), .D(n257), .Y(n207) );
  AOI22X1 U224 ( .A(\In<12> ), .B(n257), .C(\In<13> ), .D(n172), .Y(n210) );
  AOI21X1 U225 ( .A(\In<14> ), .B(n259), .C(n104), .Y(n209) );
  AOI22X1 U226 ( .A(n171), .B(n8), .C(n40), .D(n194), .Y(n220) );
  AOI22X1 U227 ( .A(\In<4> ), .B(n257), .C(\In<5> ), .D(n172), .Y(n214) );
  AOI21X1 U228 ( .A(\In<6> ), .B(n259), .C(n106), .Y(n213) );
  OR2X2 U229 ( .A(\Cnt<2> ), .B(\Cnt<3> ), .Y(n215) );
  AOI22X1 U230 ( .A(\In<0> ), .B(n257), .C(\In<1> ), .D(n172), .Y(n218) );
  AOI21X1 U231 ( .A(\In<2> ), .B(n259), .C(n108), .Y(n217) );
  AOI22X1 U232 ( .A(n173), .B(n186), .C(n280), .D(n184), .Y(n219) );
  AND2X2 U233 ( .A(n201), .B(\In<0> ), .Y(n221) );
  MUX2X1 U234 ( .B(\In<15> ), .A(n221), .S(\Cnt<0> ), .Y(n248) );
  AOI22X1 U235 ( .A(\In<9> ), .B(n257), .C(\In<10> ), .D(n172), .Y(n226) );
  AOI21X1 U236 ( .A(\In<11> ), .B(n259), .C(n110), .Y(n225) );
  AOI22X1 U237 ( .A(\In<5> ), .B(n257), .C(\In<6> ), .D(n172), .Y(n229) );
  AOI21X1 U238 ( .A(\In<7> ), .B(n259), .C(n112), .Y(n228) );
  AOI22X1 U239 ( .A(\In<1> ), .B(n257), .C(\In<2> ), .D(n172), .Y(n232) );
  AOI21X1 U240 ( .A(\In<3> ), .B(n259), .C(n114), .Y(n231) );
  AOI22X1 U241 ( .A(n173), .B(n188), .C(n280), .D(n196), .Y(n233) );
  NAND3X1 U242 ( .A(n13), .B(n55), .C(n49), .Y(\Out<1> ) );
  INVX2 U243 ( .A(\In<1> ), .Y(n234) );
  OAI21X1 U244 ( .A(n170), .B(n234), .C(n99), .Y(n235) );
  AOI22X1 U245 ( .A(\In<10> ), .B(n257), .C(\In<11> ), .D(n172), .Y(n239) );
  INVX2 U246 ( .A(\In<13> ), .Y(n237) );
  AOI21X1 U247 ( .A(\In<12> ), .B(n259), .C(n116), .Y(n238) );
  AOI22X1 U248 ( .A(\In<6> ), .B(n257), .C(\In<7> ), .D(n172), .Y(n242) );
  AOI21X1 U249 ( .A(\In<8> ), .B(n259), .C(n118), .Y(n241) );
  AOI22X1 U250 ( .A(\In<2> ), .B(n257), .C(\In<3> ), .D(n172), .Y(n245) );
  INVX2 U251 ( .A(\In<5> ), .Y(n243) );
  AOI21X1 U252 ( .A(\In<4> ), .B(n259), .C(n120), .Y(n244) );
  AOI22X1 U253 ( .A(n173), .B(n190), .C(n280), .D(n198), .Y(n246) );
  NAND3X1 U254 ( .A(n16), .B(n59), .C(n51), .Y(\Out<2> ) );
  INVX2 U255 ( .A(\In<2> ), .Y(n247) );
  AOI21X1 U256 ( .A(\In<1> ), .B(n259), .C(n122), .Y(n250) );
  OR2X2 U257 ( .A(n248), .B(\Cnt<1> ), .Y(n249) );
  OAI21X1 U258 ( .A(n38), .B(n202), .C(n249), .Y(n279) );
  AOI22X1 U259 ( .A(\In<11> ), .B(n257), .C(\In<12> ), .D(n172), .Y(n253) );
  INVX2 U260 ( .A(\In<14> ), .Y(n251) );
  AOI21X1 U261 ( .A(\In<13> ), .B(n259), .C(n124), .Y(n252) );
  AOI22X1 U262 ( .A(\In<7> ), .B(n257), .C(\In<8> ), .D(n172), .Y(n256) );
  INVX2 U263 ( .A(\In<10> ), .Y(n254) );
  AOI21X1 U264 ( .A(\In<9> ), .B(n259), .C(n18), .Y(n255) );
  AOI22X1 U265 ( .A(\In<3> ), .B(n257), .C(\In<4> ), .D(n172), .Y(n261) );
  AOI21X1 U266 ( .A(\In<5> ), .B(n259), .C(n20), .Y(n260) );
  AOI22X1 U267 ( .A(n173), .B(n192), .C(n280), .D(n200), .Y(n262) );
  AOI22X1 U268 ( .A(n280), .B(n186), .C(n194), .D(n171), .Y(n263) );
  NAND3X1 U269 ( .A(n22), .B(n39), .C(n43), .Y(\Out<4> ) );
  AOI22X1 U270 ( .A(n173), .B(n177), .C(n196), .D(n174), .Y(n265) );
  AOI22X1 U271 ( .A(n280), .B(n188), .C(n171), .D(n4), .Y(n264) );
  AOI22X1 U272 ( .A(n173), .B(n179), .C(n198), .D(n174), .Y(n267) );
  AOI22X1 U273 ( .A(n280), .B(n190), .C(n171), .D(n6), .Y(n266) );
  AOI22X1 U274 ( .A(n173), .B(n181), .C(n200), .D(n174), .Y(n269) );
  AOI22X1 U275 ( .A(n280), .B(n192), .C(n171), .D(n279), .Y(n268) );
  AOI22X1 U276 ( .A(n186), .B(n174), .C(n184), .D(n62), .Y(n271) );
  AOI22X1 U277 ( .A(n194), .B(n173), .C(n8), .D(n280), .Y(n270) );
  AOI22X1 U278 ( .A(n188), .B(n174), .C(n196), .D(n62), .Y(n272) );
  NAND3X1 U279 ( .A(n126), .B(n150), .C(n158), .Y(\Out<9> ) );
  AOI22X1 U280 ( .A(n190), .B(n174), .C(n198), .D(n62), .Y(n273) );
  NAND3X1 U281 ( .A(n128), .B(n26), .C(n160), .Y(\Out<10> ) );
  AOI22X1 U282 ( .A(n192), .B(n174), .C(n200), .D(n62), .Y(n274) );
  NAND3X1 U283 ( .A(n130), .B(n152), .C(n162), .Y(\Out<11> ) );
  AOI22X1 U284 ( .A(n186), .B(n62), .C(n184), .D(n146), .Y(n276) );
  AOI22X1 U285 ( .A(n194), .B(n280), .C(n8), .D(n174), .Y(n275) );
  AOI22X1 U286 ( .A(n188), .B(n62), .C(n196), .D(n146), .Y(n277) );
  NAND3X1 U287 ( .A(n132), .B(n154), .C(n164), .Y(\Out<13> ) );
  AOI22X1 U288 ( .A(n190), .B(n62), .C(n198), .D(n146), .Y(n278) );
  NAND3X1 U289 ( .A(n134), .B(n28), .C(n166), .Y(\Out<14> ) );
  AOI22X1 U290 ( .A(n192), .B(n62), .C(n200), .D(n146), .Y(n281) );
  NAND3X1 U291 ( .A(n136), .B(n156), .C(n168), .Y(\Out<15> ) );
endmodule


module fulladder1_31 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_30 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_29 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_28 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_27 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_26 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_25 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_24 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_23 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_22 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_21 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_20 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_19 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_18 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_17 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  AND2X2 U1 ( .A(A), .B(B), .Y(G) );
  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
endmodule


module fulladder1_16 ( A, B, Cin, S, P, G );
  input A, B, Cin;
  output S, P, G;


  XOR2X1 U2 ( .A(Cin), .B(P), .Y(S) );
  XOR2X1 U3 ( .A(A), .B(B), .Y(P) );
  AND2X1 U1 ( .A(A), .B(B), .Y(G) );
endmodule


module cla4_11 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n11,
         n13, n14, n15, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37;

  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n18), .C(n20), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n20), .C(n19), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n16), .C(\G<2> ), .Y(n11) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n13) );
  OAI21X1 U13 ( .A(n9), .B(n20), .C(n19), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n14) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n15) );
  fulladder1_44 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_45 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_46 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n35), .G(n27) );
  fulladder1_47 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  AND2X1 U1 ( .A(n21), .B(n2), .Y(n10) );
  INVX1 U2 ( .A(\G<0> ), .Y(n21) );
  AND2X1 U3 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  INVX1 U4 ( .A(\P<2> ), .Y(n18) );
  AND2X1 U5 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X1 U6 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  INVX1 U7 ( .A(\G<3> ), .Y(n19) );
  AND2X1 U9 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  INVX1 U16 ( .A(\P<3> ), .Y(n20) );
  AND2X1 U17 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U18 ( .A(n1), .Y(n2) );
  BUFX2 U19 ( .A(n15), .Y(n3) );
  INVX1 U20 ( .A(n3), .Y(n17) );
  INVX1 U21 ( .A(n13), .Y(n16) );
  INVX1 U22 ( .A(n11), .Y(n4) );
  INVX1 U23 ( .A(n4), .Y(n5) );
  AND2X1 U24 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U25 ( .A(n6), .Y(n7) );
  INVX1 U26 ( .A(n9), .Y(n8) );
  BUFX2 U27 ( .A(n14), .Y(n9) );
  INVX1 U28 ( .A(n10), .Y(n12) );
  AND2X1 U29 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U30 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U31 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U32 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U33 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U34 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U35 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U36 ( .A(n22), .B(n23), .Y(\G<0> ) );
endmodule


module cla4_10 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n8), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n6), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n10), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_43 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_42 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_41 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_40 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n9), .S(\S<3> ), .P(n38), .G(n30) );
  AND2X1 U1 ( .A(n18), .B(n2), .Y(n12) );
  INVX1 U2 ( .A(\G<0> ), .Y(n18) );
  AND2X1 U3 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  INVX1 U4 ( .A(\P<2> ), .Y(n20) );
  AND2X1 U5 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  INVX1 U6 ( .A(\G<3> ), .Y(n21) );
  AND2X1 U7 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  INVX1 U9 ( .A(\P<3> ), .Y(n22) );
  AND2X2 U16 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U17 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U18 ( .A(n1), .Y(n2) );
  BUFX2 U19 ( .A(n39), .Y(n3) );
  INVX1 U20 ( .A(n3), .Y(n17) );
  BUFX2 U21 ( .A(n41), .Y(n4) );
  INVX1 U22 ( .A(n4), .Y(n19) );
  INVX1 U23 ( .A(n42), .Y(n5) );
  INVX1 U24 ( .A(n5), .Y(n6) );
  AND2X1 U25 ( .A(\P<1> ), .B(\P<0> ), .Y(n7) );
  INVX1 U26 ( .A(n7), .Y(n8) );
  INVX1 U27 ( .A(n10), .Y(n9) );
  BUFX2 U28 ( .A(n40), .Y(n10) );
  INVX1 U29 ( .A(n12), .Y(n16) );
  AND2X1 U30 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U31 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U32 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U33 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U34 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U35 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U36 ( .A(n23), .B(n24), .Y(\G<0> ) );
endmodule


module cla4_9 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n7), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n9), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_39 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_38 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_37 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_36 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n38), .G(n30) );
  AND2X1 U1 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  AND2X1 U2 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  AND2X1 U3 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  INVX1 U4 ( .A(\P<2> ), .Y(n20) );
  INVX1 U5 ( .A(\G<3> ), .Y(n21) );
  AND2X1 U6 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  INVX1 U7 ( .A(\P<3> ), .Y(n22) );
  AND2X2 U9 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U16 ( .A(n1), .Y(n2) );
  BUFX2 U17 ( .A(n39), .Y(n3) );
  INVX1 U18 ( .A(n3), .Y(n17) );
  BUFX2 U19 ( .A(n41), .Y(n4) );
  INVX1 U20 ( .A(n4), .Y(n19) );
  BUFX2 U21 ( .A(n42), .Y(n5) );
  AND2X1 U22 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U23 ( .A(n6), .Y(n7) );
  INVX1 U24 ( .A(n10), .Y(n8) );
  INVX1 U25 ( .A(n8), .Y(n9) );
  BUFX2 U26 ( .A(n40), .Y(n10) );
  AND2X2 U27 ( .A(n2), .B(n18), .Y(n12) );
  INVX1 U28 ( .A(n12), .Y(n16) );
  AND2X1 U29 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U30 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U31 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U32 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U33 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U34 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U35 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U36 ( .A(n23), .B(n24), .Y(\G<0> ) );
  INVX2 U37 ( .A(\G<0> ), .Y(n18) );
endmodule


module cla4_8 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n19), .C(n21), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n21), .C(n20), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n18), .C(\G<2> ), .Y(n41) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n40) );
  OAI21X1 U13 ( .A(n9), .B(n21), .C(n20), .Y(Cout) );
  AOI21X1 U14 ( .A(n16), .B(\P<2> ), .C(\G<2> ), .Y(n39) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n38) );
  fulladder1_35 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_34 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_33 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n1), .S(\S<2> ), .P(n35), .G(n27) );
  fulladder1_32 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  AND2X1 U1 ( .A(Cin), .B(\P<0> ), .Y(n2) );
  AND2X1 U2 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  AND2X1 U3 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X1 U4 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  INVX1 U5 ( .A(\P<2> ), .Y(n19) );
  INVX1 U6 ( .A(\G<3> ), .Y(n20) );
  AND2X1 U7 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  INVX1 U9 ( .A(\P<3> ), .Y(n21) );
  BUFX2 U16 ( .A(n16), .Y(n1) );
  INVX1 U17 ( .A(n38), .Y(n16) );
  INVX1 U18 ( .A(n2), .Y(n3) );
  BUFX2 U19 ( .A(n40), .Y(n4) );
  INVX1 U20 ( .A(n4), .Y(n18) );
  BUFX2 U21 ( .A(n41), .Y(n5) );
  AND2X1 U22 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U23 ( .A(n6), .Y(n7) );
  INVX1 U24 ( .A(n39), .Y(n8) );
  INVX1 U25 ( .A(n8), .Y(n9) );
  AND2X2 U26 ( .A(n3), .B(n17), .Y(n10) );
  INVX1 U27 ( .A(n10), .Y(n12) );
  AND2X1 U28 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U29 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U30 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U31 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U32 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U33 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U34 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U35 ( .A(n22), .B(n23), .Y(\G<0> ) );
  INVX2 U36 ( .A(\G<0> ), .Y(n17) );
endmodule


module rf ( .read1data({\read1data<15> , \read1data<14> , \read1data<13> , 
        \read1data<12> , \read1data<11> , \read1data<10> , \read1data<9> , 
        \read1data<8> , \read1data<7> , \read1data<6> , \read1data<5> , 
        \read1data<4> , \read1data<3> , \read1data<2> , \read1data<1> , 
        \read1data<0> }), .read2data({\read2data<15> , \read2data<14> , 
        \read2data<13> , \read2data<12> , \read2data<11> , \read2data<10> , 
        \read2data<9> , \read2data<8> , \read2data<7> , \read2data<6> , 
        \read2data<5> , \read2data<4> , \read2data<3> , \read2data<2> , 
        \read2data<1> , \read2data<0> }), err, clk, rst, .read1regsel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .read2regsel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .writeregsel({
        \writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   \rf_wr_en<7> , \rf_wr_en<6> , \rf_wr_en<5> , \rf_wr_en<4> ,
         \rf_wr_en<3> , \rf_wr_en<2> , \rf_wr_en<1> , \rf_wr_en<0> ,
         \write_en<7> , \write_en<6> , \write_en<5> , \write_en<4> ,
         \write_en<3> , \write_en<2> , \write_en<1> , \write_en<0> ,
         \reg_in<127> , \reg_in<126> , \reg_in<125> , \reg_in<124> ,
         \reg_in<123> , \reg_in<122> , \reg_in<121> , \reg_in<120> ,
         \reg_in<119> , \reg_in<118> , \reg_in<117> , \reg_in<116> ,
         \reg_in<115> , \reg_in<114> , \reg_in<113> , \reg_in<112> ,
         \reg_in<111> , \reg_in<110> , \reg_in<109> , \reg_in<108> ,
         \reg_in<107> , \reg_in<106> , \reg_in<105> , \reg_in<104> ,
         \reg_in<103> , \reg_in<102> , \reg_in<101> , \reg_in<100> ,
         \reg_in<99> , \reg_in<98> , \reg_in<97> , \reg_in<96> , \reg_in<95> ,
         \reg_in<94> , \reg_in<93> , \reg_in<92> , \reg_in<91> , \reg_in<90> ,
         \reg_in<89> , \reg_in<88> , \reg_in<87> , \reg_in<86> , \reg_in<85> ,
         \reg_in<84> , \reg_in<83> , \reg_in<82> , \reg_in<81> , \reg_in<80> ,
         \reg_in<79> , \reg_in<78> , \reg_in<77> , \reg_in<76> , \reg_in<75> ,
         \reg_in<74> , \reg_in<73> , \reg_in<72> , \reg_in<71> , \reg_in<70> ,
         \reg_in<69> , \reg_in<68> , \reg_in<67> , \reg_in<66> , \reg_in<65> ,
         \reg_in<64> , \reg_in<63> , \reg_in<62> , \reg_in<61> , \reg_in<60> ,
         \reg_in<59> , \reg_in<58> , \reg_in<57> , \reg_in<56> , \reg_in<55> ,
         \reg_in<54> , \reg_in<53> , \reg_in<52> , \reg_in<51> , \reg_in<50> ,
         \reg_in<49> , \reg_in<48> , \reg_in<47> , \reg_in<46> , \reg_in<45> ,
         \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> ,
         \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> ,
         \reg_in<34> , \reg_in<33> , \reg_in<32> , \reg_in<31> , \reg_in<30> ,
         \reg_in<29> , \reg_in<28> , \reg_in<27> , \reg_in<26> , \reg_in<25> ,
         \reg_in<24> , \reg_in<23> , \reg_in<22> , \reg_in<21> , \reg_in<20> ,
         \reg_in<19> , \reg_in<18> , \reg_in<17> , \reg_in<16> , \reg_in<15> ,
         \reg_in<14> , \reg_in<13> , \reg_in<12> , \reg_in<11> , \reg_in<10> ,
         \reg_in<9> , \reg_in<8> , \reg_in<7> , \reg_in<6> , \reg_in<5> ,
         \reg_in<4> , \reg_in<3> , \reg_in<2> , \reg_in<1> , \reg_in<0> ,
         \reg_out<127> , \reg_out<126> , \reg_out<125> , \reg_out<124> ,
         \reg_out<123> , \reg_out<122> , \reg_out<121> , \reg_out<120> ,
         \reg_out<119> , \reg_out<118> , \reg_out<117> , \reg_out<116> ,
         \reg_out<115> , \reg_out<114> , \reg_out<113> , \reg_out<112> ,
         \reg_out<111> , \reg_out<110> , \reg_out<109> , \reg_out<108> ,
         \reg_out<107> , \reg_out<106> , \reg_out<105> , \reg_out<104> ,
         \reg_out<103> , \reg_out<102> , \reg_out<101> , \reg_out<100> ,
         \reg_out<99> , \reg_out<98> , \reg_out<97> , \reg_out<96> ,
         \reg_out<95> , \reg_out<94> , \reg_out<93> , \reg_out<92> ,
         \reg_out<91> , \reg_out<90> , \reg_out<89> , \reg_out<88> ,
         \reg_out<87> , \reg_out<86> , \reg_out<85> , \reg_out<84> ,
         \reg_out<83> , \reg_out<82> , \reg_out<81> , \reg_out<80> ,
         \reg_out<79> , \reg_out<78> , \reg_out<77> , \reg_out<76> ,
         \reg_out<75> , \reg_out<74> , \reg_out<73> , \reg_out<72> ,
         \reg_out<71> , \reg_out<70> , \reg_out<69> , \reg_out<68> ,
         \reg_out<67> , \reg_out<66> , \reg_out<65> , \reg_out<64> ,
         \reg_out<63> , \reg_out<62> , \reg_out<61> , \reg_out<60> ,
         \reg_out<59> , \reg_out<58> , \reg_out<57> , \reg_out<56> ,
         \reg_out<55> , \reg_out<54> , \reg_out<53> , \reg_out<52> ,
         \reg_out<51> , \reg_out<50> , \reg_out<49> , \reg_out<48> ,
         \reg_out<47> , \reg_out<46> , \reg_out<45> , \reg_out<44> ,
         \reg_out<43> , \reg_out<42> , \reg_out<41> , \reg_out<40> ,
         \reg_out<39> , \reg_out<38> , \reg_out<37> , \reg_out<36> ,
         \reg_out<35> , \reg_out<34> , \reg_out<33> , \reg_out<32> ,
         \reg_out<31> , \reg_out<30> , \reg_out<29> , \reg_out<28> ,
         \reg_out<27> , \reg_out<26> , \reg_out<25> , \reg_out<24> ,
         \reg_out<23> , \reg_out<22> , \reg_out<21> , \reg_out<20> ,
         \reg_out<19> , \reg_out<18> , \reg_out<17> , \reg_out<16> ,
         \reg_out<15> , \reg_out<14> , \reg_out<13> , \reg_out<12> ,
         \reg_out<11> , \reg_out<10> , \reg_out<9> , \reg_out<8> ,
         \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , \reg_out<3> ,
         \reg_out<2> , \reg_out<1> , \reg_out<0> , n1, n2, n3, n4;
  assign err = 1'b0;

  register16_0 \registers[0]  ( .d({\reg_in<15> , \reg_in<14> , \reg_in<13> , 
        \reg_in<12> , \reg_in<11> , \reg_in<10> , \reg_in<9> , \reg_in<8> , 
        \reg_in<7> , \reg_in<6> , \reg_in<5> , \reg_in<4> , \reg_in<3> , 
        \reg_in<2> , \reg_in<1> , \reg_in<0> }), .clk(clk), .wr_en(
        \rf_wr_en<0> ), .rst(n3), .q({\reg_out<15> , \reg_out<14> , 
        \reg_out<13> , \reg_out<12> , \reg_out<11> , \reg_out<10> , 
        \reg_out<9> , \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , 
        \reg_out<4> , \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> })
         );
  register16_1 \registers[1]  ( .d({\reg_in<31> , \reg_in<30> , \reg_in<29> , 
        \reg_in<28> , \reg_in<27> , \reg_in<26> , \reg_in<25> , \reg_in<24> , 
        \reg_in<23> , \reg_in<22> , \reg_in<21> , \reg_in<20> , \reg_in<19> , 
        \reg_in<18> , \reg_in<17> , \reg_in<16> }), .clk(clk), .wr_en(
        \rf_wr_en<1> ), .rst(n3), .q({\reg_out<31> , \reg_out<30> , 
        \reg_out<29> , \reg_out<28> , \reg_out<27> , \reg_out<26> , 
        \reg_out<25> , \reg_out<24> , \reg_out<23> , \reg_out<22> , 
        \reg_out<21> , \reg_out<20> , \reg_out<19> , \reg_out<18> , 
        \reg_out<17> , \reg_out<16> }) );
  register16_2 \registers[2]  ( .d({\reg_in<47> , \reg_in<46> , \reg_in<45> , 
        \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> , 
        \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> , 
        \reg_in<34> , \reg_in<33> , \reg_in<32> }), .clk(clk), .wr_en(
        \rf_wr_en<2> ), .rst(n3), .q({\reg_out<47> , \reg_out<46> , 
        \reg_out<45> , \reg_out<44> , \reg_out<43> , \reg_out<42> , 
        \reg_out<41> , \reg_out<40> , \reg_out<39> , \reg_out<38> , 
        \reg_out<37> , \reg_out<36> , \reg_out<35> , \reg_out<34> , 
        \reg_out<33> , \reg_out<32> }) );
  register16_3 \registers[3]  ( .d({\reg_in<63> , \reg_in<62> , \reg_in<61> , 
        \reg_in<60> , \reg_in<59> , \reg_in<58> , \reg_in<57> , \reg_in<56> , 
        \reg_in<55> , \reg_in<54> , \reg_in<53> , \reg_in<52> , \reg_in<51> , 
        \reg_in<50> , \reg_in<49> , \reg_in<48> }), .clk(clk), .wr_en(
        \rf_wr_en<3> ), .rst(n3), .q({\reg_out<63> , \reg_out<62> , 
        \reg_out<61> , \reg_out<60> , \reg_out<59> , \reg_out<58> , 
        \reg_out<57> , \reg_out<56> , \reg_out<55> , \reg_out<54> , 
        \reg_out<53> , \reg_out<52> , \reg_out<51> , \reg_out<50> , 
        \reg_out<49> , \reg_out<48> }) );
  register16_4 \registers[4]  ( .d({\reg_in<79> , \reg_in<78> , \reg_in<77> , 
        \reg_in<76> , \reg_in<75> , \reg_in<74> , \reg_in<73> , \reg_in<72> , 
        \reg_in<71> , \reg_in<70> , \reg_in<69> , \reg_in<68> , \reg_in<67> , 
        \reg_in<66> , \reg_in<65> , \reg_in<64> }), .clk(clk), .wr_en(
        \rf_wr_en<4> ), .rst(n3), .q({\reg_out<79> , \reg_out<78> , 
        \reg_out<77> , \reg_out<76> , \reg_out<75> , \reg_out<74> , 
        \reg_out<73> , \reg_out<72> , \reg_out<71> , \reg_out<70> , 
        \reg_out<69> , \reg_out<68> , \reg_out<67> , \reg_out<66> , 
        \reg_out<65> , \reg_out<64> }) );
  register16_5 \registers[5]  ( .d({\reg_in<95> , \reg_in<94> , \reg_in<93> , 
        \reg_in<92> , \reg_in<91> , \reg_in<90> , \reg_in<89> , \reg_in<88> , 
        \reg_in<87> , \reg_in<86> , \reg_in<85> , \reg_in<84> , \reg_in<83> , 
        \reg_in<82> , \reg_in<81> , \reg_in<80> }), .clk(clk), .wr_en(
        \rf_wr_en<5> ), .rst(n3), .q({\reg_out<95> , \reg_out<94> , 
        \reg_out<93> , \reg_out<92> , \reg_out<91> , \reg_out<90> , 
        \reg_out<89> , \reg_out<88> , \reg_out<87> , \reg_out<86> , 
        \reg_out<85> , \reg_out<84> , \reg_out<83> , \reg_out<82> , 
        \reg_out<81> , \reg_out<80> }) );
  register16_6 \registers[6]  ( .d({\reg_in<111> , \reg_in<110> , 
        \reg_in<109> , \reg_in<108> , \reg_in<107> , \reg_in<106> , 
        \reg_in<105> , \reg_in<104> , \reg_in<103> , \reg_in<102> , 
        \reg_in<101> , \reg_in<100> , \reg_in<99> , \reg_in<98> , \reg_in<97> , 
        \reg_in<96> }), .clk(clk), .wr_en(\rf_wr_en<6> ), .rst(n3), .q({
        \reg_out<111> , \reg_out<110> , \reg_out<109> , \reg_out<108> , 
        \reg_out<107> , \reg_out<106> , \reg_out<105> , \reg_out<104> , 
        \reg_out<103> , \reg_out<102> , \reg_out<101> , \reg_out<100> , 
        \reg_out<99> , \reg_out<98> , \reg_out<97> , \reg_out<96> }) );
  register16_7 \registers[7]  ( .d({\reg_in<127> , \reg_in<126> , 
        \reg_in<125> , \reg_in<124> , \reg_in<123> , \reg_in<122> , 
        \reg_in<121> , \reg_in<120> , \reg_in<119> , \reg_in<118> , 
        \reg_in<117> , \reg_in<116> , \reg_in<115> , \reg_in<114> , 
        \reg_in<113> , \reg_in<112> }), .clk(clk), .wr_en(\rf_wr_en<7> ), 
        .rst(n3), .q({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> }) );
  decoder3to8 wr_dec ( .In({\writeregsel<2> , \writeregsel<1> , n1}), .Out({
        \write_en<7> , \write_en<6> , \write_en<5> , \write_en<4> , 
        \write_en<3> , \write_en<2> , \write_en<1> , \write_en<0> }) );
  mux8to1_16_1 read1_mux ( .In({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> , \reg_out<111> , \reg_out<110> , \reg_out<109> , 
        \reg_out<108> , \reg_out<107> , \reg_out<106> , \reg_out<105> , 
        \reg_out<104> , \reg_out<103> , \reg_out<102> , \reg_out<101> , 
        \reg_out<100> , \reg_out<99> , \reg_out<98> , \reg_out<97> , 
        \reg_out<96> , \reg_out<95> , \reg_out<94> , \reg_out<93> , 
        \reg_out<92> , \reg_out<91> , \reg_out<90> , \reg_out<89> , 
        \reg_out<88> , \reg_out<87> , \reg_out<86> , \reg_out<85> , 
        \reg_out<84> , \reg_out<83> , \reg_out<82> , \reg_out<81> , 
        \reg_out<80> , \reg_out<79> , \reg_out<78> , \reg_out<77> , 
        \reg_out<76> , \reg_out<75> , \reg_out<74> , \reg_out<73> , 
        \reg_out<72> , \reg_out<71> , \reg_out<70> , \reg_out<69> , 
        \reg_out<68> , \reg_out<67> , \reg_out<66> , \reg_out<65> , 
        \reg_out<64> , \reg_out<63> , \reg_out<62> , \reg_out<61> , 
        \reg_out<60> , \reg_out<59> , \reg_out<58> , \reg_out<57> , 
        \reg_out<56> , \reg_out<55> , \reg_out<54> , \reg_out<53> , 
        \reg_out<52> , \reg_out<51> , \reg_out<50> , \reg_out<49> , 
        \reg_out<48> , \reg_out<47> , \reg_out<46> , \reg_out<45> , 
        \reg_out<44> , \reg_out<43> , \reg_out<42> , \reg_out<41> , 
        \reg_out<40> , \reg_out<39> , \reg_out<38> , \reg_out<37> , 
        \reg_out<36> , \reg_out<35> , \reg_out<34> , \reg_out<33> , 
        \reg_out<32> , \reg_out<31> , \reg_out<30> , \reg_out<29> , 
        \reg_out<28> , \reg_out<27> , \reg_out<26> , \reg_out<25> , 
        \reg_out<24> , \reg_out<23> , \reg_out<22> , \reg_out<21> , 
        \reg_out<20> , \reg_out<19> , \reg_out<18> , \reg_out<17> , 
        \reg_out<16> , \reg_out<15> , \reg_out<14> , \reg_out<13> , 
        \reg_out<12> , \reg_out<11> , \reg_out<10> , \reg_out<9> , 
        \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , 
        \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> }), .Sel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .Out({
        \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> , 
        \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> , 
        \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> , 
        \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> }) );
  mux8to1_16_0 read2_mux ( .In({\reg_out<127> , \reg_out<126> , \reg_out<125> , 
        \reg_out<124> , \reg_out<123> , \reg_out<122> , \reg_out<121> , 
        \reg_out<120> , \reg_out<119> , \reg_out<118> , \reg_out<117> , 
        \reg_out<116> , \reg_out<115> , \reg_out<114> , \reg_out<113> , 
        \reg_out<112> , \reg_out<111> , \reg_out<110> , \reg_out<109> , 
        \reg_out<108> , \reg_out<107> , \reg_out<106> , \reg_out<105> , 
        \reg_out<104> , \reg_out<103> , \reg_out<102> , \reg_out<101> , 
        \reg_out<100> , \reg_out<99> , \reg_out<98> , \reg_out<97> , 
        \reg_out<96> , \reg_out<95> , \reg_out<94> , \reg_out<93> , 
        \reg_out<92> , \reg_out<91> , \reg_out<90> , \reg_out<89> , 
        \reg_out<88> , \reg_out<87> , \reg_out<86> , \reg_out<85> , 
        \reg_out<84> , \reg_out<83> , \reg_out<82> , \reg_out<81> , 
        \reg_out<80> , \reg_out<79> , \reg_out<78> , \reg_out<77> , 
        \reg_out<76> , \reg_out<75> , \reg_out<74> , \reg_out<73> , 
        \reg_out<72> , \reg_out<71> , \reg_out<70> , \reg_out<69> , 
        \reg_out<68> , \reg_out<67> , \reg_out<66> , \reg_out<65> , 
        \reg_out<64> , \reg_out<63> , \reg_out<62> , \reg_out<61> , 
        \reg_out<60> , \reg_out<59> , \reg_out<58> , \reg_out<57> , 
        \reg_out<56> , \reg_out<55> , \reg_out<54> , \reg_out<53> , 
        \reg_out<52> , \reg_out<51> , \reg_out<50> , \reg_out<49> , 
        \reg_out<48> , \reg_out<47> , \reg_out<46> , \reg_out<45> , 
        \reg_out<44> , \reg_out<43> , \reg_out<42> , \reg_out<41> , 
        \reg_out<40> , \reg_out<39> , \reg_out<38> , \reg_out<37> , 
        \reg_out<36> , \reg_out<35> , \reg_out<34> , \reg_out<33> , 
        \reg_out<32> , \reg_out<31> , \reg_out<30> , \reg_out<29> , 
        \reg_out<28> , \reg_out<27> , \reg_out<26> , \reg_out<25> , 
        \reg_out<24> , \reg_out<23> , \reg_out<22> , \reg_out<21> , 
        \reg_out<20> , \reg_out<19> , \reg_out<18> , \reg_out<17> , 
        \reg_out<16> , \reg_out<15> , \reg_out<14> , \reg_out<13> , 
        \reg_out<12> , \reg_out<11> , \reg_out<10> , \reg_out<9> , 
        \reg_out<8> , \reg_out<7> , \reg_out<6> , \reg_out<5> , \reg_out<4> , 
        \reg_out<3> , \reg_out<2> , \reg_out<1> , \reg_out<0> }), .Sel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .Out({
        \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> , 
        \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> , 
        \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> , 
        \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> }) );
  demux1to8_16 wr_demux ( .In({\writedata<15> , \writedata<14> , 
        \writedata<13> , \writedata<12> , \writedata<11> , \writedata<10> , 
        \writedata<9> , \writedata<8> , \writedata<7> , \writedata<6> , 
        \writedata<5> , \writedata<4> , \writedata<3> , \writedata<2> , 
        \writedata<1> , \writedata<0> }), .S({\writeregsel<2> , 
        \writeregsel<1> , n1}), .Out0({\reg_in<15> , \reg_in<14> , 
        \reg_in<13> , \reg_in<12> , \reg_in<11> , \reg_in<10> , \reg_in<9> , 
        \reg_in<8> , \reg_in<7> , \reg_in<6> , \reg_in<5> , \reg_in<4> , 
        \reg_in<3> , \reg_in<2> , \reg_in<1> , \reg_in<0> }), .Out1({
        \reg_in<31> , \reg_in<30> , \reg_in<29> , \reg_in<28> , \reg_in<27> , 
        \reg_in<26> , \reg_in<25> , \reg_in<24> , \reg_in<23> , \reg_in<22> , 
        \reg_in<21> , \reg_in<20> , \reg_in<19> , \reg_in<18> , \reg_in<17> , 
        \reg_in<16> }), .Out2({\reg_in<47> , \reg_in<46> , \reg_in<45> , 
        \reg_in<44> , \reg_in<43> , \reg_in<42> , \reg_in<41> , \reg_in<40> , 
        \reg_in<39> , \reg_in<38> , \reg_in<37> , \reg_in<36> , \reg_in<35> , 
        \reg_in<34> , \reg_in<33> , \reg_in<32> }), .Out3({\reg_in<63> , 
        \reg_in<62> , \reg_in<61> , \reg_in<60> , \reg_in<59> , \reg_in<58> , 
        \reg_in<57> , \reg_in<56> , \reg_in<55> , \reg_in<54> , \reg_in<53> , 
        \reg_in<52> , \reg_in<51> , \reg_in<50> , \reg_in<49> , \reg_in<48> }), 
        .Out4({\reg_in<79> , \reg_in<78> , \reg_in<77> , \reg_in<76> , 
        \reg_in<75> , \reg_in<74> , \reg_in<73> , \reg_in<72> , \reg_in<71> , 
        \reg_in<70> , \reg_in<69> , \reg_in<68> , \reg_in<67> , \reg_in<66> , 
        \reg_in<65> , \reg_in<64> }), .Out5({\reg_in<95> , \reg_in<94> , 
        \reg_in<93> , \reg_in<92> , \reg_in<91> , \reg_in<90> , \reg_in<89> , 
        \reg_in<88> , \reg_in<87> , \reg_in<86> , \reg_in<85> , \reg_in<84> , 
        \reg_in<83> , \reg_in<82> , \reg_in<81> , \reg_in<80> }), .Out6({
        \reg_in<111> , \reg_in<110> , \reg_in<109> , \reg_in<108> , 
        \reg_in<107> , \reg_in<106> , \reg_in<105> , \reg_in<104> , 
        \reg_in<103> , \reg_in<102> , \reg_in<101> , \reg_in<100> , 
        \reg_in<99> , \reg_in<98> , \reg_in<97> , \reg_in<96> }), .Out7({
        \reg_in<127> , \reg_in<126> , \reg_in<125> , \reg_in<124> , 
        \reg_in<123> , \reg_in<122> , \reg_in<121> , \reg_in<120> , 
        \reg_in<119> , \reg_in<118> , \reg_in<117> , \reg_in<116> , 
        \reg_in<115> , \reg_in<114> , \reg_in<113> , \reg_in<112> }) );
  AND2X1 U2 ( .A(\write_en<0> ), .B(write), .Y(\rf_wr_en<0> ) );
  AND2X1 U3 ( .A(\write_en<1> ), .B(write), .Y(\rf_wr_en<1> ) );
  AND2X1 U4 ( .A(\write_en<2> ), .B(write), .Y(\rf_wr_en<2> ) );
  AND2X1 U5 ( .A(\write_en<3> ), .B(write), .Y(\rf_wr_en<3> ) );
  AND2X1 U6 ( .A(\write_en<4> ), .B(write), .Y(\rf_wr_en<4> ) );
  AND2X1 U7 ( .A(\write_en<5> ), .B(write), .Y(\rf_wr_en<5> ) );
  AND2X1 U8 ( .A(\write_en<6> ), .B(write), .Y(\rf_wr_en<6> ) );
  AND2X1 U9 ( .A(\write_en<7> ), .B(write), .Y(\rf_wr_en<7> ) );
  INVX2 U10 ( .A(n2), .Y(n1) );
  INVX1 U11 ( .A(\writeregsel<0> ), .Y(n2) );
  INVX2 U12 ( .A(n4), .Y(n3) );
  INVX1 U13 ( .A(rst), .Y(n4) );
endmodule


module demux1to2_16_1 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), S, .Out0({\Out0<15> , \Out0<14> , 
        \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , \Out0<9> , \Out0<8> , 
        \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , \Out0<3> , \Out0<2> , 
        \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , \Out1<14> , \Out1<13> , 
        \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , \Out1<8> , \Out1<7> , 
        \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , \Out1<2> , \Out1<1> , 
        \Out1<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , S;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> ;
  wire   n1, n2, n3;

  demux1to2_17 \d[0]  ( .In(\In<0> ), .S(n1), .Out0(\Out0<0> ), .Out1(
        \Out1<0> ) );
  demux1to2_18 \d[1]  ( .In(\In<1> ), .S(n2), .Out0(\Out0<1> ), .Out1(
        \Out1<1> ) );
  demux1to2_19 \d[2]  ( .In(\In<2> ), .S(n1), .Out0(\Out0<2> ), .Out1(
        \Out1<2> ) );
  demux1to2_20 \d[3]  ( .In(\In<3> ), .S(n1), .Out0(\Out0<3> ), .Out1(
        \Out1<3> ) );
  demux1to2_21 \d[4]  ( .In(\In<4> ), .S(S), .Out0(\Out0<4> ), .Out1(\Out1<4> ) );
  demux1to2_22 \d[5]  ( .In(\In<5> ), .S(n2), .Out0(\Out0<5> ), .Out1(
        \Out1<5> ) );
  demux1to2_23 \d[6]  ( .In(\In<6> ), .S(n1), .Out0(\Out0<6> ), .Out1(
        \Out1<6> ) );
  demux1to2_24 \d[7]  ( .In(\In<7> ), .S(n2), .Out0(\Out0<7> ), .Out1(
        \Out1<7> ) );
  demux1to2_25 \d[8]  ( .In(\In<8> ), .S(n2), .Out0(\Out0<8> ), .Out1(
        \Out1<8> ) );
  demux1to2_26 \d[9]  ( .In(\In<9> ), .S(n2), .Out0(\Out0<9> ), .Out1(
        \Out1<9> ) );
  demux1to2_27 \d[10]  ( .In(\In<10> ), .S(S), .Out0(\Out0<10> ), .Out1(
        \Out1<10> ) );
  demux1to2_28 \d[11]  ( .In(\In<11> ), .S(n2), .Out0(\Out0<11> ), .Out1(
        \Out1<11> ) );
  demux1to2_29 \d[12]  ( .In(\In<12> ), .S(S), .Out0(\Out0<12> ), .Out1(
        \Out1<12> ) );
  demux1to2_30 \d[13]  ( .In(\In<13> ), .S(n2), .Out0(\Out0<13> ), .Out1(
        \Out1<13> ) );
  demux1to2_31 \d[14]  ( .In(\In<14> ), .S(S), .Out0(\Out0<14> ), .Out1(
        \Out1<14> ) );
  demux1to2_32 \d[15]  ( .In(\In<15> ), .S(n1), .Out0(\Out0<15> ), .Out1(
        \Out1<15> ) );
  INVX8 U1 ( .A(n3), .Y(n1) );
  INVX8 U2 ( .A(n3), .Y(n2) );
  INVX8 U3 ( .A(S), .Y(n3) );
endmodule


module demux1to2_16_0 ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), S, .Out0({\Out0<15> , \Out0<14> , 
        \Out0<13> , \Out0<12> , \Out0<11> , \Out0<10> , \Out0<9> , \Out0<8> , 
        \Out0<7> , \Out0<6> , \Out0<5> , \Out0<4> , \Out0<3> , \Out0<2> , 
        \Out0<1> , \Out0<0> }), .Out1({\Out1<15> , \Out1<14> , \Out1<13> , 
        \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> , \Out1<8> , \Out1<7> , 
        \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> , \Out1<2> , \Out1<1> , 
        \Out1<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , S;
  output \Out0<15> , \Out0<14> , \Out0<13> , \Out0<12> , \Out0<11> ,
         \Out0<10> , \Out0<9> , \Out0<8> , \Out0<7> , \Out0<6> , \Out0<5> ,
         \Out0<4> , \Out0<3> , \Out0<2> , \Out0<1> , \Out0<0> , \Out1<15> ,
         \Out1<14> , \Out1<13> , \Out1<12> , \Out1<11> , \Out1<10> , \Out1<9> ,
         \Out1<8> , \Out1<7> , \Out1<6> , \Out1<5> , \Out1<4> , \Out1<3> ,
         \Out1<2> , \Out1<1> , \Out1<0> ;
  wire   n1, n2;

  demux1to2_15 \d[0]  ( .In(\In<0> ), .S(n1), .Out0(\Out0<0> ), .Out1(
        \Out1<0> ) );
  demux1to2_14 \d[1]  ( .In(\In<1> ), .S(n1), .Out0(\Out0<1> ), .Out1(
        \Out1<1> ) );
  demux1to2_13 \d[2]  ( .In(\In<2> ), .S(n1), .Out0(\Out0<2> ), .Out1(
        \Out1<2> ) );
  demux1to2_12 \d[3]  ( .In(\In<3> ), .S(n1), .Out0(\Out0<3> ), .Out1(
        \Out1<3> ) );
  demux1to2_11 \d[4]  ( .In(\In<4> ), .S(n1), .Out0(\Out0<4> ), .Out1(
        \Out1<4> ) );
  demux1to2_10 \d[5]  ( .In(\In<5> ), .S(n1), .Out0(\Out0<5> ), .Out1(
        \Out1<5> ) );
  demux1to2_9 \d[6]  ( .In(\In<6> ), .S(n1), .Out0(\Out0<6> ), .Out1(\Out1<6> ) );
  demux1to2_8 \d[7]  ( .In(\In<7> ), .S(n1), .Out0(\Out0<7> ), .Out1(\Out1<7> ) );
  demux1to2_7 \d[8]  ( .In(\In<8> ), .S(n1), .Out0(\Out0<8> ), .Out1(\Out1<8> ) );
  demux1to2_6 \d[9]  ( .In(\In<9> ), .S(n1), .Out0(\Out0<9> ), .Out1(\Out1<9> ) );
  demux1to2_5 \d[10]  ( .In(\In<10> ), .S(n1), .Out0(\Out0<10> ), .Out1(
        \Out1<10> ) );
  demux1to2_4 \d[11]  ( .In(\In<11> ), .S(n1), .Out0(\Out0<11> ), .Out1(
        \Out1<11> ) );
  demux1to2_3 \d[12]  ( .In(\In<12> ), .S(n1), .Out0(\Out0<12> ), .Out1(
        \Out1<12> ) );
  demux1to2_2 \d[13]  ( .In(\In<13> ), .S(n1), .Out0(\Out0<13> ), .Out1(
        \Out1<13> ) );
  demux1to2_1 \d[14]  ( .In(\In<14> ), .S(n1), .Out0(\Out0<14> ), .Out1(
        \Out1<14> ) );
  demux1to2_0 \d[15]  ( .In(\In<15> ), .S(n1), .Out0(\Out0<15> ), .Out1(
        \Out1<15> ) );
  INVX8 U1 ( .A(n2), .Y(n1) );
  INVX8 U2 ( .A(S), .Y(n2) );
endmodule


module cla_or_xor_and ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , 
        \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , 
        \B<3> , \B<2> , \B<1> , \B<0> }), Cin, .Op({\Op<1> , \Op<0> }), .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<1> , \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Cout;
  wire   cla_cout, \op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> ,
         \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> ,
         \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> ,
         \op0_A<1> , \op0_A<0> , \op1_A<15> , \op1_A<14> , \op1_A<13> ,
         \op1_A<12> , \op1_A<11> , \op1_A<10> , \op1_A<9> , \op1_A<8> ,
         \op1_A<7> , \op1_A<6> , \op1_A<5> , \op1_A<4> , \op1_A<3> ,
         \op1_A<2> , \op1_A<1> , \op1_A<0> , \op2_A<15> , \op2_A<14> ,
         \op2_A<13> , \op2_A<12> , \op2_A<11> , \op2_A<10> , \op2_A<9> ,
         \op2_A<8> , \op2_A<7> , \op2_A<6> , \op2_A<5> , \op2_A<4> ,
         \op2_A<3> , \op2_A<2> , \op2_A<1> , \op2_A<0> , \op3_A<15> ,
         \op3_A<14> , \op3_A<13> , \op3_A<12> , \op3_A<11> , \op3_A<10> ,
         \op3_A<9> , \op3_A<8> , \op3_A<7> , \op3_A<6> , \op3_A<5> ,
         \op3_A<4> , \op3_A<3> , \op3_A<2> , \op3_A<1> , \op3_A<0> ,
         \op0_B<15> , \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> ,
         \op0_B<10> , \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> ,
         \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , \op0_B<1> ,
         \op0_B<0> , \op1_B<15> , \op1_B<14> , \op1_B<13> , \op1_B<12> ,
         \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , \op1_B<7> ,
         \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> ,
         \op1_B<1> , \op1_B<0> , \op2_B<15> , \op2_B<14> , \op2_B<13> ,
         \op2_B<12> , \op2_B<11> , \op2_B<10> , \op2_B<9> , \op2_B<8> ,
         \op2_B<7> , \op2_B<6> , \op2_B<5> , \op2_B<4> , \op2_B<3> ,
         \op2_B<2> , \op2_B<1> , \op2_B<0> , \op3_B<15> , \op3_B<14> ,
         \op3_B<13> , \op3_B<12> , \op3_B<11> , \op3_B<10> , \op3_B<9> ,
         \op3_B<8> , \op3_B<7> , \op3_B<6> , \op3_B<5> , \op3_B<4> ,
         \op3_B<3> , \op3_B<2> , \op3_B<1> , \op3_B<0> , \op0_out<15> ,
         \op0_out<14> , \op0_out<13> , \op0_out<12> , \op0_out<11> ,
         \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , \op0_out<6> ,
         \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , \op0_out<1> ,
         \op0_out<0> , \op1_out<13> , \op1_out<12> , \op1_out<11> ,
         \op1_out<10> , \op1_out<6> , \op1_out<5> , \op2_out<15> ,
         \op2_out<14> , \op2_out<13> , \op2_out<12> , \op2_out<11> ,
         \op2_out<10> , \op2_out<9> , \op2_out<8> , \op2_out<7> , \op2_out<6> ,
         \op2_out<5> , \op2_out<4> , \op2_out<3> , \op2_out<2> , \op2_out<1> ,
         \op2_out<0> , \op3_out<15> , \op3_out<14> , \op3_out<13> ,
         \op3_out<12> , \op3_out<11> , \op3_out<10> , \op3_out<9> ,
         \op3_out<8> , \op3_out<7> , \op3_out<6> , \op3_out<5> , \op3_out<4> ,
         \op3_out<3> , \op3_out<2> , \op3_out<1> , \op3_out<0> , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50;

  AND2X2 U6 ( .A(\op3_B<5> ), .B(\op3_A<5> ), .Y(\op3_out<5> ) );
  XOR2X1 U46 ( .A(\op2_B<13> ), .B(\op2_A<13> ), .Y(\op2_out<13> ) );
  XOR2X1 U47 ( .A(\op2_B<12> ), .B(\op2_A<12> ), .Y(\op2_out<12> ) );
  XOR2X1 U48 ( .A(\op2_B<11> ), .B(\op2_A<11> ), .Y(\op2_out<11> ) );
  XOR2X1 U49 ( .A(\op2_B<10> ), .B(\op2_A<10> ), .Y(\op2_out<10> ) );
  demux1to4_16_1 demux0 ( .In({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , 
        \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , 
        \A<2> , \A<1> , \A<0> }), .S({n22, \Op<0> }), .Out0({\op0_A<15> , 
        \op0_A<14> , \op0_A<13> , \op0_A<12> , \op0_A<11> , \op0_A<10> , 
        \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , \op0_A<5> , \op0_A<4> , 
        \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .Out1({\op1_A<15> , 
        \op1_A<14> , \op1_A<13> , \op1_A<12> , \op1_A<11> , \op1_A<10> , 
        \op1_A<9> , \op1_A<8> , \op1_A<7> , \op1_A<6> , \op1_A<5> , \op1_A<4> , 
        \op1_A<3> , \op1_A<2> , \op1_A<1> , \op1_A<0> }), .Out2({\op2_A<15> , 
        \op2_A<14> , \op2_A<13> , \op2_A<12> , \op2_A<11> , \op2_A<10> , 
        \op2_A<9> , \op2_A<8> , \op2_A<7> , \op2_A<6> , \op2_A<5> , \op2_A<4> , 
        \op2_A<3> , \op2_A<2> , \op2_A<1> , \op2_A<0> }), .Out3({\op3_A<15> , 
        \op3_A<14> , \op3_A<13> , \op3_A<12> , \op3_A<11> , \op3_A<10> , 
        \op3_A<9> , \op3_A<8> , \op3_A<7> , \op3_A<6> , \op3_A<5> , \op3_A<4> , 
        \op3_A<3> , \op3_A<2> , \op3_A<1> , \op3_A<0> }) );
  demux1to4_16_0 demux1 ( .In({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , 
        \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , 
        \B<2> , \B<1> , \B<0> }), .S({n22, \Op<0> }), .Out0({\op0_B<15> , 
        \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , \op0_B<10> , 
        \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , 
        \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }), .Out1({\op1_B<15> , 
        \op1_B<14> , \op1_B<13> , \op1_B<12> , \op1_B<11> , \op1_B<10> , 
        \op1_B<9> , \op1_B<8> , \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , 
        \op1_B<3> , \op1_B<2> , \op1_B<1> , \op1_B<0> }), .Out2({\op2_B<15> , 
        \op2_B<14> , \op2_B<13> , \op2_B<12> , \op2_B<11> , \op2_B<10> , 
        \op2_B<9> , \op2_B<8> , \op2_B<7> , \op2_B<6> , \op2_B<5> , \op2_B<4> , 
        \op2_B<3> , \op2_B<2> , \op2_B<1> , \op2_B<0> }), .Out3({\op3_B<15> , 
        \op3_B<14> , \op3_B<13> , \op3_B<12> , \op3_B<11> , \op3_B<10> , 
        \op3_B<9> , \op3_B<8> , \op3_B<7> , \op3_B<6> , \op3_B<5> , \op3_B<4> , 
        \op3_B<3> , \op3_B<2> , \op3_B<1> , \op3_B<0> }) );
  cla16_0 cla0 ( .A({\op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> , n21, 
        \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , 
        \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .B({\op0_B<15> , \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , 
        \op0_B<10> , \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , 
        \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }), .Cin(Cin), .S({\op0_out<15> , \op0_out<14> , \op0_out<13> , \op0_out<12> , 
        \op0_out<11> , \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , 
        \op0_out<6> , \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , 
        \op0_out<1> , \op0_out<0> }), .Cout(cla_cout) );
  mux4to1_16_4 mux0 ( .InA({\op0_out<15> , \op0_out<14> , \op0_out<13> , 
        \op0_out<12> , \op0_out<11> , \op0_out<10> , \op0_out<9> , 
        \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , \op0_out<4> , 
        \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> }), .InB({n12, 
        n10, \op1_out<13> , \op1_out<12> , \op1_out<11> , \op1_out<10> , n8, 
        n20, n18, \op1_out<6> , \op1_out<5> , n16, n2, n14, n6, n4}), .InC({
        \op2_out<15> , \op2_out<14> , \op2_out<13> , \op2_out<12> , 
        \op2_out<11> , \op2_out<10> , \op2_out<9> , \op2_out<8> , \op2_out<7> , 
        \op2_out<6> , \op2_out<5> , \op2_out<4> , \op2_out<3> , \op2_out<2> , 
        \op2_out<1> , \op2_out<0> }), .InD({\op3_out<15> , \op3_out<14> , 
        \op3_out<13> , \op3_out<12> , \op3_out<11> , \op3_out<10> , 
        \op3_out<9> , \op3_out<8> , \op3_out<7> , \op3_out<6> , \op3_out<5> , 
        \op3_out<4> , \op3_out<3> , \op3_out<2> , \op3_out<1> , \op3_out<0> }), 
        .S({n22, \Op<0> }), .Out({\Out<15> , \Out<14> , \Out<13> , \Out<12> , 
        \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , 
        \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> }) );
  INVX1 U2 ( .A(\op1_A<7> ), .Y(n40) );
  OR2X1 U3 ( .A(\op1_A<11> ), .B(\op1_B<11> ), .Y(\op1_out<11> ) );
  AND2X1 U4 ( .A(\op3_B<11> ), .B(\op3_A<11> ), .Y(\op3_out<11> ) );
  AND2X1 U5 ( .A(\op3_A<14> ), .B(\op3_B<14> ), .Y(\op3_out<14> ) );
  OR2X1 U7 ( .A(\op1_A<10> ), .B(\op1_B<10> ), .Y(\op1_out<10> ) );
  AND2X1 U8 ( .A(\op3_B<10> ), .B(\op3_A<10> ), .Y(\op3_out<10> ) );
  AND2X1 U9 ( .A(\op3_A<7> ), .B(\op3_B<7> ), .Y(\op3_out<7> ) );
  INVX1 U10 ( .A(\op1_A<3> ), .Y(n36) );
  OR2X1 U11 ( .A(\op1_A<5> ), .B(\op1_B<5> ), .Y(\op1_out<5> ) );
  OR2X1 U12 ( .A(\op1_A<6> ), .B(\op1_B<6> ), .Y(\op1_out<6> ) );
  AND2X1 U13 ( .A(\op3_A<6> ), .B(\op3_B<6> ), .Y(\op3_out<6> ) );
  AND2X1 U14 ( .A(\op3_B<13> ), .B(\op3_A<13> ), .Y(\op3_out<13> ) );
  OR2X1 U15 ( .A(\op1_A<13> ), .B(\op1_B<13> ), .Y(\op1_out<13> ) );
  OR2X1 U16 ( .A(\op1_A<12> ), .B(\op1_B<12> ), .Y(\op1_out<12> ) );
  AND2X1 U17 ( .A(\op3_B<12> ), .B(\op3_A<12> ), .Y(\op3_out<12> ) );
  AND2X1 U18 ( .A(n37), .B(n36), .Y(n1) );
  INVX1 U19 ( .A(n1), .Y(n2) );
  AND2X1 U20 ( .A(n31), .B(n30), .Y(n3) );
  INVX1 U21 ( .A(n3), .Y(n4) );
  AND2X1 U22 ( .A(n33), .B(n32), .Y(n5) );
  INVX1 U23 ( .A(n5), .Y(n6) );
  AND2X1 U24 ( .A(n45), .B(n44), .Y(n7) );
  INVX1 U25 ( .A(n7), .Y(n8) );
  AND2X1 U26 ( .A(n47), .B(n46), .Y(n9) );
  INVX1 U27 ( .A(n9), .Y(n10) );
  AND2X1 U28 ( .A(n49), .B(n48), .Y(n11) );
  INVX1 U29 ( .A(n11), .Y(n12) );
  INVX1 U30 ( .A(cla_cout), .Y(n50) );
  INVX1 U31 ( .A(\op1_B<15> ), .Y(n49) );
  INVX1 U32 ( .A(\op1_B<14> ), .Y(n47) );
  INVX1 U33 ( .A(\op1_B<9> ), .Y(n45) );
  INVX1 U34 ( .A(\op1_B<8> ), .Y(n43) );
  INVX1 U35 ( .A(\op1_B<7> ), .Y(n41) );
  INVX1 U36 ( .A(\op1_B<4> ), .Y(n39) );
  INVX1 U37 ( .A(\op1_B<3> ), .Y(n37) );
  INVX1 U38 ( .A(\op1_B<2> ), .Y(n35) );
  INVX1 U39 ( .A(\op1_B<1> ), .Y(n33) );
  INVX1 U40 ( .A(\op1_B<0> ), .Y(n31) );
  INVX1 U41 ( .A(\op2_A<15> ), .Y(n29) );
  INVX1 U42 ( .A(\op2_A<14> ), .Y(n28) );
  INVX1 U43 ( .A(\op2_A<8> ), .Y(n27) );
  INVX1 U44 ( .A(\op2_A<4> ), .Y(n26) );
  AND2X1 U45 ( .A(n35), .B(n34), .Y(n13) );
  INVX1 U50 ( .A(n13), .Y(n14) );
  AND2X1 U51 ( .A(n39), .B(n38), .Y(n15) );
  INVX1 U52 ( .A(n15), .Y(n16) );
  AND2X1 U53 ( .A(n41), .B(n40), .Y(n17) );
  INVX1 U54 ( .A(n17), .Y(n18) );
  AND2X1 U55 ( .A(n43), .B(n42), .Y(n19) );
  INVX1 U56 ( .A(n19), .Y(n20) );
  INVX4 U57 ( .A(\Op<1> ), .Y(n23) );
  BUFX4 U58 ( .A(\op0_A<11> ), .Y(n21) );
  INVX8 U59 ( .A(n23), .Y(n22) );
  AND2X2 U60 ( .A(\op3_A<0> ), .B(\op3_B<0> ), .Y(\op3_out<0> ) );
  AND2X2 U61 ( .A(\op3_A<1> ), .B(\op3_B<1> ), .Y(\op3_out<1> ) );
  AND2X2 U62 ( .A(\op3_A<2> ), .B(\op3_B<2> ), .Y(\op3_out<2> ) );
  AND2X2 U63 ( .A(\op3_A<3> ), .B(\op3_B<3> ), .Y(\op3_out<3> ) );
  AND2X2 U64 ( .A(\op3_A<4> ), .B(\op3_B<4> ), .Y(\op3_out<4> ) );
  AND2X2 U65 ( .A(\op3_A<8> ), .B(\op3_B<8> ), .Y(\op3_out<8> ) );
  AND2X2 U66 ( .A(\op3_A<9> ), .B(\op3_B<9> ), .Y(\op3_out<9> ) );
  AND2X2 U67 ( .A(\op3_A<15> ), .B(\op3_B<15> ), .Y(\op3_out<15> ) );
  XOR2X1 U68 ( .A(\op2_A<0> ), .B(\op2_B<0> ), .Y(\op2_out<0> ) );
  INVX2 U69 ( .A(\op2_A<1> ), .Y(n24) );
  XNOR2X1 U70 ( .A(\op2_B<1> ), .B(n24), .Y(\op2_out<1> ) );
  INVX2 U71 ( .A(\op2_A<2> ), .Y(n25) );
  XNOR2X1 U72 ( .A(\op2_B<2> ), .B(n25), .Y(\op2_out<2> ) );
  XOR2X1 U73 ( .A(\op2_A<3> ), .B(\op2_B<3> ), .Y(\op2_out<3> ) );
  XNOR2X1 U74 ( .A(\op2_B<4> ), .B(n26), .Y(\op2_out<4> ) );
  XOR2X1 U75 ( .A(\op2_A<5> ), .B(\op2_B<5> ), .Y(\op2_out<5> ) );
  XOR2X1 U76 ( .A(\op2_A<6> ), .B(\op2_B<6> ), .Y(\op2_out<6> ) );
  XOR2X1 U77 ( .A(\op2_A<7> ), .B(\op2_B<7> ), .Y(\op2_out<7> ) );
  XNOR2X1 U78 ( .A(\op2_B<8> ), .B(n27), .Y(\op2_out<8> ) );
  XOR2X1 U79 ( .A(\op2_A<9> ), .B(\op2_B<9> ), .Y(\op2_out<9> ) );
  XNOR2X1 U80 ( .A(\op2_B<14> ), .B(n28), .Y(\op2_out<14> ) );
  XNOR2X1 U81 ( .A(\op2_B<15> ), .B(n29), .Y(\op2_out<15> ) );
  INVX2 U82 ( .A(\op1_A<0> ), .Y(n30) );
  INVX2 U83 ( .A(\op1_A<1> ), .Y(n32) );
  INVX2 U84 ( .A(\op1_A<2> ), .Y(n34) );
  INVX2 U85 ( .A(\op1_A<4> ), .Y(n38) );
  INVX2 U86 ( .A(\op1_A<8> ), .Y(n42) );
  INVX2 U87 ( .A(\op1_A<9> ), .Y(n44) );
  INVX2 U88 ( .A(\op1_A<14> ), .Y(n46) );
  INVX2 U89 ( .A(\op1_A<15> ), .Y(n48) );
  NOR3X1 U90 ( .A(n22), .B(\Op<0> ), .C(n50), .Y(Cout) );
endmodule


module shifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Op({\Op<1> , \Op<0> }), .Out({\Out<15> , 
        \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , 
        \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , 
        \Out<1> , \Out<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , \Op<1> ,
         \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   \ls_out<15> , \ls_out<14> , \ls_out<13> , \ls_out<12> , \ls_out<11> ,
         \ls_out<10> , \ls_out<9> , \ls_out<8> , \ls_out<7> , \ls_out<6> ,
         \ls_out<5> , \ls_out<4> , \ls_out<3> , \ls_out<2> , \ls_out<1> ,
         \ls_out<0> , \rs_out<15> , \rs_out<14> , \rs_out<13> , \rs_out<12> ,
         \rs_out<11> , \rs_out<10> , \rs_out<9> , \rs_out<8> , \rs_out<7> ,
         \rs_out<6> , \rs_out<5> , \rs_out<4> , \rs_out<3> , \rs_out<2> ,
         \rs_out<1> , \rs_out<0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33;

  lshifter ls ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Rot_sel(n1), .Out({\ls_out<15> , \ls_out<14> , 
        \ls_out<13> , \ls_out<12> , \ls_out<11> , \ls_out<10> , \ls_out<9> , 
        \ls_out<8> , \ls_out<7> , \ls_out<6> , \ls_out<5> , \ls_out<4> , 
        \ls_out<3> , \ls_out<2> , \ls_out<1> , \ls_out<0> }) );
  rshifter rs ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Rot_sel(n1), .Out({\rs_out<15> , \rs_out<14> , 
        \rs_out<13> , \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> , 
        \rs_out<8> , \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> , 
        \rs_out<3> , \rs_out<2> , \rs_out<1> , \rs_out<0> }) );
  INVX1 U1 ( .A(\rs_out<1> ), .Y(n4) );
  INVX1 U2 ( .A(\rs_out<3> ), .Y(n8) );
  INVX1 U3 ( .A(\rs_out<4> ), .Y(n10) );
  INVX1 U4 ( .A(\rs_out<9> ), .Y(n20) );
  INVX1 U5 ( .A(\rs_out<10> ), .Y(n22) );
  INVX1 U6 ( .A(\rs_out<11> ), .Y(n24) );
  INVX1 U7 ( .A(\rs_out<13> ), .Y(n28) );
  INVX1 U8 ( .A(\rs_out<14> ), .Y(n30) );
  INVX1 U9 ( .A(\rs_out<15> ), .Y(n32) );
  INVX1 U10 ( .A(\ls_out<4> ), .Y(n11) );
  INVX1 U11 ( .A(\ls_out<6> ), .Y(n15) );
  INVX1 U12 ( .A(\ls_out<9> ), .Y(n21) );
  INVX1 U13 ( .A(\ls_out<10> ), .Y(n23) );
  INVX1 U14 ( .A(\ls_out<13> ), .Y(n29) );
  INVX1 U15 ( .A(\ls_out<14> ), .Y(n31) );
  INVX1 U16 ( .A(\rs_out<0> ), .Y(n2) );
  INVX1 U17 ( .A(\rs_out<6> ), .Y(n14) );
  INVX1 U18 ( .A(\rs_out<7> ), .Y(n16) );
  INVX1 U19 ( .A(\rs_out<8> ), .Y(n18) );
  INVX1 U20 ( .A(\rs_out<12> ), .Y(n26) );
  INVX1 U21 ( .A(\ls_out<0> ), .Y(n3) );
  INVX1 U22 ( .A(\ls_out<1> ), .Y(n5) );
  INVX1 U23 ( .A(\ls_out<3> ), .Y(n9) );
  INVX1 U24 ( .A(\ls_out<7> ), .Y(n17) );
  INVX1 U25 ( .A(\ls_out<8> ), .Y(n19) );
  INVX1 U26 ( .A(\ls_out<11> ), .Y(n25) );
  INVX1 U27 ( .A(\ls_out<12> ), .Y(n27) );
  INVX1 U28 ( .A(\ls_out<15> ), .Y(n33) );
  INVX1 U29 ( .A(\ls_out<2> ), .Y(n7) );
  INVX1 U30 ( .A(\rs_out<5> ), .Y(n12) );
  INVX1 U31 ( .A(\ls_out<5> ), .Y(n13) );
  INVX1 U32 ( .A(\rs_out<2> ), .Y(n6) );
  INVX1 U33 ( .A(\Op<0> ), .Y(n1) );
  MUX2X1 U34 ( .B(n3), .A(n2), .S(\Op<1> ), .Y(\Out<0> ) );
  MUX2X1 U35 ( .B(n5), .A(n4), .S(\Op<1> ), .Y(\Out<1> ) );
  MUX2X1 U36 ( .B(n7), .A(n6), .S(\Op<1> ), .Y(\Out<2> ) );
  MUX2X1 U37 ( .B(n9), .A(n8), .S(\Op<1> ), .Y(\Out<3> ) );
  MUX2X1 U38 ( .B(n11), .A(n10), .S(\Op<1> ), .Y(\Out<4> ) );
  MUX2X1 U39 ( .B(n13), .A(n12), .S(\Op<1> ), .Y(\Out<5> ) );
  MUX2X1 U40 ( .B(n15), .A(n14), .S(\Op<1> ), .Y(\Out<6> ) );
  MUX2X1 U41 ( .B(n17), .A(n16), .S(\Op<1> ), .Y(\Out<7> ) );
  MUX2X1 U42 ( .B(n19), .A(n18), .S(\Op<1> ), .Y(\Out<8> ) );
  MUX2X1 U43 ( .B(n21), .A(n20), .S(\Op<1> ), .Y(\Out<9> ) );
  MUX2X1 U44 ( .B(n23), .A(n22), .S(\Op<1> ), .Y(\Out<10> ) );
  MUX2X1 U45 ( .B(n25), .A(n24), .S(\Op<1> ), .Y(\Out<11> ) );
  MUX2X1 U46 ( .B(n27), .A(n26), .S(\Op<1> ), .Y(\Out<12> ) );
  MUX2X1 U47 ( .B(n29), .A(n28), .S(\Op<1> ), .Y(\Out<13> ) );
  MUX2X1 U48 ( .B(n31), .A(n30), .S(\Op<1> ), .Y(\Out<14> ) );
  MUX2X1 U49 ( .B(n33), .A(n32), .S(\Op<1> ), .Y(\Out<15> ) );
endmodule


module cla4_7 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n22) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n24) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n26) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n28) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n30) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n32) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n34) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n36) );
  NOR3X1 U8 ( .A(n7), .B(n19), .C(n21), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n21), .C(n20), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n18), .C(\G<2> ), .Y(n41) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n40) );
  OAI21X1 U13 ( .A(n9), .B(n21), .C(n20), .Y(Cout) );
  AOI21X1 U14 ( .A(n16), .B(\P<2> ), .C(\G<2> ), .Y(n39) );
  AOI21X1 U15 ( .A(n12), .B(\P<1> ), .C(\G<1> ), .Y(n38) );
  fulladder1_31 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n31), .G(n23) );
  fulladder1_30 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n12), .S(\S<1> ), .P(
        n33), .G(n25) );
  fulladder1_29 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n16), .S(\S<2> ), .P(
        n35), .G(n27) );
  fulladder1_28 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n37), .G(n29) );
  INVX1 U1 ( .A(\P<2> ), .Y(n19) );
  AND2X1 U2 ( .A(n17), .B(n2), .Y(n10) );
  INVX1 U3 ( .A(\G<0> ), .Y(n17) );
  INVX1 U4 ( .A(\G<3> ), .Y(n20) );
  INVX1 U5 ( .A(\P<3> ), .Y(n21) );
  AND2X1 U6 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  BUFX2 U9 ( .A(n38), .Y(n3) );
  INVX1 U16 ( .A(n3), .Y(n16) );
  INVX1 U17 ( .A(n41), .Y(n4) );
  INVX1 U18 ( .A(n4), .Y(n5) );
  INVX1 U19 ( .A(n40), .Y(n18) );
  AND2X1 U20 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U21 ( .A(n6), .Y(n7) );
  INVX1 U22 ( .A(n9), .Y(n8) );
  BUFX2 U23 ( .A(n39), .Y(n9) );
  INVX1 U24 ( .A(n10), .Y(n12) );
  AND2X1 U25 ( .A(n36), .B(n37), .Y(\P<3> ) );
  AND2X1 U26 ( .A(n34), .B(n35), .Y(\P<2> ) );
  AND2X1 U27 ( .A(n32), .B(n33), .Y(\P<1> ) );
  AND2X1 U28 ( .A(n30), .B(n31), .Y(\P<0> ) );
  AND2X1 U29 ( .A(n28), .B(n29), .Y(\G<3> ) );
  AND2X1 U30 ( .A(n26), .B(n27), .Y(\G<2> ) );
  AND2X1 U31 ( .A(n24), .B(n25), .Y(\G<1> ) );
  AND2X1 U32 ( .A(n22), .B(n23), .Y(\G<0> ) );
endmodule


module cla4_6 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n7), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n9), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_27 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_26 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_25 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_24 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n38), .G(n30) );
  INVX1 U1 ( .A(\P<2> ), .Y(n20) );
  INVX1 U2 ( .A(\G<3> ), .Y(n21) );
  INVX1 U3 ( .A(\P<3> ), .Y(n22) );
  AND2X1 U4 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  BUFX2 U6 ( .A(n39), .Y(n3) );
  INVX1 U7 ( .A(n3), .Y(n17) );
  BUFX2 U9 ( .A(n41), .Y(n4) );
  INVX1 U16 ( .A(n4), .Y(n19) );
  BUFX2 U17 ( .A(n42), .Y(n5) );
  AND2X1 U18 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U19 ( .A(n6), .Y(n7) );
  INVX1 U20 ( .A(n10), .Y(n8) );
  INVX1 U21 ( .A(n8), .Y(n9) );
  BUFX2 U22 ( .A(n40), .Y(n10) );
  AND2X2 U23 ( .A(n18), .B(n2), .Y(n12) );
  INVX1 U24 ( .A(n12), .Y(n16) );
  AND2X1 U25 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U26 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U27 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U28 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U29 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U30 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U31 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U32 ( .A(n23), .B(n24), .Y(\G<0> ) );
  INVX2 U33 ( .A(\G<0> ), .Y(n18) );
endmodule


module cla4_5 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n23) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n25) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n27) );
  AND2X2 C24 ( .A(\A<3> ), .B(\B<3> ), .Y(n29) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n31) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n33) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n35) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n37) );
  NOR3X1 U8 ( .A(n7), .B(n20), .C(n22), .Y(PG) );
  OAI21X1 U10 ( .A(n5), .B(n22), .C(n21), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n19), .C(\G<2> ), .Y(n42) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n41) );
  OAI21X1 U13 ( .A(n9), .B(n22), .C(n21), .Y(Cout) );
  AOI21X1 U14 ( .A(n17), .B(\P<2> ), .C(\G<2> ), .Y(n40) );
  AOI21X1 U15 ( .A(n16), .B(\P<1> ), .C(\G<1> ), .Y(n39) );
  fulladder1_23 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n32), .G(n24) );
  fulladder1_22 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n16), .S(\S<1> ), .P(
        n34), .G(n26) );
  fulladder1_21 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n17), .S(\S<2> ), .P(
        n36), .G(n28) );
  fulladder1_20 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n8), .S(\S<3> ), .P(n38), .G(n30) );
  INVX1 U1 ( .A(\G<0> ), .Y(n18) );
  INVX1 U2 ( .A(\P<2> ), .Y(n20) );
  INVX1 U3 ( .A(\G<3> ), .Y(n21) );
  INVX1 U4 ( .A(\P<3> ), .Y(n22) );
  AND2X2 U5 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
  BUFX2 U7 ( .A(n39), .Y(n3) );
  INVX1 U9 ( .A(n3), .Y(n17) );
  BUFX2 U16 ( .A(n41), .Y(n4) );
  INVX1 U17 ( .A(n4), .Y(n19) );
  BUFX2 U18 ( .A(n42), .Y(n5) );
  AND2X1 U19 ( .A(\P<1> ), .B(\P<0> ), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(n7) );
  INVX1 U21 ( .A(n10), .Y(n8) );
  INVX1 U22 ( .A(n8), .Y(n9) );
  BUFX2 U23 ( .A(n40), .Y(n10) );
  AND2X2 U24 ( .A(n18), .B(n2), .Y(n12) );
  INVX1 U25 ( .A(n12), .Y(n16) );
  AND2X1 U26 ( .A(n37), .B(n38), .Y(\P<3> ) );
  AND2X1 U27 ( .A(n35), .B(n36), .Y(\P<2> ) );
  AND2X1 U28 ( .A(n33), .B(n34), .Y(\P<1> ) );
  AND2X1 U29 ( .A(n31), .B(n32), .Y(\P<0> ) );
  AND2X1 U30 ( .A(n29), .B(n30), .Y(\G<3> ) );
  AND2X1 U31 ( .A(n27), .B(n28), .Y(\G<2> ) );
  AND2X1 U32 ( .A(n25), .B(n26), .Y(\G<1> ) );
  AND2X1 U33 ( .A(n23), .B(n24), .Y(\G<0> ) );
endmodule


module cla4_4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, .S({\S<3> , \S<2> , \S<1> , \S<0> }), Cout, PG, 
        GG );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<3> , \S<2> , \S<1> , \S<0> , Cout, PG, GG;
  wire   \P<3> , \P<2> , \P<1> , \P<0> , \G<3> , \G<2> , \G<1> , \G<0> , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  AND2X2 C27 ( .A(\A<0> ), .B(\B<0> ), .Y(n21) );
  AND2X2 C26 ( .A(\A<1> ), .B(\B<1> ), .Y(n23) );
  AND2X2 C25 ( .A(\A<2> ), .B(\B<2> ), .Y(n25) );
  XOR2X1 C23 ( .A(\A<0> ), .B(\B<0> ), .Y(n29) );
  XOR2X1 C22 ( .A(\A<1> ), .B(\B<1> ), .Y(n31) );
  XOR2X1 C21 ( .A(\A<2> ), .B(\B<2> ), .Y(n33) );
  XOR2X1 C20 ( .A(\A<3> ), .B(\B<3> ), .Y(n35) );
  NOR3X1 U8 ( .A(n6), .B(n18), .C(n20), .Y(PG) );
  OAI21X1 U10 ( .A(n4), .B(n20), .C(n19), .Y(GG) );
  AOI21X1 U11 ( .A(\P<2> ), .B(n17), .C(\G<2> ), .Y(n40) );
  AOI21X1 U12 ( .A(\P<1> ), .B(\G<0> ), .C(\G<1> ), .Y(n39) );
  OAI21X1 U13 ( .A(n8), .B(n20), .C(n19), .Y(Cout) );
  AOI21X1 U14 ( .A(n12), .B(\P<2> ), .C(\G<2> ), .Y(n38) );
  AOI21X1 U15 ( .A(n10), .B(\P<1> ), .C(\G<1> ), .Y(n37) );
  fulladder1_19 \fa[0]  ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .S(\S<0> ), .P(
        n30), .G(n22) );
  fulladder1_18 \fa[1]  ( .A(\A<1> ), .B(\B<1> ), .Cin(n10), .S(\S<1> ), .P(
        n32), .G(n24) );
  fulladder1_17 \fa[2]  ( .A(\A<2> ), .B(\B<2> ), .Cin(n12), .S(\S<2> ), .P(
        n34), .G(n26) );
  fulladder1_16 \fa[3]  ( .A(\A<3> ), .B(\B<3> ), .Cin(n7), .S(\S<3> ), .P(n36), .G(n28) );
  AND2X1 U1 ( .A(Cin), .B(\P<0> ), .Y(n1) );
  INVX1 U2 ( .A(\P<2> ), .Y(n18) );
  INVX1 U3 ( .A(\G<3> ), .Y(n19) );
  AND2X1 U4 ( .A(\A<3> ), .B(\B<3> ), .Y(n27) );
  INVX1 U5 ( .A(\P<3> ), .Y(n20) );
  INVX1 U6 ( .A(n37), .Y(n12) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  BUFX2 U9 ( .A(n39), .Y(n3) );
  INVX1 U16 ( .A(n3), .Y(n17) );
  BUFX2 U17 ( .A(n40), .Y(n4) );
  AND2X1 U18 ( .A(\P<1> ), .B(\P<0> ), .Y(n5) );
  INVX1 U19 ( .A(n5), .Y(n6) );
  INVX1 U20 ( .A(n38), .Y(n7) );
  INVX1 U21 ( .A(n7), .Y(n8) );
  AND2X2 U22 ( .A(n2), .B(n16), .Y(n9) );
  INVX1 U23 ( .A(n9), .Y(n10) );
  AND2X1 U24 ( .A(n35), .B(n36), .Y(\P<3> ) );
  AND2X1 U25 ( .A(n33), .B(n34), .Y(\P<2> ) );
  AND2X1 U26 ( .A(n31), .B(n32), .Y(\P<1> ) );
  AND2X1 U27 ( .A(n29), .B(n30), .Y(\P<0> ) );
  AND2X1 U28 ( .A(n27), .B(n28), .Y(\G<3> ) );
  AND2X1 U29 ( .A(n25), .B(n26), .Y(\G<2> ) );
  AND2X1 U30 ( .A(n23), .B(n24), .Y(\G<1> ) );
  AND2X1 U31 ( .A(n21), .B(n22), .Y(\G<0> ) );
  INVX2 U32 ( .A(\G<0> ), .Y(n16) );
endmodule


module dff_388 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_389 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_390 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_391 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_392 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_393 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_394 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_395 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_396 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_397 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_398 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_399 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_400 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_401 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_402 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_403 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_372 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_373 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_374 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_375 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_376 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_377 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_378 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_379 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_380 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_381 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_382 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_383 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_384 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_385 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_386 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_387 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_404 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memory2c_1 ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, \mem<0><7> , \mem<0><6> , \mem<0><5> ,
         \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> ,
         \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> ,
         \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> ,
         \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> ,
         \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> ,
         \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> ,
         \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> ,
         \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> ,
         \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> ,
         \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> ,
         \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> ,
         \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> ,
         \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> ,
         \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> ,
         \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> ,
         \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> ,
         \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> ,
         \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> ,
         \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> ,
         \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> ,
         \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> ,
         \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> ,
         \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> ,
         \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> ,
         \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> ,
         \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> ,
         \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> ,
         \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> ,
         \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> ,
         \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> ,
         \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> ,
         \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> ,
         \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> ,
         \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> ,
         \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> ,
         \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> ,
         \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> ,
         \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> ,
         \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> , \mem<33><4> ,
         \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> , \mem<34><7> ,
         \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> , \mem<34><2> ,
         \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> , \mem<35><5> ,
         \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> , \mem<35><0> ,
         \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> , \mem<36><3> ,
         \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> , \mem<37><6> ,
         \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> , \mem<37><1> ,
         \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> , \mem<38><4> ,
         \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> , \mem<39><7> ,
         \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> , \mem<39><2> ,
         \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> , \mem<40><5> ,
         \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> , \mem<40><0> ,
         \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> , \mem<41><3> ,
         \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> , \mem<42><6> ,
         \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> , \mem<42><1> ,
         \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> , \mem<43><4> ,
         \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> , \mem<44><7> ,
         \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> , \mem<44><2> ,
         \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> , \mem<45><5> ,
         \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> , \mem<45><0> ,
         \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> , \mem<46><3> ,
         \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> , \mem<47><6> ,
         \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> , \mem<47><1> ,
         \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> , \mem<48><4> ,
         \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> , \mem<49><7> ,
         \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> , \mem<49><2> ,
         \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> , \mem<50><5> ,
         \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> , \mem<50><0> ,
         \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> , \mem<51><3> ,
         \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> , \mem<52><6> ,
         \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> , \mem<52><1> ,
         \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> , \mem<53><4> ,
         \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> , \mem<54><7> ,
         \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> , \mem<54><2> ,
         \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> , \mem<55><5> ,
         \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> , \mem<55><0> ,
         \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> , \mem<56><3> ,
         \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> , \mem<57><6> ,
         \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> , \mem<57><1> ,
         \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> , \mem<58><4> ,
         \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> , \mem<59><7> ,
         \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> , \mem<59><2> ,
         \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> , \mem<60><5> ,
         \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> , \mem<60><0> ,
         \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> , \mem<61><3> ,
         \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> , \mem<62><6> ,
         \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> , \mem<62><1> ,
         \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> , \mem<63><4> ,
         \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> , N185, N186,
         N187, N188, N189, N190, N191, N192, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n610, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1367, n1368,
         n1370, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1772, n1774, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1797,
         n1798, n1799, n1800, n1801, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n609, n611, n624, n637, n649, n661, n673, n685, n697,
         n709, n721, n733, n745, n757, n769, n781, n793, n805, n817, n829,
         n841, n853, n865, n877, n889, n901, n913, n925, n937, n949, n961,
         n973, n985, n997, n1009, n1021, n1033, n1045, n1057, n1069, n1081,
         n1093, n1105, n1117, n1129, n1141, n1153, n1165, n1177, n1189, n1201,
         n1213, n1225, n1237, n1249, n1261, n1273, n1285, n1297, n1309, n1321,
         n1333, n1345, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1369, n1371, n1372, n1383, n1384, n1396, n1397, n1409,
         n1410, n1424, n1425, n1436, n1437, n1449, n1450, n1461, n1462, n1476,
         n1477, n1488, n1489, n1501, n1502, n1513, n1514, n1528, n1529, n1540,
         n1541, n1553, n1554, n1565, n1566, n1580, n1581, n1592, n1593, n1605,
         n1606, n1617, n1618, n1632, n1633, n1644, n1645, n1657, n1658, n1669,
         n1670, n1684, n1685, n1696, n1697, n1709, n1710, n1721, n1722, n1736,
         n1737, n1758, n1759, n1771, n1773, n1775, n1776, n1793, n1794, n1795,
         n1796, n1802, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n2327), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2326), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2325), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2324), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2323), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2322), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2321), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2320), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2319), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2318), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2317), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2316), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2315), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2314), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2313), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2312), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2311), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2310), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2309), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2308), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2307), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2306), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2305), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2304), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2303), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2302), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2301), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2300), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2299), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2298), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2297), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2296), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2295), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2294), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2293), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2292), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2291), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2290), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2289), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2288), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2287), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2286), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2285), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2284), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2283), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2282), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2281), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2280), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2279), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2278), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2277), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2276), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2275), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2274), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2273), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2272), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2271), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2270), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2269), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2268), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2267), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2266), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2265), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2264), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2263), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2262), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2261), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2260), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2259), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2258), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2257), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2256), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2255), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2254), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2253), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2252), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2251), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2250), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2249), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2248), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2247), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2246), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2245), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2244), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2243), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2242), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2241), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2240), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2239), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2238), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2237), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2236), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2235), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2234), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2233), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2232), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2231), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2230), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2229), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2228), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2227), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2226), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2225), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2224), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2223), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2222), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2221), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2220), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2219), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2218), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2217), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2216), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2215), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2214), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2213), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2212), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2211), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2210), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2209), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2208), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2207), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2206), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2205), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2204), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2203), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2202), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2201), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2200), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2199), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2198), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2197), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2196), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2195), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2194), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2193), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2192), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2191), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2190), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2189), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2188), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2187), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2186), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2185), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2184), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2183), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2182), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2181), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2180), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2179), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2178), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2177), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2176), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2175), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2174), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2173), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2172), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2171), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2170), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2169), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2168), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2167), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2166), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2165), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2164), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2163), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2162), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2161), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2160), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2159), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2158), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2157), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2156), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2155), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2154), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2153), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2152), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2151), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2150), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2149), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2148), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2147), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2146), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2145), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2144), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2143), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2142), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2141), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2140), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2139), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2138), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2137), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2136), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2135), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2134), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2133), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2132), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2131), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2130), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2129), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2128), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2127), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2126), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2125), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2124), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2123), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2122), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2121), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2120), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2119), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2118), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2117), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2116), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2115), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2114), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2113), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2112), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2111), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2110), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2109), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2108), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2107), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2106), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2105), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2104), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2103), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2102), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2101), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2100), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2099), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2098), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2097), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2096), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2095), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2094), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2093), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2092), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2091), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2090), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2089), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2088), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2087), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2086), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2085), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2084), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2083), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2082), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2081), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2080), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2079), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2078), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2077), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2076), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2075), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2074), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2073), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2072), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n2071), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n2070), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n2069), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n2068), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n2067), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n2066), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n2065), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n2064), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n2063), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n2062), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n2061), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n2060), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n2059), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n2058), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n2057), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n2056), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n2055), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n2054), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n2053), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n2052), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n2051), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n2050), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n2049), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n2048), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n2047), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n2046), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n2045), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n2044), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n2043), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n2042), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n2041), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n2040), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n2039), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n2038), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n2037), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n2036), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n2035), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n2034), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n2033), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n2032), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n2031), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n2030), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n2029), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n2028), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n2027), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n2026), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n2025), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n2024), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n2023), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n2022), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n2021), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n2020), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n2019), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n2018), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n2017), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n2016), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n2015), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n2014), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n2013), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n2012), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n2011), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n2010), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n2009), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n2008), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n2007), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n2006), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n2005), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n2004), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n2003), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n2002), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n2001), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n2000), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n1999), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n1998), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n1997), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n1996), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n1995), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n1994), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n1993), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n1992), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n1991), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n1990), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n1989), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n1988), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n1987), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n1986), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n1985), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n1984), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n1983), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n1982), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n1981), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n1980), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n1979), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n1978), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n1977), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n1976), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n1975), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n1974), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n1973), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n1972), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n1971), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n1970), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n1969), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n1968), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n1967), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n1966), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n1965), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n1964), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n1963), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n1962), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n1961), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n1960), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n1959), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n1958), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n1957), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n1956), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n1955), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n1954), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n1953), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n1952), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n1951), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n1950), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n1949), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n1948), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n1947), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n1946), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n1945), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n1944), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n1943), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n1942), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n1941), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n1940), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n1939), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n1938), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n1937), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n1936), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n1935), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n1934), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n1933), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n1932), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n1931), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n1930), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n1929), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n1928), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n1927), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n1926), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n1925), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n1924), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n1923), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n1922), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n1921), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n1920), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n1919), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n1918), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n1917), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n1916), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n1915), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n1914), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n1913), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n1912), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n1911), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n1910), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n1909), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n1908), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n1907), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n1906), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n1905), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n1904), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n1903), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n1902), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n1901), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n1900), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n1899), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n1898), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n1897), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n1896), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n1895), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n1894), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n1893), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n1892), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n1891), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n1890), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n1889), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n1888), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n1887), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n1886), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n1885), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n1884), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n1883), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n1882), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n1881), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n1880), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n1879), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n1878), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n1877), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n1876), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n1875), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n1874), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n1873), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n1872), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n1871), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n1870), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n1869), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n1868), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n1867), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n1866), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n1865), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n1864), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n1863), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n1862), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n1861), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n1860), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n1859), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n1858), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n1857), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n1856), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n1855), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n1854), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n1853), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n1852), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n1851), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n1850), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n1849), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n1848), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n1847), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n1846), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n1845), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n1844), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n1843), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n1842), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n1841), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n1840), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n1839), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n1838), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n1837), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n1836), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n1835), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n1834), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n1833), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n1832), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n1831), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n1830), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n1829), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n1828), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n1827), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n1826), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n1825), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n1824), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n1823), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n1822), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n1821), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n1820), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n1819), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n1818), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n1817), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n1816), .CLK(clk), .Q(\mem<63><0> ) );
  AND2X2 U132 ( .A(n1376), .B(n1377), .Y(n1375) );
  AND2X2 U133 ( .A(n1381), .B(n1382), .Y(n1380) );
  AND2X2 U135 ( .A(n1388), .B(n1389), .Y(n1387) );
  AND2X2 U136 ( .A(n1393), .B(n1394), .Y(n1392) );
  AND2X2 U137 ( .A(n1401), .B(n1402), .Y(n1400) );
  AND2X2 U138 ( .A(n1407), .B(n1408), .Y(n1406) );
  AND2X2 U140 ( .A(n1414), .B(n1415), .Y(n1413) );
  AND2X2 U141 ( .A(n1419), .B(n1420), .Y(n1418) );
  AND2X2 U142 ( .A(n1429), .B(n1430), .Y(n1428) );
  AND2X2 U143 ( .A(n1434), .B(n1435), .Y(n1433) );
  AND2X2 U145 ( .A(n1441), .B(n1442), .Y(n1440) );
  AND2X2 U146 ( .A(n1446), .B(n1447), .Y(n1445) );
  AND2X2 U147 ( .A(n1454), .B(n1455), .Y(n1453) );
  AND2X2 U148 ( .A(n1459), .B(n1460), .Y(n1458) );
  AND2X2 U150 ( .A(n1466), .B(n1467), .Y(n1465) );
  AND2X2 U151 ( .A(n1471), .B(n1472), .Y(n1470) );
  AND2X2 U152 ( .A(n1481), .B(n1482), .Y(n1480) );
  AND2X2 U153 ( .A(n1486), .B(n1487), .Y(n1485) );
  AND2X2 U155 ( .A(n1493), .B(n1494), .Y(n1492) );
  AND2X2 U156 ( .A(n1498), .B(n1499), .Y(n1497) );
  AND2X2 U157 ( .A(n1506), .B(n1507), .Y(n1505) );
  AND2X2 U158 ( .A(n1511), .B(n1512), .Y(n1510) );
  AND2X2 U160 ( .A(n1518), .B(n1519), .Y(n1517) );
  AND2X2 U161 ( .A(n1523), .B(n1524), .Y(n1522) );
  AND2X2 U162 ( .A(n1533), .B(n1534), .Y(n1532) );
  AND2X2 U163 ( .A(n1538), .B(n1539), .Y(n1537) );
  AND2X2 U165 ( .A(n1545), .B(n1546), .Y(n1544) );
  AND2X2 U166 ( .A(n1550), .B(n1551), .Y(n1549) );
  AND2X2 U167 ( .A(n1558), .B(n1559), .Y(n1557) );
  AND2X2 U168 ( .A(n1563), .B(n1564), .Y(n1562) );
  AND2X2 U170 ( .A(n1570), .B(n1571), .Y(n1569) );
  AND2X2 U171 ( .A(n1575), .B(n1576), .Y(n1574) );
  AND2X2 U172 ( .A(n1585), .B(n1586), .Y(n1584) );
  AND2X2 U173 ( .A(n1590), .B(n1591), .Y(n1589) );
  AND2X2 U175 ( .A(n1597), .B(n1598), .Y(n1596) );
  AND2X2 U176 ( .A(n1602), .B(n1603), .Y(n1601) );
  AND2X2 U177 ( .A(n1610), .B(n1611), .Y(n1609) );
  AND2X2 U178 ( .A(n1615), .B(n1616), .Y(n1614) );
  AND2X2 U180 ( .A(n1622), .B(n1623), .Y(n1621) );
  AND2X2 U181 ( .A(n1627), .B(n1628), .Y(n1626) );
  AND2X2 U182 ( .A(n1637), .B(n1638), .Y(n1636) );
  AND2X2 U183 ( .A(n1642), .B(n1643), .Y(n1641) );
  AND2X2 U185 ( .A(n1649), .B(n1650), .Y(n1648) );
  AND2X2 U186 ( .A(n1654), .B(n1655), .Y(n1653) );
  AND2X2 U187 ( .A(n1662), .B(n1663), .Y(n1661) );
  AND2X2 U188 ( .A(n1667), .B(n1668), .Y(n1666) );
  AND2X2 U190 ( .A(n1674), .B(n1675), .Y(n1673) );
  AND2X2 U191 ( .A(n1679), .B(n1680), .Y(n1678) );
  AND2X2 U192 ( .A(n1689), .B(n1690), .Y(n1688) );
  AND2X2 U193 ( .A(n1694), .B(n1695), .Y(n1693) );
  AND2X2 U195 ( .A(n1701), .B(n1702), .Y(n1700) );
  AND2X2 U196 ( .A(n1706), .B(n1707), .Y(n1705) );
  AND2X2 U197 ( .A(n1714), .B(n1715), .Y(n1713) );
  AND2X2 U198 ( .A(n1719), .B(n1720), .Y(n1718) );
  AND2X2 U200 ( .A(n1726), .B(n1727), .Y(n1725) );
  AND2X2 U201 ( .A(n1731), .B(n1732), .Y(n1730) );
  AND2X2 U208 ( .A(n1741), .B(n1742), .Y(n1740) );
  AND2X2 U209 ( .A(n1753), .B(n1754), .Y(n1752) );
  AND2X2 U212 ( .A(n1763), .B(n1764), .Y(n1762) );
  AND2X2 U213 ( .A(n1768), .B(n1769), .Y(n1767) );
  AND2X2 U214 ( .A(n1780), .B(n1781), .Y(n1779) );
  OR2X2 U215 ( .A(n1785), .B(n1786), .Y(n1784) );
  AND2X2 U216 ( .A(n1791), .B(n1792), .Y(n1790) );
  AND2X2 U218 ( .A(n1800), .B(n1801), .Y(n1799) );
  AND2X2 U219 ( .A(n1806), .B(n1807), .Y(n1805) );
  OAI21X1 U817 ( .A(n598), .B(n3707), .C(n1776), .Y(n1816) );
  AOI22X1 U818 ( .A(\data_in<8> ), .B(n600), .C(\data_in<0> ), .D(n601), .Y(
        n599) );
  OAI21X1 U819 ( .A(n598), .B(n3706), .C(n1775), .Y(n1817) );
  AOI22X1 U820 ( .A(\data_in<9> ), .B(n600), .C(\data_in<1> ), .D(n601), .Y(
        n602) );
  OAI21X1 U821 ( .A(n598), .B(n3705), .C(n1773), .Y(n1818) );
  AOI22X1 U822 ( .A(\data_in<10> ), .B(n600), .C(\data_in<2> ), .D(n601), .Y(
        n603) );
  OAI21X1 U823 ( .A(n598), .B(n3704), .C(n1771), .Y(n1819) );
  AOI22X1 U824 ( .A(\data_in<11> ), .B(n600), .C(\data_in<3> ), .D(n601), .Y(
        n604) );
  OAI21X1 U825 ( .A(n598), .B(n3703), .C(n1759), .Y(n1820) );
  AOI22X1 U826 ( .A(\data_in<12> ), .B(n600), .C(\data_in<4> ), .D(n601), .Y(
        n605) );
  OAI21X1 U827 ( .A(n598), .B(n3702), .C(n1758), .Y(n1821) );
  AOI22X1 U828 ( .A(\data_in<13> ), .B(n600), .C(\data_in<5> ), .D(n601), .Y(
        n606) );
  OAI21X1 U829 ( .A(n598), .B(n3701), .C(n1737), .Y(n1822) );
  AOI22X1 U830 ( .A(\data_in<14> ), .B(n600), .C(\data_in<6> ), .D(n601), .Y(
        n607) );
  OAI21X1 U831 ( .A(n598), .B(n3700), .C(n1736), .Y(n1823) );
  AOI22X1 U832 ( .A(\data_in<15> ), .B(n600), .C(\data_in<7> ), .D(n601), .Y(
        n608) );
  OAI21X1 U833 ( .A(n2454), .B(n612), .C(n2460), .Y(n610) );
  OAI21X1 U834 ( .A(n3174), .B(n3699), .C(n1722), .Y(n1824) );
  AOI22X1 U835 ( .A(n615), .B(\data_in<8> ), .C(n616), .D(\data_in<0> ), .Y(
        n614) );
  OAI21X1 U836 ( .A(n3174), .B(n3698), .C(n1721), .Y(n1825) );
  AOI22X1 U837 ( .A(n615), .B(\data_in<9> ), .C(n616), .D(\data_in<1> ), .Y(
        n617) );
  OAI21X1 U838 ( .A(n3174), .B(n3697), .C(n1710), .Y(n1826) );
  AOI22X1 U839 ( .A(n615), .B(\data_in<10> ), .C(n616), .D(\data_in<2> ), .Y(
        n618) );
  OAI21X1 U840 ( .A(n3174), .B(n3696), .C(n1709), .Y(n1827) );
  AOI22X1 U841 ( .A(n615), .B(\data_in<11> ), .C(n616), .D(\data_in<3> ), .Y(
        n619) );
  OAI21X1 U842 ( .A(n3174), .B(n3695), .C(n1697), .Y(n1828) );
  AOI22X1 U843 ( .A(n615), .B(\data_in<12> ), .C(n616), .D(\data_in<4> ), .Y(
        n620) );
  OAI21X1 U844 ( .A(n3174), .B(n3694), .C(n1696), .Y(n1829) );
  AOI22X1 U845 ( .A(n615), .B(\data_in<13> ), .C(n616), .D(\data_in<5> ), .Y(
        n621) );
  OAI21X1 U846 ( .A(n3174), .B(n3693), .C(n1685), .Y(n1830) );
  AOI22X1 U847 ( .A(n615), .B(\data_in<14> ), .C(n616), .D(\data_in<6> ), .Y(
        n622) );
  OAI21X1 U848 ( .A(n3174), .B(n3692), .C(n1684), .Y(n1831) );
  AOI22X1 U849 ( .A(n615), .B(\data_in<15> ), .C(n616), .D(\data_in<7> ), .Y(
        n623) );
  AOI21X1 U850 ( .A(n2460), .B(n2564), .C(n2452), .Y(n613) );
  OAI21X1 U851 ( .A(n3173), .B(n3691), .C(n1670), .Y(n1832) );
  AOI22X1 U852 ( .A(n628), .B(\data_in<8> ), .C(n629), .D(\data_in<0> ), .Y(
        n627) );
  OAI21X1 U853 ( .A(n3173), .B(n3690), .C(n1669), .Y(n1833) );
  AOI22X1 U854 ( .A(n628), .B(\data_in<9> ), .C(n629), .D(\data_in<1> ), .Y(
        n630) );
  OAI21X1 U855 ( .A(n3173), .B(n3689), .C(n1658), .Y(n1834) );
  AOI22X1 U856 ( .A(n628), .B(\data_in<10> ), .C(n629), .D(\data_in<2> ), .Y(
        n631) );
  OAI21X1 U857 ( .A(n3173), .B(n3688), .C(n1657), .Y(n1835) );
  AOI22X1 U858 ( .A(n628), .B(\data_in<11> ), .C(n629), .D(\data_in<3> ), .Y(
        n632) );
  OAI21X1 U859 ( .A(n3173), .B(n3687), .C(n1645), .Y(n1836) );
  AOI22X1 U860 ( .A(n628), .B(\data_in<12> ), .C(n629), .D(\data_in<4> ), .Y(
        n633) );
  OAI21X1 U861 ( .A(n3173), .B(n3686), .C(n1644), .Y(n1837) );
  AOI22X1 U862 ( .A(n628), .B(\data_in<13> ), .C(n629), .D(\data_in<5> ), .Y(
        n634) );
  OAI21X1 U863 ( .A(n3173), .B(n3685), .C(n1633), .Y(n1838) );
  AOI22X1 U864 ( .A(n628), .B(\data_in<14> ), .C(n629), .D(\data_in<6> ), .Y(
        n635) );
  OAI21X1 U865 ( .A(n3173), .B(n3684), .C(n1632), .Y(n1839) );
  AOI22X1 U866 ( .A(n628), .B(\data_in<15> ), .C(n629), .D(\data_in<7> ), .Y(
        n636) );
  AOI21X1 U867 ( .A(n2564), .B(n2560), .C(n2452), .Y(n626) );
  OAI21X1 U868 ( .A(n3172), .B(n3683), .C(n1618), .Y(n1840) );
  AOI22X1 U869 ( .A(n640), .B(\data_in<8> ), .C(n641), .D(\data_in<0> ), .Y(
        n639) );
  OAI21X1 U870 ( .A(n3172), .B(n3682), .C(n1617), .Y(n1841) );
  AOI22X1 U871 ( .A(n640), .B(\data_in<9> ), .C(n641), .D(\data_in<1> ), .Y(
        n642) );
  OAI21X1 U872 ( .A(n3172), .B(n3681), .C(n1606), .Y(n1842) );
  AOI22X1 U873 ( .A(n640), .B(\data_in<10> ), .C(n641), .D(\data_in<2> ), .Y(
        n643) );
  OAI21X1 U874 ( .A(n3172), .B(n3680), .C(n1605), .Y(n1843) );
  AOI22X1 U875 ( .A(n640), .B(\data_in<11> ), .C(n641), .D(\data_in<3> ), .Y(
        n644) );
  OAI21X1 U876 ( .A(n3172), .B(n3679), .C(n1593), .Y(n1844) );
  AOI22X1 U877 ( .A(n640), .B(\data_in<12> ), .C(n641), .D(\data_in<4> ), .Y(
        n645) );
  OAI21X1 U878 ( .A(n3172), .B(n3678), .C(n1592), .Y(n1845) );
  AOI22X1 U879 ( .A(n640), .B(\data_in<13> ), .C(n641), .D(\data_in<5> ), .Y(
        n646) );
  OAI21X1 U880 ( .A(n3172), .B(n3677), .C(n1581), .Y(n1846) );
  AOI22X1 U881 ( .A(n640), .B(\data_in<14> ), .C(n641), .D(\data_in<6> ), .Y(
        n647) );
  OAI21X1 U882 ( .A(n3172), .B(n3676), .C(n1580), .Y(n1847) );
  AOI22X1 U883 ( .A(n640), .B(\data_in<15> ), .C(n641), .D(\data_in<7> ), .Y(
        n648) );
  AOI21X1 U884 ( .A(n2560), .B(n2562), .C(n2452), .Y(n638) );
  OAI21X1 U885 ( .A(n3171), .B(n3675), .C(n1566), .Y(n1848) );
  AOI22X1 U886 ( .A(n652), .B(\data_in<8> ), .C(n653), .D(\data_in<0> ), .Y(
        n651) );
  OAI21X1 U887 ( .A(n3171), .B(n3674), .C(n1565), .Y(n1849) );
  AOI22X1 U888 ( .A(n652), .B(\data_in<9> ), .C(n653), .D(\data_in<1> ), .Y(
        n654) );
  OAI21X1 U889 ( .A(n3171), .B(n3673), .C(n1554), .Y(n1850) );
  AOI22X1 U890 ( .A(n652), .B(\data_in<10> ), .C(n653), .D(\data_in<2> ), .Y(
        n655) );
  OAI21X1 U891 ( .A(n3171), .B(n3672), .C(n1553), .Y(n1851) );
  AOI22X1 U892 ( .A(n652), .B(\data_in<11> ), .C(n653), .D(\data_in<3> ), .Y(
        n656) );
  OAI21X1 U893 ( .A(n3171), .B(n3671), .C(n1541), .Y(n1852) );
  AOI22X1 U894 ( .A(n652), .B(\data_in<12> ), .C(n653), .D(\data_in<4> ), .Y(
        n657) );
  OAI21X1 U895 ( .A(n3171), .B(n3670), .C(n1540), .Y(n1853) );
  AOI22X1 U896 ( .A(n652), .B(\data_in<13> ), .C(n653), .D(\data_in<5> ), .Y(
        n658) );
  OAI21X1 U897 ( .A(n3171), .B(n3669), .C(n1529), .Y(n1854) );
  AOI22X1 U898 ( .A(n652), .B(\data_in<14> ), .C(n653), .D(\data_in<6> ), .Y(
        n659) );
  OAI21X1 U899 ( .A(n3171), .B(n3668), .C(n1528), .Y(n1855) );
  AOI22X1 U900 ( .A(n652), .B(\data_in<15> ), .C(n653), .D(\data_in<7> ), .Y(
        n660) );
  AOI21X1 U901 ( .A(n2562), .B(n2556), .C(n2452), .Y(n650) );
  OAI21X1 U902 ( .A(n3170), .B(n3667), .C(n1514), .Y(n1856) );
  AOI22X1 U903 ( .A(n664), .B(\data_in<8> ), .C(n665), .D(\data_in<0> ), .Y(
        n663) );
  OAI21X1 U904 ( .A(n3170), .B(n3666), .C(n1513), .Y(n1857) );
  AOI22X1 U905 ( .A(n664), .B(\data_in<9> ), .C(n665), .D(\data_in<1> ), .Y(
        n666) );
  OAI21X1 U906 ( .A(n3170), .B(n3665), .C(n1502), .Y(n1858) );
  AOI22X1 U907 ( .A(n664), .B(\data_in<10> ), .C(n665), .D(\data_in<2> ), .Y(
        n667) );
  OAI21X1 U908 ( .A(n3170), .B(n3664), .C(n1501), .Y(n1859) );
  AOI22X1 U909 ( .A(n664), .B(\data_in<11> ), .C(n665), .D(\data_in<3> ), .Y(
        n668) );
  OAI21X1 U910 ( .A(n3170), .B(n3663), .C(n1489), .Y(n1860) );
  AOI22X1 U911 ( .A(n664), .B(\data_in<12> ), .C(n665), .D(\data_in<4> ), .Y(
        n669) );
  OAI21X1 U912 ( .A(n3170), .B(n3662), .C(n1488), .Y(n1861) );
  AOI22X1 U913 ( .A(n664), .B(\data_in<13> ), .C(n665), .D(\data_in<5> ), .Y(
        n670) );
  OAI21X1 U914 ( .A(n3170), .B(n3661), .C(n1477), .Y(n1862) );
  AOI22X1 U915 ( .A(n664), .B(\data_in<14> ), .C(n665), .D(\data_in<6> ), .Y(
        n671) );
  OAI21X1 U916 ( .A(n3170), .B(n3660), .C(n1476), .Y(n1863) );
  AOI22X1 U917 ( .A(n664), .B(\data_in<15> ), .C(n665), .D(\data_in<7> ), .Y(
        n672) );
  AOI21X1 U918 ( .A(n2556), .B(n2558), .C(n2452), .Y(n662) );
  OAI21X1 U919 ( .A(n3169), .B(n3659), .C(n1462), .Y(n1864) );
  AOI22X1 U920 ( .A(n676), .B(\data_in<8> ), .C(n677), .D(\data_in<0> ), .Y(
        n675) );
  OAI21X1 U921 ( .A(n3169), .B(n3658), .C(n1461), .Y(n1865) );
  AOI22X1 U922 ( .A(n676), .B(\data_in<9> ), .C(n677), .D(\data_in<1> ), .Y(
        n678) );
  OAI21X1 U923 ( .A(n3169), .B(n3657), .C(n1450), .Y(n1866) );
  AOI22X1 U924 ( .A(n676), .B(\data_in<10> ), .C(n677), .D(\data_in<2> ), .Y(
        n679) );
  OAI21X1 U925 ( .A(n3169), .B(n3656), .C(n1449), .Y(n1867) );
  AOI22X1 U926 ( .A(n676), .B(\data_in<11> ), .C(n677), .D(\data_in<3> ), .Y(
        n680) );
  OAI21X1 U927 ( .A(n3169), .B(n3655), .C(n1437), .Y(n1868) );
  AOI22X1 U928 ( .A(n676), .B(\data_in<12> ), .C(n677), .D(\data_in<4> ), .Y(
        n681) );
  OAI21X1 U929 ( .A(n3169), .B(n3654), .C(n1436), .Y(n1869) );
  AOI22X1 U930 ( .A(n676), .B(\data_in<13> ), .C(n677), .D(\data_in<5> ), .Y(
        n682) );
  OAI21X1 U931 ( .A(n3169), .B(n3653), .C(n1425), .Y(n1870) );
  AOI22X1 U932 ( .A(n676), .B(\data_in<14> ), .C(n677), .D(\data_in<6> ), .Y(
        n683) );
  OAI21X1 U933 ( .A(n3169), .B(n3652), .C(n1424), .Y(n1871) );
  AOI22X1 U934 ( .A(n676), .B(\data_in<15> ), .C(n677), .D(\data_in<7> ), .Y(
        n684) );
  AOI21X1 U935 ( .A(n2558), .B(n2552), .C(n2452), .Y(n674) );
  OAI21X1 U936 ( .A(n3168), .B(n3651), .C(n1410), .Y(n1872) );
  AOI22X1 U937 ( .A(n688), .B(\data_in<8> ), .C(n689), .D(\data_in<0> ), .Y(
        n687) );
  OAI21X1 U938 ( .A(n3168), .B(n3650), .C(n1409), .Y(n1873) );
  AOI22X1 U939 ( .A(n688), .B(\data_in<9> ), .C(n689), .D(\data_in<1> ), .Y(
        n690) );
  OAI21X1 U940 ( .A(n3168), .B(n3649), .C(n1397), .Y(n1874) );
  AOI22X1 U941 ( .A(n688), .B(\data_in<10> ), .C(n689), .D(\data_in<2> ), .Y(
        n691) );
  OAI21X1 U942 ( .A(n3168), .B(n3648), .C(n1396), .Y(n1875) );
  AOI22X1 U943 ( .A(n688), .B(\data_in<11> ), .C(n689), .D(\data_in<3> ), .Y(
        n692) );
  OAI21X1 U944 ( .A(n3168), .B(n3647), .C(n1384), .Y(n1876) );
  AOI22X1 U945 ( .A(n688), .B(\data_in<12> ), .C(n689), .D(\data_in<4> ), .Y(
        n693) );
  OAI21X1 U946 ( .A(n3168), .B(n3646), .C(n1383), .Y(n1877) );
  AOI22X1 U947 ( .A(n688), .B(\data_in<13> ), .C(n689), .D(\data_in<5> ), .Y(
        n694) );
  OAI21X1 U948 ( .A(n3168), .B(n3645), .C(n1372), .Y(n1878) );
  AOI22X1 U949 ( .A(n688), .B(\data_in<14> ), .C(n689), .D(\data_in<6> ), .Y(
        n695) );
  OAI21X1 U950 ( .A(n3168), .B(n3644), .C(n1371), .Y(n1879) );
  AOI22X1 U951 ( .A(n688), .B(\data_in<15> ), .C(n689), .D(\data_in<7> ), .Y(
        n696) );
  AOI21X1 U952 ( .A(n2552), .B(n2554), .C(n2452), .Y(n686) );
  OAI21X1 U953 ( .A(n3167), .B(n3643), .C(n1369), .Y(n1880) );
  AOI22X1 U954 ( .A(n700), .B(\data_in<8> ), .C(n701), .D(\data_in<0> ), .Y(
        n699) );
  OAI21X1 U955 ( .A(n3167), .B(n3642), .C(n1366), .Y(n1881) );
  AOI22X1 U956 ( .A(n700), .B(\data_in<9> ), .C(n701), .D(\data_in<1> ), .Y(
        n702) );
  OAI21X1 U957 ( .A(n3167), .B(n3641), .C(n1365), .Y(n1882) );
  AOI22X1 U958 ( .A(n700), .B(\data_in<10> ), .C(n701), .D(\data_in<2> ), .Y(
        n703) );
  OAI21X1 U959 ( .A(n3167), .B(n3640), .C(n1364), .Y(n1883) );
  AOI22X1 U960 ( .A(n700), .B(\data_in<11> ), .C(n701), .D(\data_in<3> ), .Y(
        n704) );
  OAI21X1 U961 ( .A(n3167), .B(n3639), .C(n1363), .Y(n1884) );
  AOI22X1 U962 ( .A(n700), .B(\data_in<12> ), .C(n701), .D(\data_in<4> ), .Y(
        n705) );
  OAI21X1 U963 ( .A(n3167), .B(n3638), .C(n1362), .Y(n1885) );
  AOI22X1 U964 ( .A(n700), .B(\data_in<13> ), .C(n701), .D(\data_in<5> ), .Y(
        n706) );
  OAI21X1 U965 ( .A(n3167), .B(n3637), .C(n1361), .Y(n1886) );
  AOI22X1 U966 ( .A(n700), .B(\data_in<14> ), .C(n701), .D(\data_in<6> ), .Y(
        n707) );
  OAI21X1 U967 ( .A(n3167), .B(n3636), .C(n1360), .Y(n1887) );
  AOI22X1 U968 ( .A(n700), .B(\data_in<15> ), .C(n701), .D(\data_in<7> ), .Y(
        n708) );
  AOI21X1 U969 ( .A(n2554), .B(n2578), .C(n2452), .Y(n698) );
  OAI21X1 U970 ( .A(n3166), .B(n3635), .C(n1359), .Y(n1888) );
  AOI22X1 U971 ( .A(n712), .B(\data_in<8> ), .C(n713), .D(\data_in<0> ), .Y(
        n711) );
  OAI21X1 U972 ( .A(n3166), .B(n3634), .C(n1358), .Y(n1889) );
  AOI22X1 U973 ( .A(n712), .B(\data_in<9> ), .C(n713), .D(\data_in<1> ), .Y(
        n714) );
  OAI21X1 U974 ( .A(n3166), .B(n3633), .C(n1357), .Y(n1890) );
  AOI22X1 U975 ( .A(n712), .B(\data_in<10> ), .C(n713), .D(\data_in<2> ), .Y(
        n715) );
  OAI21X1 U976 ( .A(n3166), .B(n3632), .C(n1345), .Y(n1891) );
  AOI22X1 U977 ( .A(n712), .B(\data_in<11> ), .C(n713), .D(\data_in<3> ), .Y(
        n716) );
  OAI21X1 U978 ( .A(n3166), .B(n3631), .C(n1333), .Y(n1892) );
  AOI22X1 U979 ( .A(n712), .B(\data_in<12> ), .C(n713), .D(\data_in<4> ), .Y(
        n717) );
  OAI21X1 U980 ( .A(n3166), .B(n3630), .C(n1321), .Y(n1893) );
  AOI22X1 U981 ( .A(n712), .B(\data_in<13> ), .C(n713), .D(\data_in<5> ), .Y(
        n718) );
  OAI21X1 U982 ( .A(n3166), .B(n3629), .C(n1309), .Y(n1894) );
  AOI22X1 U983 ( .A(n712), .B(\data_in<14> ), .C(n713), .D(\data_in<6> ), .Y(
        n719) );
  OAI21X1 U984 ( .A(n3166), .B(n3628), .C(n1297), .Y(n1895) );
  AOI22X1 U985 ( .A(n712), .B(\data_in<15> ), .C(n713), .D(\data_in<7> ), .Y(
        n720) );
  AOI21X1 U986 ( .A(n2578), .B(n2580), .C(n2452), .Y(n710) );
  OAI21X1 U987 ( .A(n3165), .B(n3627), .C(n1285), .Y(n1896) );
  AOI22X1 U988 ( .A(n724), .B(\data_in<8> ), .C(n725), .D(\data_in<0> ), .Y(
        n723) );
  OAI21X1 U989 ( .A(n3165), .B(n3626), .C(n1273), .Y(n1897) );
  AOI22X1 U990 ( .A(n724), .B(\data_in<9> ), .C(n725), .D(\data_in<1> ), .Y(
        n726) );
  OAI21X1 U991 ( .A(n3165), .B(n3625), .C(n1261), .Y(n1898) );
  AOI22X1 U992 ( .A(n724), .B(\data_in<10> ), .C(n725), .D(\data_in<2> ), .Y(
        n727) );
  OAI21X1 U993 ( .A(n3165), .B(n3624), .C(n1249), .Y(n1899) );
  AOI22X1 U994 ( .A(n724), .B(\data_in<11> ), .C(n725), .D(\data_in<3> ), .Y(
        n728) );
  OAI21X1 U995 ( .A(n3165), .B(n3623), .C(n1237), .Y(n1900) );
  AOI22X1 U996 ( .A(n724), .B(\data_in<12> ), .C(n725), .D(\data_in<4> ), .Y(
        n729) );
  OAI21X1 U997 ( .A(n3165), .B(n3622), .C(n1225), .Y(n1901) );
  AOI22X1 U998 ( .A(n724), .B(\data_in<13> ), .C(n725), .D(\data_in<5> ), .Y(
        n730) );
  OAI21X1 U999 ( .A(n3165), .B(n3621), .C(n1213), .Y(n1902) );
  AOI22X1 U1000 ( .A(n724), .B(\data_in<14> ), .C(n725), .D(\data_in<6> ), .Y(
        n731) );
  OAI21X1 U1001 ( .A(n3165), .B(n3620), .C(n1201), .Y(n1903) );
  AOI22X1 U1002 ( .A(n724), .B(\data_in<15> ), .C(n725), .D(\data_in<7> ), .Y(
        n732) );
  AOI21X1 U1003 ( .A(n2580), .B(n2574), .C(n2452), .Y(n722) );
  OAI21X1 U1004 ( .A(n3164), .B(n3619), .C(n1189), .Y(n1904) );
  AOI22X1 U1005 ( .A(n736), .B(\data_in<8> ), .C(n737), .D(\data_in<0> ), .Y(
        n735) );
  OAI21X1 U1006 ( .A(n3164), .B(n3618), .C(n1177), .Y(n1905) );
  AOI22X1 U1007 ( .A(n736), .B(\data_in<9> ), .C(n737), .D(\data_in<1> ), .Y(
        n738) );
  OAI21X1 U1008 ( .A(n3164), .B(n3617), .C(n1165), .Y(n1906) );
  AOI22X1 U1009 ( .A(n736), .B(\data_in<10> ), .C(n737), .D(\data_in<2> ), .Y(
        n739) );
  OAI21X1 U1010 ( .A(n3164), .B(n3616), .C(n1153), .Y(n1907) );
  AOI22X1 U1011 ( .A(n736), .B(\data_in<11> ), .C(n737), .D(\data_in<3> ), .Y(
        n740) );
  OAI21X1 U1012 ( .A(n3164), .B(n3615), .C(n1141), .Y(n1908) );
  AOI22X1 U1013 ( .A(n736), .B(\data_in<12> ), .C(n737), .D(\data_in<4> ), .Y(
        n741) );
  OAI21X1 U1014 ( .A(n3164), .B(n3614), .C(n1129), .Y(n1909) );
  AOI22X1 U1015 ( .A(n736), .B(\data_in<13> ), .C(n737), .D(\data_in<5> ), .Y(
        n742) );
  OAI21X1 U1016 ( .A(n3164), .B(n3613), .C(n1117), .Y(n1910) );
  AOI22X1 U1017 ( .A(n736), .B(\data_in<14> ), .C(n737), .D(\data_in<6> ), .Y(
        n743) );
  OAI21X1 U1018 ( .A(n3164), .B(n3612), .C(n1105), .Y(n1911) );
  AOI22X1 U1019 ( .A(n736), .B(\data_in<15> ), .C(n737), .D(\data_in<7> ), .Y(
        n744) );
  AOI21X1 U1020 ( .A(n2574), .B(n2576), .C(n2452), .Y(n734) );
  OAI21X1 U1021 ( .A(n3163), .B(n3611), .C(n1093), .Y(n1912) );
  AOI22X1 U1022 ( .A(n748), .B(\data_in<8> ), .C(n749), .D(\data_in<0> ), .Y(
        n747) );
  OAI21X1 U1023 ( .A(n3163), .B(n3610), .C(n1081), .Y(n1913) );
  AOI22X1 U1024 ( .A(n748), .B(\data_in<9> ), .C(n749), .D(\data_in<1> ), .Y(
        n750) );
  OAI21X1 U1025 ( .A(n3163), .B(n3609), .C(n1069), .Y(n1914) );
  AOI22X1 U1026 ( .A(n748), .B(\data_in<10> ), .C(n749), .D(\data_in<2> ), .Y(
        n751) );
  OAI21X1 U1027 ( .A(n3163), .B(n3608), .C(n1057), .Y(n1915) );
  AOI22X1 U1028 ( .A(n748), .B(\data_in<11> ), .C(n749), .D(\data_in<3> ), .Y(
        n752) );
  OAI21X1 U1029 ( .A(n3163), .B(n3607), .C(n1045), .Y(n1916) );
  AOI22X1 U1030 ( .A(n748), .B(\data_in<12> ), .C(n749), .D(\data_in<4> ), .Y(
        n753) );
  OAI21X1 U1031 ( .A(n3163), .B(n3606), .C(n1033), .Y(n1917) );
  AOI22X1 U1032 ( .A(n748), .B(\data_in<13> ), .C(n749), .D(\data_in<5> ), .Y(
        n754) );
  OAI21X1 U1033 ( .A(n3163), .B(n3605), .C(n1021), .Y(n1918) );
  AOI22X1 U1034 ( .A(n748), .B(\data_in<14> ), .C(n749), .D(\data_in<6> ), .Y(
        n755) );
  OAI21X1 U1035 ( .A(n3163), .B(n3604), .C(n1009), .Y(n1919) );
  AOI22X1 U1036 ( .A(n748), .B(\data_in<15> ), .C(n749), .D(\data_in<7> ), .Y(
        n756) );
  AOI21X1 U1037 ( .A(n2576), .B(n2570), .C(n2452), .Y(n746) );
  OAI21X1 U1038 ( .A(n3162), .B(n3603), .C(n997), .Y(n1920) );
  AOI22X1 U1039 ( .A(n760), .B(\data_in<8> ), .C(n761), .D(\data_in<0> ), .Y(
        n759) );
  OAI21X1 U1040 ( .A(n3162), .B(n3602), .C(n985), .Y(n1921) );
  AOI22X1 U1041 ( .A(n760), .B(\data_in<9> ), .C(n761), .D(\data_in<1> ), .Y(
        n762) );
  OAI21X1 U1042 ( .A(n3162), .B(n3601), .C(n973), .Y(n1922) );
  AOI22X1 U1043 ( .A(n760), .B(\data_in<10> ), .C(n761), .D(\data_in<2> ), .Y(
        n763) );
  OAI21X1 U1044 ( .A(n3162), .B(n3600), .C(n961), .Y(n1923) );
  AOI22X1 U1045 ( .A(n760), .B(\data_in<11> ), .C(n761), .D(\data_in<3> ), .Y(
        n764) );
  OAI21X1 U1046 ( .A(n3162), .B(n3599), .C(n949), .Y(n1924) );
  AOI22X1 U1047 ( .A(n760), .B(\data_in<12> ), .C(n761), .D(\data_in<4> ), .Y(
        n765) );
  OAI21X1 U1048 ( .A(n3162), .B(n3598), .C(n937), .Y(n1925) );
  AOI22X1 U1049 ( .A(n760), .B(\data_in<13> ), .C(n761), .D(\data_in<5> ), .Y(
        n766) );
  OAI21X1 U1050 ( .A(n3162), .B(n3597), .C(n925), .Y(n1926) );
  AOI22X1 U1051 ( .A(n760), .B(\data_in<14> ), .C(n761), .D(\data_in<6> ), .Y(
        n767) );
  OAI21X1 U1052 ( .A(n3162), .B(n3596), .C(n913), .Y(n1927) );
  AOI22X1 U1053 ( .A(n760), .B(\data_in<15> ), .C(n761), .D(\data_in<7> ), .Y(
        n768) );
  AOI21X1 U1054 ( .A(n2570), .B(n2572), .C(n2452), .Y(n758) );
  OAI21X1 U1055 ( .A(n3161), .B(n3595), .C(n901), .Y(n1928) );
  AOI22X1 U1056 ( .A(n772), .B(\data_in<8> ), .C(n773), .D(\data_in<0> ), .Y(
        n771) );
  OAI21X1 U1057 ( .A(n3161), .B(n3594), .C(n889), .Y(n1929) );
  AOI22X1 U1058 ( .A(n772), .B(\data_in<9> ), .C(n773), .D(\data_in<1> ), .Y(
        n774) );
  OAI21X1 U1059 ( .A(n3161), .B(n3593), .C(n877), .Y(n1930) );
  AOI22X1 U1060 ( .A(n772), .B(\data_in<10> ), .C(n773), .D(\data_in<2> ), .Y(
        n775) );
  OAI21X1 U1061 ( .A(n3161), .B(n3592), .C(n865), .Y(n1931) );
  AOI22X1 U1062 ( .A(n772), .B(\data_in<11> ), .C(n773), .D(\data_in<3> ), .Y(
        n776) );
  OAI21X1 U1063 ( .A(n3161), .B(n3591), .C(n853), .Y(n1932) );
  AOI22X1 U1064 ( .A(n772), .B(\data_in<12> ), .C(n773), .D(\data_in<4> ), .Y(
        n777) );
  OAI21X1 U1065 ( .A(n3161), .B(n3590), .C(n841), .Y(n1933) );
  AOI22X1 U1066 ( .A(n772), .B(\data_in<13> ), .C(n773), .D(\data_in<5> ), .Y(
        n778) );
  OAI21X1 U1067 ( .A(n3161), .B(n3589), .C(n829), .Y(n1934) );
  AOI22X1 U1068 ( .A(n772), .B(\data_in<14> ), .C(n773), .D(\data_in<6> ), .Y(
        n779) );
  OAI21X1 U1069 ( .A(n3161), .B(n3588), .C(n817), .Y(n1935) );
  AOI22X1 U1070 ( .A(n772), .B(\data_in<15> ), .C(n773), .D(\data_in<7> ), .Y(
        n780) );
  AOI21X1 U1071 ( .A(n2572), .B(n2566), .C(n2452), .Y(n770) );
  OAI21X1 U1072 ( .A(n3160), .B(n3587), .C(n805), .Y(n1936) );
  AOI22X1 U1073 ( .A(n784), .B(\data_in<8> ), .C(n785), .D(\data_in<0> ), .Y(
        n783) );
  OAI21X1 U1074 ( .A(n3160), .B(n3586), .C(n793), .Y(n1937) );
  AOI22X1 U1075 ( .A(n784), .B(\data_in<9> ), .C(n785), .D(\data_in<1> ), .Y(
        n786) );
  OAI21X1 U1076 ( .A(n3160), .B(n3585), .C(n781), .Y(n1938) );
  AOI22X1 U1077 ( .A(n784), .B(\data_in<10> ), .C(n785), .D(\data_in<2> ), .Y(
        n787) );
  OAI21X1 U1078 ( .A(n3160), .B(n3584), .C(n769), .Y(n1939) );
  AOI22X1 U1079 ( .A(n784), .B(\data_in<11> ), .C(n785), .D(\data_in<3> ), .Y(
        n788) );
  OAI21X1 U1080 ( .A(n3160), .B(n3583), .C(n757), .Y(n1940) );
  AOI22X1 U1081 ( .A(n784), .B(\data_in<12> ), .C(n785), .D(\data_in<4> ), .Y(
        n789) );
  OAI21X1 U1082 ( .A(n3160), .B(n3582), .C(n745), .Y(n1941) );
  AOI22X1 U1083 ( .A(n784), .B(\data_in<13> ), .C(n785), .D(\data_in<5> ), .Y(
        n790) );
  OAI21X1 U1084 ( .A(n3160), .B(n3581), .C(n733), .Y(n1942) );
  AOI22X1 U1085 ( .A(n784), .B(\data_in<14> ), .C(n785), .D(\data_in<6> ), .Y(
        n791) );
  OAI21X1 U1086 ( .A(n3160), .B(n3580), .C(n721), .Y(n1943) );
  AOI22X1 U1087 ( .A(n784), .B(\data_in<15> ), .C(n785), .D(\data_in<7> ), .Y(
        n792) );
  AOI21X1 U1088 ( .A(n2566), .B(n2568), .C(n2452), .Y(n782) );
  OAI21X1 U1089 ( .A(n3159), .B(n3579), .C(n709), .Y(n1944) );
  AOI22X1 U1090 ( .A(n796), .B(\data_in<8> ), .C(n797), .D(\data_in<0> ), .Y(
        n795) );
  OAI21X1 U1091 ( .A(n3159), .B(n3578), .C(n697), .Y(n1945) );
  AOI22X1 U1092 ( .A(n796), .B(\data_in<9> ), .C(n797), .D(\data_in<1> ), .Y(
        n798) );
  OAI21X1 U1093 ( .A(n3159), .B(n3577), .C(n685), .Y(n1946) );
  AOI22X1 U1094 ( .A(n796), .B(\data_in<10> ), .C(n797), .D(\data_in<2> ), .Y(
        n799) );
  OAI21X1 U1095 ( .A(n3159), .B(n3576), .C(n673), .Y(n1947) );
  AOI22X1 U1096 ( .A(n796), .B(\data_in<11> ), .C(n797), .D(\data_in<3> ), .Y(
        n800) );
  OAI21X1 U1097 ( .A(n3159), .B(n3575), .C(n661), .Y(n1948) );
  AOI22X1 U1098 ( .A(n796), .B(\data_in<12> ), .C(n797), .D(\data_in<4> ), .Y(
        n801) );
  OAI21X1 U1099 ( .A(n3159), .B(n3574), .C(n649), .Y(n1949) );
  AOI22X1 U1100 ( .A(n796), .B(\data_in<13> ), .C(n797), .D(\data_in<5> ), .Y(
        n802) );
  OAI21X1 U1101 ( .A(n3159), .B(n3573), .C(n637), .Y(n1950) );
  AOI22X1 U1102 ( .A(n796), .B(\data_in<14> ), .C(n797), .D(\data_in<6> ), .Y(
        n803) );
  OAI21X1 U1103 ( .A(n3159), .B(n3572), .C(n624), .Y(n1951) );
  AOI22X1 U1104 ( .A(n796), .B(\data_in<15> ), .C(n797), .D(\data_in<7> ), .Y(
        n804) );
  AOI21X1 U1105 ( .A(n2568), .B(n2532), .C(n2452), .Y(n794) );
  OAI21X1 U1106 ( .A(n3158), .B(n3571), .C(n611), .Y(n1952) );
  AOI22X1 U1107 ( .A(n808), .B(\data_in<8> ), .C(n809), .D(\data_in<0> ), .Y(
        n807) );
  OAI21X1 U1108 ( .A(n3158), .B(n3570), .C(n609), .Y(n1953) );
  AOI22X1 U1109 ( .A(n808), .B(\data_in<9> ), .C(n809), .D(\data_in<1> ), .Y(
        n810) );
  OAI21X1 U1110 ( .A(n3158), .B(n3569), .C(n597), .Y(n1954) );
  AOI22X1 U1111 ( .A(n808), .B(\data_in<10> ), .C(n809), .D(\data_in<2> ), .Y(
        n811) );
  OAI21X1 U1112 ( .A(n3158), .B(n3568), .C(n596), .Y(n1955) );
  AOI22X1 U1113 ( .A(n808), .B(\data_in<11> ), .C(n809), .D(\data_in<3> ), .Y(
        n812) );
  OAI21X1 U1114 ( .A(n3158), .B(n3567), .C(n595), .Y(n1956) );
  AOI22X1 U1115 ( .A(n808), .B(\data_in<12> ), .C(n809), .D(\data_in<4> ), .Y(
        n813) );
  OAI21X1 U1116 ( .A(n3158), .B(n3566), .C(n594), .Y(n1957) );
  AOI22X1 U1117 ( .A(n808), .B(\data_in<13> ), .C(n809), .D(\data_in<5> ), .Y(
        n814) );
  OAI21X1 U1118 ( .A(n3158), .B(n3565), .C(n593), .Y(n1958) );
  AOI22X1 U1119 ( .A(n808), .B(\data_in<14> ), .C(n809), .D(\data_in<6> ), .Y(
        n815) );
  OAI21X1 U1120 ( .A(n3158), .B(n3564), .C(n592), .Y(n1959) );
  AOI22X1 U1121 ( .A(n808), .B(\data_in<15> ), .C(n809), .D(\data_in<7> ), .Y(
        n816) );
  AOI21X1 U1122 ( .A(n2532), .B(n2534), .C(n2452), .Y(n806) );
  OAI21X1 U1123 ( .A(n3157), .B(n3563), .C(n591), .Y(n1960) );
  AOI22X1 U1124 ( .A(n820), .B(\data_in<8> ), .C(n821), .D(\data_in<0> ), .Y(
        n819) );
  OAI21X1 U1125 ( .A(n3157), .B(n3562), .C(n590), .Y(n1961) );
  AOI22X1 U1126 ( .A(n820), .B(\data_in<9> ), .C(n821), .D(\data_in<1> ), .Y(
        n822) );
  OAI21X1 U1127 ( .A(n3157), .B(n3561), .C(n589), .Y(n1962) );
  AOI22X1 U1128 ( .A(n820), .B(\data_in<10> ), .C(n821), .D(\data_in<2> ), .Y(
        n823) );
  OAI21X1 U1129 ( .A(n3157), .B(n3560), .C(n588), .Y(n1963) );
  AOI22X1 U1130 ( .A(n820), .B(\data_in<11> ), .C(n821), .D(\data_in<3> ), .Y(
        n824) );
  OAI21X1 U1131 ( .A(n3157), .B(n3559), .C(n587), .Y(n1964) );
  AOI22X1 U1132 ( .A(n820), .B(\data_in<12> ), .C(n821), .D(\data_in<4> ), .Y(
        n825) );
  OAI21X1 U1133 ( .A(n3157), .B(n3558), .C(n586), .Y(n1965) );
  AOI22X1 U1134 ( .A(n820), .B(\data_in<13> ), .C(n821), .D(\data_in<5> ), .Y(
        n826) );
  OAI21X1 U1135 ( .A(n3157), .B(n3557), .C(n585), .Y(n1966) );
  AOI22X1 U1136 ( .A(n820), .B(\data_in<14> ), .C(n821), .D(\data_in<6> ), .Y(
        n827) );
  OAI21X1 U1137 ( .A(n3157), .B(n3556), .C(n584), .Y(n1967) );
  AOI22X1 U1138 ( .A(n820), .B(\data_in<15> ), .C(n821), .D(\data_in<7> ), .Y(
        n828) );
  AOI21X1 U1139 ( .A(n2534), .B(n2528), .C(n2452), .Y(n818) );
  OAI21X1 U1140 ( .A(n3156), .B(n3555), .C(n583), .Y(n1968) );
  AOI22X1 U1141 ( .A(n832), .B(\data_in<8> ), .C(n833), .D(\data_in<0> ), .Y(
        n831) );
  OAI21X1 U1142 ( .A(n3156), .B(n3554), .C(n582), .Y(n1969) );
  AOI22X1 U1143 ( .A(n832), .B(\data_in<9> ), .C(n833), .D(\data_in<1> ), .Y(
        n834) );
  OAI21X1 U1144 ( .A(n3156), .B(n3553), .C(n581), .Y(n1970) );
  AOI22X1 U1145 ( .A(n832), .B(\data_in<10> ), .C(n833), .D(\data_in<2> ), .Y(
        n835) );
  OAI21X1 U1146 ( .A(n3156), .B(n3552), .C(n580), .Y(n1971) );
  AOI22X1 U1147 ( .A(n832), .B(\data_in<11> ), .C(n833), .D(\data_in<3> ), .Y(
        n836) );
  OAI21X1 U1148 ( .A(n3156), .B(n3551), .C(n579), .Y(n1972) );
  AOI22X1 U1149 ( .A(n832), .B(\data_in<12> ), .C(n833), .D(\data_in<4> ), .Y(
        n837) );
  OAI21X1 U1150 ( .A(n3156), .B(n3550), .C(n578), .Y(n1973) );
  AOI22X1 U1151 ( .A(n832), .B(\data_in<13> ), .C(n833), .D(\data_in<5> ), .Y(
        n838) );
  OAI21X1 U1152 ( .A(n3156), .B(n3549), .C(n577), .Y(n1974) );
  AOI22X1 U1153 ( .A(n832), .B(\data_in<14> ), .C(n833), .D(\data_in<6> ), .Y(
        n839) );
  OAI21X1 U1154 ( .A(n3156), .B(n3548), .C(n576), .Y(n1975) );
  AOI22X1 U1155 ( .A(n832), .B(\data_in<15> ), .C(n833), .D(\data_in<7> ), .Y(
        n840) );
  AOI21X1 U1156 ( .A(n2528), .B(n2530), .C(n2452), .Y(n830) );
  OAI21X1 U1157 ( .A(n3155), .B(n3547), .C(n575), .Y(n1976) );
  AOI22X1 U1158 ( .A(n844), .B(\data_in<8> ), .C(n845), .D(\data_in<0> ), .Y(
        n843) );
  OAI21X1 U1159 ( .A(n3155), .B(n3546), .C(n574), .Y(n1977) );
  AOI22X1 U1160 ( .A(n844), .B(\data_in<9> ), .C(n845), .D(\data_in<1> ), .Y(
        n846) );
  OAI21X1 U1161 ( .A(n3155), .B(n3545), .C(n573), .Y(n1978) );
  AOI22X1 U1162 ( .A(n844), .B(\data_in<10> ), .C(n845), .D(\data_in<2> ), .Y(
        n847) );
  OAI21X1 U1163 ( .A(n3155), .B(n3544), .C(n572), .Y(n1979) );
  AOI22X1 U1164 ( .A(n844), .B(\data_in<11> ), .C(n845), .D(\data_in<3> ), .Y(
        n848) );
  OAI21X1 U1165 ( .A(n3155), .B(n3543), .C(n571), .Y(n1980) );
  AOI22X1 U1166 ( .A(n844), .B(\data_in<12> ), .C(n845), .D(\data_in<4> ), .Y(
        n849) );
  OAI21X1 U1167 ( .A(n3155), .B(n3542), .C(n570), .Y(n1981) );
  AOI22X1 U1168 ( .A(n844), .B(\data_in<13> ), .C(n845), .D(\data_in<5> ), .Y(
        n850) );
  OAI21X1 U1169 ( .A(n3155), .B(n3541), .C(n569), .Y(n1982) );
  AOI22X1 U1170 ( .A(n844), .B(\data_in<14> ), .C(n845), .D(\data_in<6> ), .Y(
        n851) );
  OAI21X1 U1171 ( .A(n3155), .B(n3540), .C(n568), .Y(n1983) );
  AOI22X1 U1172 ( .A(n844), .B(\data_in<15> ), .C(n845), .D(\data_in<7> ), .Y(
        n852) );
  AOI21X1 U1173 ( .A(n2530), .B(n2524), .C(n2452), .Y(n842) );
  OAI21X1 U1174 ( .A(n3154), .B(n3539), .C(n567), .Y(n1984) );
  AOI22X1 U1175 ( .A(n856), .B(\data_in<8> ), .C(n857), .D(\data_in<0> ), .Y(
        n855) );
  OAI21X1 U1176 ( .A(n3154), .B(n3538), .C(n566), .Y(n1985) );
  AOI22X1 U1177 ( .A(n856), .B(\data_in<9> ), .C(n857), .D(\data_in<1> ), .Y(
        n858) );
  OAI21X1 U1178 ( .A(n3154), .B(n3537), .C(n565), .Y(n1986) );
  AOI22X1 U1179 ( .A(n856), .B(\data_in<10> ), .C(n857), .D(\data_in<2> ), .Y(
        n859) );
  OAI21X1 U1180 ( .A(n3154), .B(n3536), .C(n564), .Y(n1987) );
  AOI22X1 U1181 ( .A(n856), .B(\data_in<11> ), .C(n857), .D(\data_in<3> ), .Y(
        n860) );
  OAI21X1 U1182 ( .A(n3154), .B(n3535), .C(n563), .Y(n1988) );
  AOI22X1 U1183 ( .A(n856), .B(\data_in<12> ), .C(n857), .D(\data_in<4> ), .Y(
        n861) );
  OAI21X1 U1184 ( .A(n3154), .B(n3534), .C(n562), .Y(n1989) );
  AOI22X1 U1185 ( .A(n856), .B(\data_in<13> ), .C(n857), .D(\data_in<5> ), .Y(
        n862) );
  OAI21X1 U1186 ( .A(n3154), .B(n3533), .C(n561), .Y(n1990) );
  AOI22X1 U1187 ( .A(n856), .B(\data_in<14> ), .C(n857), .D(\data_in<6> ), .Y(
        n863) );
  OAI21X1 U1188 ( .A(n3154), .B(n3532), .C(n560), .Y(n1991) );
  AOI22X1 U1189 ( .A(n856), .B(\data_in<15> ), .C(n857), .D(\data_in<7> ), .Y(
        n864) );
  AOI21X1 U1190 ( .A(n2524), .B(n2526), .C(n3177), .Y(n854) );
  OAI21X1 U1191 ( .A(n3153), .B(n3531), .C(n559), .Y(n1992) );
  AOI22X1 U1192 ( .A(n868), .B(\data_in<8> ), .C(n869), .D(\data_in<0> ), .Y(
        n867) );
  OAI21X1 U1193 ( .A(n3153), .B(n3530), .C(n558), .Y(n1993) );
  AOI22X1 U1194 ( .A(n868), .B(\data_in<9> ), .C(n869), .D(\data_in<1> ), .Y(
        n870) );
  OAI21X1 U1195 ( .A(n3153), .B(n3529), .C(n557), .Y(n1994) );
  AOI22X1 U1196 ( .A(n868), .B(\data_in<10> ), .C(n869), .D(\data_in<2> ), .Y(
        n871) );
  OAI21X1 U1197 ( .A(n3153), .B(n3528), .C(n556), .Y(n1995) );
  AOI22X1 U1198 ( .A(n868), .B(\data_in<11> ), .C(n869), .D(\data_in<3> ), .Y(
        n872) );
  OAI21X1 U1199 ( .A(n3153), .B(n3527), .C(n555), .Y(n1996) );
  AOI22X1 U1200 ( .A(n868), .B(\data_in<12> ), .C(n869), .D(\data_in<4> ), .Y(
        n873) );
  OAI21X1 U1201 ( .A(n3153), .B(n3526), .C(n554), .Y(n1997) );
  AOI22X1 U1202 ( .A(n868), .B(\data_in<13> ), .C(n869), .D(\data_in<5> ), .Y(
        n874) );
  OAI21X1 U1203 ( .A(n3153), .B(n3525), .C(n553), .Y(n1998) );
  AOI22X1 U1204 ( .A(n868), .B(\data_in<14> ), .C(n869), .D(\data_in<6> ), .Y(
        n875) );
  OAI21X1 U1205 ( .A(n3153), .B(n3524), .C(n552), .Y(n1999) );
  AOI22X1 U1206 ( .A(n868), .B(\data_in<15> ), .C(n869), .D(\data_in<7> ), .Y(
        n876) );
  AOI21X1 U1207 ( .A(n2526), .B(n2520), .C(n3177), .Y(n866) );
  OAI21X1 U1208 ( .A(n3152), .B(n3523), .C(n551), .Y(n2000) );
  AOI22X1 U1209 ( .A(n880), .B(\data_in<8> ), .C(n881), .D(\data_in<0> ), .Y(
        n879) );
  OAI21X1 U1210 ( .A(n3152), .B(n3522), .C(n550), .Y(n2001) );
  AOI22X1 U1211 ( .A(n880), .B(\data_in<9> ), .C(n881), .D(\data_in<1> ), .Y(
        n882) );
  OAI21X1 U1212 ( .A(n3152), .B(n3521), .C(n549), .Y(n2002) );
  AOI22X1 U1213 ( .A(n880), .B(\data_in<10> ), .C(n881), .D(\data_in<2> ), .Y(
        n883) );
  OAI21X1 U1214 ( .A(n3152), .B(n3520), .C(n548), .Y(n2003) );
  AOI22X1 U1215 ( .A(n880), .B(\data_in<11> ), .C(n881), .D(\data_in<3> ), .Y(
        n884) );
  OAI21X1 U1216 ( .A(n3152), .B(n3519), .C(n547), .Y(n2004) );
  AOI22X1 U1217 ( .A(n880), .B(\data_in<12> ), .C(n881), .D(\data_in<4> ), .Y(
        n885) );
  OAI21X1 U1218 ( .A(n3152), .B(n3518), .C(n546), .Y(n2005) );
  AOI22X1 U1219 ( .A(n880), .B(\data_in<13> ), .C(n881), .D(\data_in<5> ), .Y(
        n886) );
  OAI21X1 U1220 ( .A(n3152), .B(n3517), .C(n545), .Y(n2006) );
  AOI22X1 U1221 ( .A(n880), .B(\data_in<14> ), .C(n881), .D(\data_in<6> ), .Y(
        n887) );
  OAI21X1 U1222 ( .A(n3152), .B(n3516), .C(n544), .Y(n2007) );
  AOI22X1 U1223 ( .A(n880), .B(\data_in<15> ), .C(n881), .D(\data_in<7> ), .Y(
        n888) );
  AOI21X1 U1224 ( .A(n2520), .B(n2522), .C(n3177), .Y(n878) );
  OAI21X1 U1225 ( .A(n3151), .B(n3515), .C(n543), .Y(n2008) );
  AOI22X1 U1226 ( .A(n892), .B(\data_in<8> ), .C(n893), .D(\data_in<0> ), .Y(
        n891) );
  OAI21X1 U1227 ( .A(n3151), .B(n3514), .C(n542), .Y(n2009) );
  AOI22X1 U1228 ( .A(n892), .B(\data_in<9> ), .C(n893), .D(\data_in<1> ), .Y(
        n894) );
  OAI21X1 U1229 ( .A(n3151), .B(n3513), .C(n541), .Y(n2010) );
  AOI22X1 U1230 ( .A(n892), .B(\data_in<10> ), .C(n893), .D(\data_in<2> ), .Y(
        n895) );
  OAI21X1 U1231 ( .A(n3151), .B(n3512), .C(n540), .Y(n2011) );
  AOI22X1 U1232 ( .A(n892), .B(\data_in<11> ), .C(n893), .D(\data_in<3> ), .Y(
        n896) );
  OAI21X1 U1233 ( .A(n3151), .B(n3511), .C(n539), .Y(n2012) );
  AOI22X1 U1234 ( .A(n892), .B(\data_in<12> ), .C(n893), .D(\data_in<4> ), .Y(
        n897) );
  OAI21X1 U1235 ( .A(n3151), .B(n3510), .C(n538), .Y(n2013) );
  AOI22X1 U1236 ( .A(n892), .B(\data_in<13> ), .C(n893), .D(\data_in<5> ), .Y(
        n898) );
  OAI21X1 U1237 ( .A(n3151), .B(n3509), .C(n537), .Y(n2014) );
  AOI22X1 U1238 ( .A(n892), .B(\data_in<14> ), .C(n893), .D(\data_in<6> ), .Y(
        n899) );
  OAI21X1 U1239 ( .A(n3151), .B(n3508), .C(n536), .Y(n2015) );
  AOI22X1 U1240 ( .A(n892), .B(\data_in<15> ), .C(n893), .D(\data_in<7> ), .Y(
        n900) );
  AOI21X1 U1241 ( .A(n2522), .B(n2548), .C(n3177), .Y(n890) );
  OAI21X1 U1242 ( .A(n3150), .B(n3507), .C(n535), .Y(n2016) );
  AOI22X1 U1243 ( .A(n904), .B(\data_in<8> ), .C(n905), .D(\data_in<0> ), .Y(
        n903) );
  OAI21X1 U1244 ( .A(n3150), .B(n3506), .C(n534), .Y(n2017) );
  AOI22X1 U1245 ( .A(n904), .B(\data_in<9> ), .C(n905), .D(\data_in<1> ), .Y(
        n906) );
  OAI21X1 U1246 ( .A(n3150), .B(n3505), .C(n533), .Y(n2018) );
  AOI22X1 U1247 ( .A(n904), .B(\data_in<10> ), .C(n905), .D(\data_in<2> ), .Y(
        n907) );
  OAI21X1 U1248 ( .A(n3150), .B(n3504), .C(n532), .Y(n2019) );
  AOI22X1 U1249 ( .A(n904), .B(\data_in<11> ), .C(n905), .D(\data_in<3> ), .Y(
        n908) );
  OAI21X1 U1250 ( .A(n3150), .B(n3503), .C(n531), .Y(n2020) );
  AOI22X1 U1251 ( .A(n904), .B(\data_in<12> ), .C(n905), .D(\data_in<4> ), .Y(
        n909) );
  OAI21X1 U1252 ( .A(n3150), .B(n3502), .C(n530), .Y(n2021) );
  AOI22X1 U1253 ( .A(n904), .B(\data_in<13> ), .C(n905), .D(\data_in<5> ), .Y(
        n910) );
  OAI21X1 U1254 ( .A(n3150), .B(n3501), .C(n529), .Y(n2022) );
  AOI22X1 U1255 ( .A(n904), .B(\data_in<14> ), .C(n905), .D(\data_in<6> ), .Y(
        n911) );
  OAI21X1 U1256 ( .A(n3150), .B(n3500), .C(n528), .Y(n2023) );
  AOI22X1 U1257 ( .A(n904), .B(\data_in<15> ), .C(n905), .D(\data_in<7> ), .Y(
        n912) );
  AOI21X1 U1258 ( .A(n2548), .B(n2550), .C(n3177), .Y(n902) );
  OAI21X1 U1259 ( .A(n3149), .B(n3499), .C(n527), .Y(n2024) );
  AOI22X1 U1260 ( .A(n916), .B(\data_in<8> ), .C(n917), .D(\data_in<0> ), .Y(
        n915) );
  OAI21X1 U1261 ( .A(n3149), .B(n3498), .C(n526), .Y(n2025) );
  AOI22X1 U1262 ( .A(n916), .B(\data_in<9> ), .C(n917), .D(\data_in<1> ), .Y(
        n918) );
  OAI21X1 U1263 ( .A(n3149), .B(n3497), .C(n525), .Y(n2026) );
  AOI22X1 U1264 ( .A(n916), .B(\data_in<10> ), .C(n917), .D(\data_in<2> ), .Y(
        n919) );
  OAI21X1 U1265 ( .A(n3149), .B(n3496), .C(n524), .Y(n2027) );
  AOI22X1 U1266 ( .A(n916), .B(\data_in<11> ), .C(n917), .D(\data_in<3> ), .Y(
        n920) );
  OAI21X1 U1267 ( .A(n3149), .B(n3495), .C(n523), .Y(n2028) );
  AOI22X1 U1268 ( .A(n916), .B(\data_in<12> ), .C(n917), .D(\data_in<4> ), .Y(
        n921) );
  OAI21X1 U1269 ( .A(n3149), .B(n3494), .C(n522), .Y(n2029) );
  AOI22X1 U1270 ( .A(n916), .B(\data_in<13> ), .C(n917), .D(\data_in<5> ), .Y(
        n922) );
  OAI21X1 U1271 ( .A(n3149), .B(n3493), .C(n521), .Y(n2030) );
  AOI22X1 U1272 ( .A(n916), .B(\data_in<14> ), .C(n917), .D(\data_in<6> ), .Y(
        n923) );
  OAI21X1 U1273 ( .A(n3149), .B(n3492), .C(n520), .Y(n2031) );
  AOI22X1 U1274 ( .A(n916), .B(\data_in<15> ), .C(n917), .D(\data_in<7> ), .Y(
        n924) );
  AOI21X1 U1275 ( .A(n2550), .B(n2544), .C(n3177), .Y(n914) );
  OAI21X1 U1276 ( .A(n3148), .B(n3491), .C(n519), .Y(n2032) );
  AOI22X1 U1277 ( .A(n928), .B(\data_in<8> ), .C(n929), .D(\data_in<0> ), .Y(
        n927) );
  OAI21X1 U1278 ( .A(n3148), .B(n3490), .C(n518), .Y(n2033) );
  AOI22X1 U1279 ( .A(n928), .B(\data_in<9> ), .C(n929), .D(\data_in<1> ), .Y(
        n930) );
  OAI21X1 U1280 ( .A(n3148), .B(n3489), .C(n517), .Y(n2034) );
  AOI22X1 U1281 ( .A(n928), .B(\data_in<10> ), .C(n929), .D(\data_in<2> ), .Y(
        n931) );
  OAI21X1 U1282 ( .A(n3148), .B(n3488), .C(n516), .Y(n2035) );
  AOI22X1 U1283 ( .A(n928), .B(\data_in<11> ), .C(n929), .D(\data_in<3> ), .Y(
        n932) );
  OAI21X1 U1284 ( .A(n3148), .B(n3487), .C(n515), .Y(n2036) );
  AOI22X1 U1285 ( .A(n928), .B(\data_in<12> ), .C(n929), .D(\data_in<4> ), .Y(
        n933) );
  OAI21X1 U1286 ( .A(n3148), .B(n3486), .C(n514), .Y(n2037) );
  AOI22X1 U1287 ( .A(n928), .B(\data_in<13> ), .C(n929), .D(\data_in<5> ), .Y(
        n934) );
  OAI21X1 U1288 ( .A(n3148), .B(n3485), .C(n513), .Y(n2038) );
  AOI22X1 U1289 ( .A(n928), .B(\data_in<14> ), .C(n929), .D(\data_in<6> ), .Y(
        n935) );
  OAI21X1 U1290 ( .A(n3148), .B(n3484), .C(n512), .Y(n2039) );
  AOI22X1 U1291 ( .A(n928), .B(\data_in<15> ), .C(n929), .D(\data_in<7> ), .Y(
        n936) );
  AOI21X1 U1292 ( .A(n2544), .B(n2546), .C(n3177), .Y(n926) );
  OAI21X1 U1293 ( .A(n3147), .B(n3483), .C(n511), .Y(n2040) );
  AOI22X1 U1294 ( .A(n940), .B(\data_in<8> ), .C(n941), .D(\data_in<0> ), .Y(
        n939) );
  OAI21X1 U1295 ( .A(n3147), .B(n3482), .C(n510), .Y(n2041) );
  AOI22X1 U1296 ( .A(n940), .B(\data_in<9> ), .C(n941), .D(\data_in<1> ), .Y(
        n942) );
  OAI21X1 U1297 ( .A(n3147), .B(n3481), .C(n509), .Y(n2042) );
  AOI22X1 U1298 ( .A(n940), .B(\data_in<10> ), .C(n941), .D(\data_in<2> ), .Y(
        n943) );
  OAI21X1 U1299 ( .A(n3147), .B(n3480), .C(n508), .Y(n2043) );
  AOI22X1 U1300 ( .A(n940), .B(\data_in<11> ), .C(n941), .D(\data_in<3> ), .Y(
        n944) );
  OAI21X1 U1301 ( .A(n3147), .B(n3479), .C(n507), .Y(n2044) );
  AOI22X1 U1302 ( .A(n940), .B(\data_in<12> ), .C(n941), .D(\data_in<4> ), .Y(
        n945) );
  OAI21X1 U1303 ( .A(n3147), .B(n3478), .C(n506), .Y(n2045) );
  AOI22X1 U1304 ( .A(n940), .B(\data_in<13> ), .C(n941), .D(\data_in<5> ), .Y(
        n946) );
  OAI21X1 U1305 ( .A(n3147), .B(n3477), .C(n505), .Y(n2046) );
  AOI22X1 U1306 ( .A(n940), .B(\data_in<14> ), .C(n941), .D(\data_in<6> ), .Y(
        n947) );
  OAI21X1 U1307 ( .A(n3147), .B(n3476), .C(n504), .Y(n2047) );
  AOI22X1 U1308 ( .A(n940), .B(\data_in<15> ), .C(n941), .D(\data_in<7> ), .Y(
        n948) );
  AOI21X1 U1309 ( .A(n2546), .B(n2540), .C(n3177), .Y(n938) );
  OAI21X1 U1310 ( .A(n3146), .B(n3475), .C(n503), .Y(n2048) );
  AOI22X1 U1311 ( .A(n952), .B(\data_in<8> ), .C(n953), .D(\data_in<0> ), .Y(
        n951) );
  OAI21X1 U1312 ( .A(n3146), .B(n3474), .C(n502), .Y(n2049) );
  AOI22X1 U1313 ( .A(n952), .B(\data_in<9> ), .C(n953), .D(\data_in<1> ), .Y(
        n954) );
  OAI21X1 U1314 ( .A(n3146), .B(n3473), .C(n501), .Y(n2050) );
  AOI22X1 U1315 ( .A(n952), .B(\data_in<10> ), .C(n953), .D(\data_in<2> ), .Y(
        n955) );
  OAI21X1 U1316 ( .A(n3146), .B(n3472), .C(n500), .Y(n2051) );
  AOI22X1 U1317 ( .A(n952), .B(\data_in<11> ), .C(n953), .D(\data_in<3> ), .Y(
        n956) );
  OAI21X1 U1318 ( .A(n3146), .B(n3471), .C(n499), .Y(n2052) );
  AOI22X1 U1319 ( .A(n952), .B(\data_in<12> ), .C(n953), .D(\data_in<4> ), .Y(
        n957) );
  OAI21X1 U1320 ( .A(n3146), .B(n3470), .C(n498), .Y(n2053) );
  AOI22X1 U1321 ( .A(n952), .B(\data_in<13> ), .C(n953), .D(\data_in<5> ), .Y(
        n958) );
  OAI21X1 U1322 ( .A(n3146), .B(n3469), .C(n497), .Y(n2054) );
  AOI22X1 U1323 ( .A(n952), .B(\data_in<14> ), .C(n953), .D(\data_in<6> ), .Y(
        n959) );
  OAI21X1 U1324 ( .A(n3146), .B(n3468), .C(n496), .Y(n2055) );
  AOI22X1 U1325 ( .A(n952), .B(\data_in<15> ), .C(n953), .D(\data_in<7> ), .Y(
        n960) );
  AOI21X1 U1326 ( .A(n2540), .B(n2542), .C(n3177), .Y(n950) );
  OAI21X1 U1327 ( .A(n3145), .B(n3467), .C(n495), .Y(n2056) );
  AOI22X1 U1328 ( .A(n964), .B(\data_in<8> ), .C(n965), .D(\data_in<0> ), .Y(
        n963) );
  OAI21X1 U1329 ( .A(n3145), .B(n3466), .C(n494), .Y(n2057) );
  AOI22X1 U1330 ( .A(n964), .B(\data_in<9> ), .C(n965), .D(\data_in<1> ), .Y(
        n966) );
  OAI21X1 U1331 ( .A(n3145), .B(n3465), .C(n493), .Y(n2058) );
  AOI22X1 U1332 ( .A(n964), .B(\data_in<10> ), .C(n965), .D(\data_in<2> ), .Y(
        n967) );
  OAI21X1 U1333 ( .A(n3145), .B(n3464), .C(n492), .Y(n2059) );
  AOI22X1 U1334 ( .A(n964), .B(\data_in<11> ), .C(n965), .D(\data_in<3> ), .Y(
        n968) );
  OAI21X1 U1335 ( .A(n3145), .B(n3463), .C(n491), .Y(n2060) );
  AOI22X1 U1336 ( .A(n964), .B(\data_in<12> ), .C(n965), .D(\data_in<4> ), .Y(
        n969) );
  OAI21X1 U1337 ( .A(n3145), .B(n3462), .C(n490), .Y(n2061) );
  AOI22X1 U1338 ( .A(n964), .B(\data_in<13> ), .C(n965), .D(\data_in<5> ), .Y(
        n970) );
  OAI21X1 U1339 ( .A(n3145), .B(n3461), .C(n489), .Y(n2062) );
  AOI22X1 U1340 ( .A(n964), .B(\data_in<14> ), .C(n965), .D(\data_in<6> ), .Y(
        n971) );
  OAI21X1 U1341 ( .A(n3145), .B(n3460), .C(n488), .Y(n2063) );
  AOI22X1 U1342 ( .A(n964), .B(\data_in<15> ), .C(n965), .D(\data_in<7> ), .Y(
        n972) );
  AOI21X1 U1343 ( .A(n2542), .B(n2535), .C(n3177), .Y(n962) );
  OAI21X1 U1344 ( .A(n3144), .B(n3459), .C(n487), .Y(n2064) );
  AOI22X1 U1345 ( .A(n976), .B(\data_in<8> ), .C(n977), .D(\data_in<0> ), .Y(
        n975) );
  OAI21X1 U1346 ( .A(n3144), .B(n3458), .C(n486), .Y(n2065) );
  AOI22X1 U1347 ( .A(n976), .B(\data_in<9> ), .C(n977), .D(\data_in<1> ), .Y(
        n978) );
  OAI21X1 U1348 ( .A(n3144), .B(n3457), .C(n485), .Y(n2066) );
  AOI22X1 U1349 ( .A(n976), .B(\data_in<10> ), .C(n977), .D(\data_in<2> ), .Y(
        n979) );
  OAI21X1 U1350 ( .A(n3144), .B(n3456), .C(n484), .Y(n2067) );
  AOI22X1 U1351 ( .A(n976), .B(\data_in<11> ), .C(n977), .D(\data_in<3> ), .Y(
        n980) );
  OAI21X1 U1352 ( .A(n3144), .B(n3455), .C(n483), .Y(n2068) );
  AOI22X1 U1353 ( .A(n976), .B(\data_in<12> ), .C(n977), .D(\data_in<4> ), .Y(
        n981) );
  OAI21X1 U1354 ( .A(n3144), .B(n3454), .C(n482), .Y(n2069) );
  AOI22X1 U1355 ( .A(n976), .B(\data_in<13> ), .C(n977), .D(\data_in<5> ), .Y(
        n982) );
  OAI21X1 U1356 ( .A(n3144), .B(n3453), .C(n481), .Y(n2070) );
  AOI22X1 U1357 ( .A(n976), .B(\data_in<14> ), .C(n977), .D(\data_in<6> ), .Y(
        n983) );
  OAI21X1 U1358 ( .A(n3144), .B(n3452), .C(n480), .Y(n2071) );
  AOI22X1 U1359 ( .A(n976), .B(\data_in<15> ), .C(n977), .D(\data_in<7> ), .Y(
        n984) );
  AOI21X1 U1360 ( .A(n2535), .B(n2538), .C(n3177), .Y(n974) );
  OAI21X1 U1361 ( .A(n3143), .B(n3451), .C(n479), .Y(n2072) );
  AOI22X1 U1362 ( .A(n988), .B(\data_in<8> ), .C(n989), .D(\data_in<0> ), .Y(
        n987) );
  OAI21X1 U1363 ( .A(n3143), .B(n3450), .C(n478), .Y(n2073) );
  AOI22X1 U1364 ( .A(n988), .B(\data_in<9> ), .C(n989), .D(\data_in<1> ), .Y(
        n990) );
  OAI21X1 U1365 ( .A(n3143), .B(n3449), .C(n477), .Y(n2074) );
  AOI22X1 U1366 ( .A(n988), .B(\data_in<10> ), .C(n989), .D(\data_in<2> ), .Y(
        n991) );
  OAI21X1 U1367 ( .A(n3143), .B(n3448), .C(n476), .Y(n2075) );
  AOI22X1 U1368 ( .A(n988), .B(\data_in<11> ), .C(n989), .D(\data_in<3> ), .Y(
        n992) );
  OAI21X1 U1369 ( .A(n3143), .B(n3447), .C(n475), .Y(n2076) );
  AOI22X1 U1370 ( .A(n988), .B(\data_in<12> ), .C(n989), .D(\data_in<4> ), .Y(
        n993) );
  OAI21X1 U1371 ( .A(n3143), .B(n3446), .C(n474), .Y(n2077) );
  AOI22X1 U1372 ( .A(n988), .B(\data_in<13> ), .C(n989), .D(\data_in<5> ), .Y(
        n994) );
  OAI21X1 U1373 ( .A(n3143), .B(n3445), .C(n473), .Y(n2078) );
  AOI22X1 U1374 ( .A(n988), .B(\data_in<14> ), .C(n989), .D(\data_in<6> ), .Y(
        n995) );
  OAI21X1 U1375 ( .A(n3143), .B(n3444), .C(n472), .Y(n2079) );
  AOI22X1 U1376 ( .A(n988), .B(\data_in<15> ), .C(n989), .D(\data_in<7> ), .Y(
        n996) );
  AOI21X1 U1377 ( .A(n2538), .B(n2474), .C(n3177), .Y(n986) );
  OAI21X1 U1378 ( .A(n3142), .B(n3443), .C(n471), .Y(n2080) );
  AOI22X1 U1379 ( .A(n1000), .B(\data_in<8> ), .C(n1001), .D(\data_in<0> ), 
        .Y(n999) );
  OAI21X1 U1380 ( .A(n3142), .B(n3442), .C(n470), .Y(n2081) );
  AOI22X1 U1381 ( .A(n1000), .B(\data_in<9> ), .C(n1001), .D(\data_in<1> ), 
        .Y(n1002) );
  OAI21X1 U1382 ( .A(n3142), .B(n3441), .C(n469), .Y(n2082) );
  AOI22X1 U1383 ( .A(n1000), .B(\data_in<10> ), .C(n1001), .D(\data_in<2> ), 
        .Y(n1003) );
  OAI21X1 U1384 ( .A(n3142), .B(n3440), .C(n468), .Y(n2083) );
  AOI22X1 U1385 ( .A(n1000), .B(\data_in<11> ), .C(n1001), .D(\data_in<3> ), 
        .Y(n1004) );
  OAI21X1 U1386 ( .A(n3142), .B(n3439), .C(n467), .Y(n2084) );
  AOI22X1 U1387 ( .A(n1000), .B(\data_in<12> ), .C(n1001), .D(\data_in<4> ), 
        .Y(n1005) );
  OAI21X1 U1388 ( .A(n3142), .B(n3438), .C(n466), .Y(n2085) );
  AOI22X1 U1389 ( .A(n1000), .B(\data_in<13> ), .C(n1001), .D(\data_in<5> ), 
        .Y(n1006) );
  OAI21X1 U1390 ( .A(n3142), .B(n3437), .C(n465), .Y(n2086) );
  AOI22X1 U1391 ( .A(n1000), .B(\data_in<14> ), .C(n1001), .D(\data_in<6> ), 
        .Y(n1007) );
  OAI21X1 U1392 ( .A(n3142), .B(n3436), .C(n464), .Y(n2087) );
  AOI22X1 U1393 ( .A(n1000), .B(\data_in<15> ), .C(n1001), .D(\data_in<7> ), 
        .Y(n1008) );
  AOI21X1 U1394 ( .A(n2474), .B(n2476), .C(n3177), .Y(n998) );
  OAI21X1 U1395 ( .A(n3141), .B(n3435), .C(n463), .Y(n2088) );
  AOI22X1 U1396 ( .A(n1012), .B(\data_in<8> ), .C(n1013), .D(\data_in<0> ), 
        .Y(n1011) );
  OAI21X1 U1397 ( .A(n3141), .B(n3434), .C(n462), .Y(n2089) );
  AOI22X1 U1398 ( .A(n1012), .B(\data_in<9> ), .C(n1013), .D(\data_in<1> ), 
        .Y(n1014) );
  OAI21X1 U1399 ( .A(n3141), .B(n3433), .C(n461), .Y(n2090) );
  AOI22X1 U1400 ( .A(n1012), .B(\data_in<10> ), .C(n1013), .D(\data_in<2> ), 
        .Y(n1015) );
  OAI21X1 U1401 ( .A(n3141), .B(n3432), .C(n460), .Y(n2091) );
  AOI22X1 U1402 ( .A(n1012), .B(\data_in<11> ), .C(n1013), .D(\data_in<3> ), 
        .Y(n1016) );
  OAI21X1 U1403 ( .A(n3141), .B(n3431), .C(n459), .Y(n2092) );
  AOI22X1 U1404 ( .A(n1012), .B(\data_in<12> ), .C(n1013), .D(\data_in<4> ), 
        .Y(n1017) );
  OAI21X1 U1405 ( .A(n3141), .B(n3430), .C(n458), .Y(n2093) );
  AOI22X1 U1406 ( .A(n1012), .B(\data_in<13> ), .C(n1013), .D(\data_in<5> ), 
        .Y(n1018) );
  OAI21X1 U1407 ( .A(n3141), .B(n3429), .C(n457), .Y(n2094) );
  AOI22X1 U1408 ( .A(n1012), .B(\data_in<14> ), .C(n1013), .D(\data_in<6> ), 
        .Y(n1019) );
  OAI21X1 U1409 ( .A(n3141), .B(n3428), .C(n456), .Y(n2095) );
  AOI22X1 U1410 ( .A(n1012), .B(\data_in<15> ), .C(n1013), .D(\data_in<7> ), 
        .Y(n1020) );
  AOI21X1 U1411 ( .A(n2476), .B(n2470), .C(n3177), .Y(n1010) );
  OAI21X1 U1412 ( .A(n3140), .B(n3427), .C(n455), .Y(n2096) );
  AOI22X1 U1413 ( .A(n1024), .B(\data_in<8> ), .C(n1025), .D(\data_in<0> ), 
        .Y(n1023) );
  OAI21X1 U1414 ( .A(n3140), .B(n3426), .C(n454), .Y(n2097) );
  AOI22X1 U1415 ( .A(n1024), .B(\data_in<9> ), .C(n1025), .D(\data_in<1> ), 
        .Y(n1026) );
  OAI21X1 U1416 ( .A(n3140), .B(n3425), .C(n453), .Y(n2098) );
  AOI22X1 U1417 ( .A(n1024), .B(\data_in<10> ), .C(n1025), .D(\data_in<2> ), 
        .Y(n1027) );
  OAI21X1 U1418 ( .A(n3140), .B(n3424), .C(n452), .Y(n2099) );
  AOI22X1 U1419 ( .A(n1024), .B(\data_in<11> ), .C(n1025), .D(\data_in<3> ), 
        .Y(n1028) );
  OAI21X1 U1420 ( .A(n3140), .B(n3423), .C(n451), .Y(n2100) );
  AOI22X1 U1421 ( .A(n1024), .B(\data_in<12> ), .C(n1025), .D(\data_in<4> ), 
        .Y(n1029) );
  OAI21X1 U1422 ( .A(n3140), .B(n3422), .C(n450), .Y(n2101) );
  AOI22X1 U1423 ( .A(n1024), .B(\data_in<13> ), .C(n1025), .D(\data_in<5> ), 
        .Y(n1030) );
  OAI21X1 U1424 ( .A(n3140), .B(n3421), .C(n449), .Y(n2102) );
  AOI22X1 U1425 ( .A(n1024), .B(\data_in<14> ), .C(n1025), .D(\data_in<6> ), 
        .Y(n1031) );
  OAI21X1 U1426 ( .A(n3140), .B(n3420), .C(n448), .Y(n2103) );
  AOI22X1 U1427 ( .A(n1024), .B(\data_in<15> ), .C(n1025), .D(\data_in<7> ), 
        .Y(n1032) );
  AOI21X1 U1428 ( .A(n2470), .B(n2472), .C(n3176), .Y(n1022) );
  OAI21X1 U1429 ( .A(n3139), .B(n3419), .C(n447), .Y(n2104) );
  AOI22X1 U1430 ( .A(n1036), .B(\data_in<8> ), .C(n1037), .D(\data_in<0> ), 
        .Y(n1035) );
  OAI21X1 U1431 ( .A(n3139), .B(n3418), .C(n446), .Y(n2105) );
  AOI22X1 U1432 ( .A(n1036), .B(\data_in<9> ), .C(n1037), .D(\data_in<1> ), 
        .Y(n1038) );
  OAI21X1 U1433 ( .A(n3139), .B(n3417), .C(n445), .Y(n2106) );
  AOI22X1 U1434 ( .A(n1036), .B(\data_in<10> ), .C(n1037), .D(\data_in<2> ), 
        .Y(n1039) );
  OAI21X1 U1435 ( .A(n3139), .B(n3416), .C(n444), .Y(n2107) );
  AOI22X1 U1436 ( .A(n1036), .B(\data_in<11> ), .C(n1037), .D(\data_in<3> ), 
        .Y(n1040) );
  OAI21X1 U1437 ( .A(n3139), .B(n3415), .C(n443), .Y(n2108) );
  AOI22X1 U1438 ( .A(n1036), .B(\data_in<12> ), .C(n1037), .D(\data_in<4> ), 
        .Y(n1041) );
  OAI21X1 U1439 ( .A(n3139), .B(n3414), .C(n442), .Y(n2109) );
  AOI22X1 U1440 ( .A(n1036), .B(\data_in<13> ), .C(n1037), .D(\data_in<5> ), 
        .Y(n1042) );
  OAI21X1 U1441 ( .A(n3139), .B(n3413), .C(n441), .Y(n2110) );
  AOI22X1 U1442 ( .A(n1036), .B(\data_in<14> ), .C(n1037), .D(\data_in<6> ), 
        .Y(n1043) );
  OAI21X1 U1443 ( .A(n3139), .B(n3412), .C(n440), .Y(n2111) );
  AOI22X1 U1444 ( .A(n1036), .B(\data_in<15> ), .C(n1037), .D(\data_in<7> ), 
        .Y(n1044) );
  AOI21X1 U1445 ( .A(n2472), .B(n2466), .C(n3176), .Y(n1034) );
  OAI21X1 U1446 ( .A(n3138), .B(n3411), .C(n439), .Y(n2112) );
  AOI22X1 U1447 ( .A(n1048), .B(\data_in<8> ), .C(n1049), .D(\data_in<0> ), 
        .Y(n1047) );
  OAI21X1 U1448 ( .A(n3138), .B(n3410), .C(n438), .Y(n2113) );
  AOI22X1 U1449 ( .A(n1048), .B(\data_in<9> ), .C(n1049), .D(\data_in<1> ), 
        .Y(n1050) );
  OAI21X1 U1450 ( .A(n3138), .B(n3409), .C(n437), .Y(n2114) );
  AOI22X1 U1451 ( .A(n1048), .B(\data_in<10> ), .C(n1049), .D(\data_in<2> ), 
        .Y(n1051) );
  OAI21X1 U1452 ( .A(n3138), .B(n3408), .C(n436), .Y(n2115) );
  AOI22X1 U1453 ( .A(n1048), .B(\data_in<11> ), .C(n1049), .D(\data_in<3> ), 
        .Y(n1052) );
  OAI21X1 U1454 ( .A(n3138), .B(n3407), .C(n435), .Y(n2116) );
  AOI22X1 U1455 ( .A(n1048), .B(\data_in<12> ), .C(n1049), .D(\data_in<4> ), 
        .Y(n1053) );
  OAI21X1 U1456 ( .A(n3138), .B(n3406), .C(n434), .Y(n2117) );
  AOI22X1 U1457 ( .A(n1048), .B(\data_in<13> ), .C(n1049), .D(\data_in<5> ), 
        .Y(n1054) );
  OAI21X1 U1458 ( .A(n3138), .B(n3405), .C(n433), .Y(n2118) );
  AOI22X1 U1459 ( .A(n1048), .B(\data_in<14> ), .C(n1049), .D(\data_in<6> ), 
        .Y(n1055) );
  OAI21X1 U1460 ( .A(n3138), .B(n3404), .C(n432), .Y(n2119) );
  AOI22X1 U1461 ( .A(n1048), .B(\data_in<15> ), .C(n1049), .D(\data_in<7> ), 
        .Y(n1056) );
  AOI21X1 U1462 ( .A(n2466), .B(n2468), .C(n3176), .Y(n1046) );
  OAI21X1 U1463 ( .A(n3137), .B(n3403), .C(n431), .Y(n2120) );
  AOI22X1 U1464 ( .A(n1060), .B(\data_in<8> ), .C(n1061), .D(\data_in<0> ), 
        .Y(n1059) );
  OAI21X1 U1465 ( .A(n3137), .B(n3402), .C(n430), .Y(n2121) );
  AOI22X1 U1466 ( .A(n1060), .B(\data_in<9> ), .C(n1061), .D(\data_in<1> ), 
        .Y(n1062) );
  OAI21X1 U1467 ( .A(n3137), .B(n3401), .C(n429), .Y(n2122) );
  AOI22X1 U1468 ( .A(n1060), .B(\data_in<10> ), .C(n1061), .D(\data_in<2> ), 
        .Y(n1063) );
  OAI21X1 U1469 ( .A(n3137), .B(n3400), .C(n428), .Y(n2123) );
  AOI22X1 U1470 ( .A(n1060), .B(\data_in<11> ), .C(n1061), .D(\data_in<3> ), 
        .Y(n1064) );
  OAI21X1 U1471 ( .A(n3137), .B(n3399), .C(n427), .Y(n2124) );
  AOI22X1 U1472 ( .A(n1060), .B(\data_in<12> ), .C(n1061), .D(\data_in<4> ), 
        .Y(n1065) );
  OAI21X1 U1473 ( .A(n3137), .B(n3398), .C(n426), .Y(n2125) );
  AOI22X1 U1474 ( .A(n1060), .B(\data_in<13> ), .C(n1061), .D(\data_in<5> ), 
        .Y(n1066) );
  OAI21X1 U1475 ( .A(n3137), .B(n3397), .C(n425), .Y(n2126) );
  AOI22X1 U1476 ( .A(n1060), .B(\data_in<14> ), .C(n1061), .D(\data_in<6> ), 
        .Y(n1067) );
  OAI21X1 U1477 ( .A(n3137), .B(n3396), .C(n424), .Y(n2127) );
  AOI22X1 U1478 ( .A(n1060), .B(\data_in<15> ), .C(n1061), .D(\data_in<7> ), 
        .Y(n1068) );
  AOI21X1 U1479 ( .A(n2468), .B(n2462), .C(n3176), .Y(n1058) );
  OAI21X1 U1480 ( .A(n3136), .B(n3395), .C(n423), .Y(n2128) );
  AOI22X1 U1481 ( .A(n1072), .B(\data_in<8> ), .C(n1073), .D(\data_in<0> ), 
        .Y(n1071) );
  OAI21X1 U1482 ( .A(n3136), .B(n3394), .C(n422), .Y(n2129) );
  AOI22X1 U1483 ( .A(n1072), .B(\data_in<9> ), .C(n1073), .D(\data_in<1> ), 
        .Y(n1074) );
  OAI21X1 U1484 ( .A(n3136), .B(n3393), .C(n421), .Y(n2130) );
  AOI22X1 U1485 ( .A(n1072), .B(\data_in<10> ), .C(n1073), .D(\data_in<2> ), 
        .Y(n1075) );
  OAI21X1 U1486 ( .A(n3136), .B(n3392), .C(n420), .Y(n2131) );
  AOI22X1 U1487 ( .A(n1072), .B(\data_in<11> ), .C(n1073), .D(\data_in<3> ), 
        .Y(n1076) );
  OAI21X1 U1488 ( .A(n3136), .B(n3391), .C(n419), .Y(n2132) );
  AOI22X1 U1489 ( .A(n1072), .B(\data_in<12> ), .C(n1073), .D(\data_in<4> ), 
        .Y(n1077) );
  OAI21X1 U1490 ( .A(n3136), .B(n3390), .C(n418), .Y(n2133) );
  AOI22X1 U1491 ( .A(n1072), .B(\data_in<13> ), .C(n1073), .D(\data_in<5> ), 
        .Y(n1078) );
  OAI21X1 U1492 ( .A(n3136), .B(n3389), .C(n417), .Y(n2134) );
  AOI22X1 U1493 ( .A(n1072), .B(\data_in<14> ), .C(n1073), .D(\data_in<6> ), 
        .Y(n1079) );
  OAI21X1 U1494 ( .A(n3136), .B(n3388), .C(n416), .Y(n2135) );
  AOI22X1 U1495 ( .A(n1072), .B(\data_in<15> ), .C(n1073), .D(\data_in<7> ), 
        .Y(n1080) );
  AOI21X1 U1496 ( .A(n2462), .B(n2464), .C(n3176), .Y(n1070) );
  OAI21X1 U1497 ( .A(n3135), .B(n3387), .C(n415), .Y(n2136) );
  AOI22X1 U1498 ( .A(n1084), .B(\data_in<8> ), .C(n1085), .D(\data_in<0> ), 
        .Y(n1083) );
  OAI21X1 U1499 ( .A(n3135), .B(n3386), .C(n414), .Y(n2137) );
  AOI22X1 U1500 ( .A(n1084), .B(\data_in<9> ), .C(n1085), .D(\data_in<1> ), 
        .Y(n1086) );
  OAI21X1 U1501 ( .A(n3135), .B(n3385), .C(n413), .Y(n2138) );
  AOI22X1 U1502 ( .A(n1084), .B(\data_in<10> ), .C(n1085), .D(\data_in<2> ), 
        .Y(n1087) );
  OAI21X1 U1503 ( .A(n3135), .B(n3384), .C(n412), .Y(n2139) );
  AOI22X1 U1504 ( .A(n1084), .B(\data_in<11> ), .C(n1085), .D(\data_in<3> ), 
        .Y(n1088) );
  OAI21X1 U1505 ( .A(n3135), .B(n3383), .C(n411), .Y(n2140) );
  AOI22X1 U1506 ( .A(n1084), .B(\data_in<12> ), .C(n1085), .D(\data_in<4> ), 
        .Y(n1089) );
  OAI21X1 U1507 ( .A(n3135), .B(n3382), .C(n410), .Y(n2141) );
  AOI22X1 U1508 ( .A(n1084), .B(\data_in<13> ), .C(n1085), .D(\data_in<5> ), 
        .Y(n1090) );
  OAI21X1 U1509 ( .A(n3135), .B(n3381), .C(n409), .Y(n2142) );
  AOI22X1 U1510 ( .A(n1084), .B(\data_in<14> ), .C(n1085), .D(\data_in<6> ), 
        .Y(n1091) );
  OAI21X1 U1511 ( .A(n3135), .B(n3380), .C(n408), .Y(n2143) );
  AOI22X1 U1512 ( .A(n1084), .B(\data_in<15> ), .C(n1085), .D(\data_in<7> ), 
        .Y(n1092) );
  AOI21X1 U1513 ( .A(n2464), .B(n2490), .C(n3176), .Y(n1082) );
  OAI21X1 U1514 ( .A(n3134), .B(n3379), .C(n407), .Y(n2144) );
  AOI22X1 U1515 ( .A(n1096), .B(\data_in<8> ), .C(n1097), .D(\data_in<0> ), 
        .Y(n1095) );
  OAI21X1 U1516 ( .A(n3134), .B(n3378), .C(n406), .Y(n2145) );
  AOI22X1 U1517 ( .A(n1096), .B(\data_in<9> ), .C(n1097), .D(\data_in<1> ), 
        .Y(n1098) );
  OAI21X1 U1518 ( .A(n3134), .B(n3377), .C(n405), .Y(n2146) );
  AOI22X1 U1519 ( .A(n1096), .B(\data_in<10> ), .C(n1097), .D(\data_in<2> ), 
        .Y(n1099) );
  OAI21X1 U1520 ( .A(n3134), .B(n3376), .C(n404), .Y(n2147) );
  AOI22X1 U1521 ( .A(n1096), .B(\data_in<11> ), .C(n1097), .D(\data_in<3> ), 
        .Y(n1100) );
  OAI21X1 U1522 ( .A(n3134), .B(n3375), .C(n403), .Y(n2148) );
  AOI22X1 U1523 ( .A(n1096), .B(\data_in<12> ), .C(n1097), .D(\data_in<4> ), 
        .Y(n1101) );
  OAI21X1 U1524 ( .A(n3134), .B(n3374), .C(n402), .Y(n2149) );
  AOI22X1 U1525 ( .A(n1096), .B(\data_in<13> ), .C(n1097), .D(\data_in<5> ), 
        .Y(n1102) );
  OAI21X1 U1526 ( .A(n3134), .B(n3373), .C(n401), .Y(n2150) );
  AOI22X1 U1527 ( .A(n1096), .B(\data_in<14> ), .C(n1097), .D(\data_in<6> ), 
        .Y(n1103) );
  OAI21X1 U1528 ( .A(n3134), .B(n3372), .C(n400), .Y(n2151) );
  AOI22X1 U1529 ( .A(n1096), .B(\data_in<15> ), .C(n1097), .D(\data_in<7> ), 
        .Y(n1104) );
  AOI21X1 U1530 ( .A(n2490), .B(n2492), .C(n3176), .Y(n1094) );
  OAI21X1 U1531 ( .A(n3133), .B(n3371), .C(n399), .Y(n2152) );
  AOI22X1 U1532 ( .A(n1108), .B(\data_in<8> ), .C(n1109), .D(\data_in<0> ), 
        .Y(n1107) );
  OAI21X1 U1533 ( .A(n3133), .B(n3370), .C(n398), .Y(n2153) );
  AOI22X1 U1534 ( .A(n1108), .B(\data_in<9> ), .C(n1109), .D(\data_in<1> ), 
        .Y(n1110) );
  OAI21X1 U1535 ( .A(n3133), .B(n3369), .C(n397), .Y(n2154) );
  AOI22X1 U1536 ( .A(n1108), .B(\data_in<10> ), .C(n1109), .D(\data_in<2> ), 
        .Y(n1111) );
  OAI21X1 U1537 ( .A(n3133), .B(n3368), .C(n396), .Y(n2155) );
  AOI22X1 U1538 ( .A(n1108), .B(\data_in<11> ), .C(n1109), .D(\data_in<3> ), 
        .Y(n1112) );
  OAI21X1 U1539 ( .A(n3133), .B(n3367), .C(n395), .Y(n2156) );
  AOI22X1 U1540 ( .A(n1108), .B(\data_in<12> ), .C(n1109), .D(\data_in<4> ), 
        .Y(n1113) );
  OAI21X1 U1541 ( .A(n3133), .B(n3366), .C(n394), .Y(n2157) );
  AOI22X1 U1542 ( .A(n1108), .B(\data_in<13> ), .C(n1109), .D(\data_in<5> ), 
        .Y(n1114) );
  OAI21X1 U1543 ( .A(n3133), .B(n3365), .C(n393), .Y(n2158) );
  AOI22X1 U1544 ( .A(n1108), .B(\data_in<14> ), .C(n1109), .D(\data_in<6> ), 
        .Y(n1115) );
  OAI21X1 U1545 ( .A(n3133), .B(n3364), .C(n392), .Y(n2159) );
  AOI22X1 U1546 ( .A(n1108), .B(\data_in<15> ), .C(n1109), .D(\data_in<7> ), 
        .Y(n1116) );
  AOI21X1 U1547 ( .A(n2492), .B(n2486), .C(n3176), .Y(n1106) );
  OAI21X1 U1548 ( .A(n3132), .B(n3363), .C(n391), .Y(n2160) );
  AOI22X1 U1549 ( .A(n1120), .B(\data_in<8> ), .C(n1121), .D(\data_in<0> ), 
        .Y(n1119) );
  OAI21X1 U1550 ( .A(n3132), .B(n3362), .C(n390), .Y(n2161) );
  AOI22X1 U1551 ( .A(n1120), .B(\data_in<9> ), .C(n1121), .D(\data_in<1> ), 
        .Y(n1122) );
  OAI21X1 U1552 ( .A(n3132), .B(n3361), .C(n389), .Y(n2162) );
  AOI22X1 U1553 ( .A(n1120), .B(\data_in<10> ), .C(n1121), .D(\data_in<2> ), 
        .Y(n1123) );
  OAI21X1 U1554 ( .A(n3132), .B(n3360), .C(n388), .Y(n2163) );
  AOI22X1 U1555 ( .A(n1120), .B(\data_in<11> ), .C(n1121), .D(\data_in<3> ), 
        .Y(n1124) );
  OAI21X1 U1556 ( .A(n3132), .B(n3359), .C(n387), .Y(n2164) );
  AOI22X1 U1557 ( .A(n1120), .B(\data_in<12> ), .C(n1121), .D(\data_in<4> ), 
        .Y(n1125) );
  OAI21X1 U1558 ( .A(n3132), .B(n3358), .C(n386), .Y(n2165) );
  AOI22X1 U1559 ( .A(n1120), .B(\data_in<13> ), .C(n1121), .D(\data_in<5> ), 
        .Y(n1126) );
  OAI21X1 U1560 ( .A(n3132), .B(n3357), .C(n385), .Y(n2166) );
  AOI22X1 U1561 ( .A(n1120), .B(\data_in<14> ), .C(n1121), .D(\data_in<6> ), 
        .Y(n1127) );
  OAI21X1 U1562 ( .A(n3132), .B(n3356), .C(n384), .Y(n2167) );
  AOI22X1 U1563 ( .A(n1120), .B(\data_in<15> ), .C(n1121), .D(\data_in<7> ), 
        .Y(n1128) );
  AOI21X1 U1564 ( .A(n2486), .B(n2488), .C(n3176), .Y(n1118) );
  OAI21X1 U1565 ( .A(n3131), .B(n3355), .C(n383), .Y(n2168) );
  AOI22X1 U1566 ( .A(n1132), .B(\data_in<8> ), .C(n1133), .D(\data_in<0> ), 
        .Y(n1131) );
  OAI21X1 U1567 ( .A(n3131), .B(n3354), .C(n382), .Y(n2169) );
  AOI22X1 U1568 ( .A(n1132), .B(\data_in<9> ), .C(n1133), .D(\data_in<1> ), 
        .Y(n1134) );
  OAI21X1 U1569 ( .A(n3131), .B(n3353), .C(n381), .Y(n2170) );
  AOI22X1 U1570 ( .A(n1132), .B(\data_in<10> ), .C(n1133), .D(\data_in<2> ), 
        .Y(n1135) );
  OAI21X1 U1571 ( .A(n3131), .B(n3352), .C(n380), .Y(n2171) );
  AOI22X1 U1572 ( .A(n1132), .B(\data_in<11> ), .C(n1133), .D(\data_in<3> ), 
        .Y(n1136) );
  OAI21X1 U1573 ( .A(n3131), .B(n3351), .C(n379), .Y(n2172) );
  AOI22X1 U1574 ( .A(n1132), .B(\data_in<12> ), .C(n1133), .D(\data_in<4> ), 
        .Y(n1137) );
  OAI21X1 U1575 ( .A(n3131), .B(n3350), .C(n378), .Y(n2173) );
  AOI22X1 U1576 ( .A(n1132), .B(\data_in<13> ), .C(n1133), .D(\data_in<5> ), 
        .Y(n1138) );
  OAI21X1 U1577 ( .A(n3131), .B(n3349), .C(n377), .Y(n2174) );
  AOI22X1 U1578 ( .A(n1132), .B(\data_in<14> ), .C(n1133), .D(\data_in<6> ), 
        .Y(n1139) );
  OAI21X1 U1579 ( .A(n3131), .B(n3348), .C(n376), .Y(n2175) );
  AOI22X1 U1580 ( .A(n1132), .B(\data_in<15> ), .C(n1133), .D(\data_in<7> ), 
        .Y(n1140) );
  AOI21X1 U1581 ( .A(n2488), .B(n2482), .C(n3176), .Y(n1130) );
  OAI21X1 U1582 ( .A(n3130), .B(n3347), .C(n375), .Y(n2176) );
  AOI22X1 U1583 ( .A(n1144), .B(\data_in<8> ), .C(n1145), .D(\data_in<0> ), 
        .Y(n1143) );
  OAI21X1 U1584 ( .A(n3130), .B(n3346), .C(n374), .Y(n2177) );
  AOI22X1 U1585 ( .A(n1144), .B(\data_in<9> ), .C(n1145), .D(\data_in<1> ), 
        .Y(n1146) );
  OAI21X1 U1586 ( .A(n3130), .B(n3345), .C(n373), .Y(n2178) );
  AOI22X1 U1587 ( .A(n1144), .B(\data_in<10> ), .C(n1145), .D(\data_in<2> ), 
        .Y(n1147) );
  OAI21X1 U1588 ( .A(n3130), .B(n3344), .C(n372), .Y(n2179) );
  AOI22X1 U1589 ( .A(n1144), .B(\data_in<11> ), .C(n1145), .D(\data_in<3> ), 
        .Y(n1148) );
  OAI21X1 U1590 ( .A(n3130), .B(n3343), .C(n371), .Y(n2180) );
  AOI22X1 U1591 ( .A(n1144), .B(\data_in<12> ), .C(n1145), .D(\data_in<4> ), 
        .Y(n1149) );
  OAI21X1 U1592 ( .A(n3130), .B(n3342), .C(n370), .Y(n2181) );
  AOI22X1 U1593 ( .A(n1144), .B(\data_in<13> ), .C(n1145), .D(\data_in<5> ), 
        .Y(n1150) );
  OAI21X1 U1594 ( .A(n3130), .B(n3341), .C(n369), .Y(n2182) );
  AOI22X1 U1595 ( .A(n1144), .B(\data_in<14> ), .C(n1145), .D(\data_in<6> ), 
        .Y(n1151) );
  OAI21X1 U1596 ( .A(n3130), .B(n3340), .C(n368), .Y(n2183) );
  AOI22X1 U1597 ( .A(n1144), .B(\data_in<15> ), .C(n1145), .D(\data_in<7> ), 
        .Y(n1152) );
  AOI21X1 U1598 ( .A(n2482), .B(n2484), .C(n3176), .Y(n1142) );
  OAI21X1 U1599 ( .A(n3129), .B(n3339), .C(n367), .Y(n2184) );
  AOI22X1 U1600 ( .A(n1156), .B(\data_in<8> ), .C(n1157), .D(\data_in<0> ), 
        .Y(n1155) );
  OAI21X1 U1601 ( .A(n3129), .B(n3338), .C(n366), .Y(n2185) );
  AOI22X1 U1602 ( .A(n1156), .B(\data_in<9> ), .C(n1157), .D(\data_in<1> ), 
        .Y(n1158) );
  OAI21X1 U1603 ( .A(n3129), .B(n3337), .C(n365), .Y(n2186) );
  AOI22X1 U1604 ( .A(n1156), .B(\data_in<10> ), .C(n1157), .D(\data_in<2> ), 
        .Y(n1159) );
  OAI21X1 U1605 ( .A(n3129), .B(n3336), .C(n364), .Y(n2187) );
  AOI22X1 U1606 ( .A(n1156), .B(\data_in<11> ), .C(n1157), .D(\data_in<3> ), 
        .Y(n1160) );
  OAI21X1 U1607 ( .A(n3129), .B(n3335), .C(n363), .Y(n2188) );
  AOI22X1 U1608 ( .A(n1156), .B(\data_in<12> ), .C(n1157), .D(\data_in<4> ), 
        .Y(n1161) );
  OAI21X1 U1609 ( .A(n3129), .B(n3334), .C(n362), .Y(n2189) );
  AOI22X1 U1610 ( .A(n1156), .B(\data_in<13> ), .C(n1157), .D(\data_in<5> ), 
        .Y(n1162) );
  OAI21X1 U1611 ( .A(n3129), .B(n3333), .C(n361), .Y(n2190) );
  AOI22X1 U1612 ( .A(n1156), .B(\data_in<14> ), .C(n1157), .D(\data_in<6> ), 
        .Y(n1163) );
  OAI21X1 U1613 ( .A(n3129), .B(n3332), .C(n360), .Y(n2191) );
  AOI22X1 U1614 ( .A(n1156), .B(\data_in<15> ), .C(n1157), .D(\data_in<7> ), 
        .Y(n1164) );
  AOI21X1 U1615 ( .A(n2484), .B(n2478), .C(n3176), .Y(n1154) );
  OAI21X1 U1616 ( .A(n3128), .B(n3331), .C(n359), .Y(n2192) );
  AOI22X1 U1617 ( .A(n1168), .B(\data_in<8> ), .C(n1169), .D(\data_in<0> ), 
        .Y(n1167) );
  OAI21X1 U1618 ( .A(n3128), .B(n3330), .C(n358), .Y(n2193) );
  AOI22X1 U1619 ( .A(n1168), .B(\data_in<9> ), .C(n1169), .D(\data_in<1> ), 
        .Y(n1170) );
  OAI21X1 U1620 ( .A(n3128), .B(n3329), .C(n357), .Y(n2194) );
  AOI22X1 U1621 ( .A(n1168), .B(\data_in<10> ), .C(n1169), .D(\data_in<2> ), 
        .Y(n1171) );
  OAI21X1 U1622 ( .A(n3128), .B(n3328), .C(n356), .Y(n2195) );
  AOI22X1 U1623 ( .A(n1168), .B(\data_in<11> ), .C(n1169), .D(\data_in<3> ), 
        .Y(n1172) );
  OAI21X1 U1624 ( .A(n3128), .B(n3327), .C(n355), .Y(n2196) );
  AOI22X1 U1625 ( .A(n1168), .B(\data_in<12> ), .C(n1169), .D(\data_in<4> ), 
        .Y(n1173) );
  OAI21X1 U1626 ( .A(n3128), .B(n3326), .C(n354), .Y(n2197) );
  AOI22X1 U1627 ( .A(n1168), .B(\data_in<13> ), .C(n1169), .D(\data_in<5> ), 
        .Y(n1174) );
  OAI21X1 U1628 ( .A(n3128), .B(n3325), .C(n353), .Y(n2198) );
  AOI22X1 U1629 ( .A(n1168), .B(\data_in<14> ), .C(n1169), .D(\data_in<6> ), 
        .Y(n1175) );
  OAI21X1 U1630 ( .A(n3128), .B(n3324), .C(n352), .Y(n2199) );
  AOI22X1 U1631 ( .A(n1168), .B(\data_in<15> ), .C(n1169), .D(\data_in<7> ), 
        .Y(n1176) );
  AOI21X1 U1632 ( .A(n2478), .B(n2480), .C(n3176), .Y(n1166) );
  OAI21X1 U1633 ( .A(n3127), .B(n3323), .C(n351), .Y(n2200) );
  AOI22X1 U1634 ( .A(n1180), .B(\data_in<8> ), .C(n1181), .D(\data_in<0> ), 
        .Y(n1179) );
  OAI21X1 U1635 ( .A(n3127), .B(n3322), .C(n350), .Y(n2201) );
  AOI22X1 U1636 ( .A(n1180), .B(\data_in<9> ), .C(n1181), .D(\data_in<1> ), 
        .Y(n1182) );
  OAI21X1 U1637 ( .A(n3127), .B(n3321), .C(n349), .Y(n2202) );
  AOI22X1 U1638 ( .A(n1180), .B(\data_in<10> ), .C(n1181), .D(\data_in<2> ), 
        .Y(n1183) );
  OAI21X1 U1639 ( .A(n3127), .B(n3320), .C(n348), .Y(n2203) );
  AOI22X1 U1640 ( .A(n1180), .B(\data_in<11> ), .C(n1181), .D(\data_in<3> ), 
        .Y(n1184) );
  OAI21X1 U1641 ( .A(n3127), .B(n3319), .C(n347), .Y(n2204) );
  AOI22X1 U1642 ( .A(n1180), .B(\data_in<12> ), .C(n1181), .D(\data_in<4> ), 
        .Y(n1185) );
  OAI21X1 U1643 ( .A(n3127), .B(n3318), .C(n346), .Y(n2205) );
  AOI22X1 U1644 ( .A(n1180), .B(\data_in<13> ), .C(n1181), .D(\data_in<5> ), 
        .Y(n1186) );
  OAI21X1 U1645 ( .A(n3127), .B(n3317), .C(n345), .Y(n2206) );
  AOI22X1 U1646 ( .A(n1180), .B(\data_in<14> ), .C(n1181), .D(\data_in<6> ), 
        .Y(n1187) );
  OAI21X1 U1647 ( .A(n3127), .B(n3316), .C(n344), .Y(n2207) );
  AOI22X1 U1648 ( .A(n1180), .B(\data_in<15> ), .C(n1181), .D(\data_in<7> ), 
        .Y(n1188) );
  AOI21X1 U1649 ( .A(n2480), .B(n2506), .C(n3176), .Y(n1178) );
  OAI21X1 U1650 ( .A(n3126), .B(n3315), .C(n343), .Y(n2208) );
  AOI22X1 U1651 ( .A(n1192), .B(\data_in<8> ), .C(n1193), .D(\data_in<0> ), 
        .Y(n1191) );
  OAI21X1 U1652 ( .A(n3126), .B(n3314), .C(n342), .Y(n2209) );
  AOI22X1 U1653 ( .A(n1192), .B(\data_in<9> ), .C(n1193), .D(\data_in<1> ), 
        .Y(n1194) );
  OAI21X1 U1654 ( .A(n3126), .B(n3313), .C(n341), .Y(n2210) );
  AOI22X1 U1655 ( .A(n1192), .B(\data_in<10> ), .C(n1193), .D(\data_in<2> ), 
        .Y(n1195) );
  OAI21X1 U1656 ( .A(n3126), .B(n3312), .C(n340), .Y(n2211) );
  AOI22X1 U1657 ( .A(n1192), .B(\data_in<11> ), .C(n1193), .D(\data_in<3> ), 
        .Y(n1196) );
  OAI21X1 U1658 ( .A(n3126), .B(n3311), .C(n339), .Y(n2212) );
  AOI22X1 U1659 ( .A(n1192), .B(\data_in<12> ), .C(n1193), .D(\data_in<4> ), 
        .Y(n1197) );
  OAI21X1 U1660 ( .A(n3126), .B(n3310), .C(n338), .Y(n2213) );
  AOI22X1 U1661 ( .A(n1192), .B(\data_in<13> ), .C(n1193), .D(\data_in<5> ), 
        .Y(n1198) );
  OAI21X1 U1662 ( .A(n3126), .B(n3309), .C(n337), .Y(n2214) );
  AOI22X1 U1663 ( .A(n1192), .B(\data_in<14> ), .C(n1193), .D(\data_in<6> ), 
        .Y(n1199) );
  OAI21X1 U1664 ( .A(n3126), .B(n3308), .C(n336), .Y(n2215) );
  AOI22X1 U1665 ( .A(n1192), .B(\data_in<15> ), .C(n1193), .D(\data_in<7> ), 
        .Y(n1200) );
  AOI21X1 U1666 ( .A(n2506), .B(n2508), .C(n3175), .Y(n1190) );
  OAI21X1 U1667 ( .A(n3125), .B(n3307), .C(n335), .Y(n2216) );
  AOI22X1 U1668 ( .A(n1204), .B(\data_in<8> ), .C(n1205), .D(\data_in<0> ), 
        .Y(n1203) );
  OAI21X1 U1669 ( .A(n3125), .B(n3306), .C(n334), .Y(n2217) );
  AOI22X1 U1670 ( .A(n1204), .B(\data_in<9> ), .C(n1205), .D(\data_in<1> ), 
        .Y(n1206) );
  OAI21X1 U1671 ( .A(n3125), .B(n3305), .C(n333), .Y(n2218) );
  AOI22X1 U1672 ( .A(n1204), .B(\data_in<10> ), .C(n1205), .D(\data_in<2> ), 
        .Y(n1207) );
  OAI21X1 U1673 ( .A(n3125), .B(n3304), .C(n332), .Y(n2219) );
  AOI22X1 U1674 ( .A(n1204), .B(\data_in<11> ), .C(n1205), .D(\data_in<3> ), 
        .Y(n1208) );
  OAI21X1 U1675 ( .A(n3125), .B(n3303), .C(n331), .Y(n2220) );
  AOI22X1 U1676 ( .A(n1204), .B(\data_in<12> ), .C(n1205), .D(\data_in<4> ), 
        .Y(n1209) );
  OAI21X1 U1677 ( .A(n3125), .B(n3302), .C(n330), .Y(n2221) );
  AOI22X1 U1678 ( .A(n1204), .B(\data_in<13> ), .C(n1205), .D(\data_in<5> ), 
        .Y(n1210) );
  OAI21X1 U1679 ( .A(n3125), .B(n3301), .C(n329), .Y(n2222) );
  AOI22X1 U1680 ( .A(n1204), .B(\data_in<14> ), .C(n1205), .D(\data_in<6> ), 
        .Y(n1211) );
  OAI21X1 U1681 ( .A(n3125), .B(n3300), .C(n328), .Y(n2223) );
  AOI22X1 U1682 ( .A(n1204), .B(\data_in<15> ), .C(n1205), .D(\data_in<7> ), 
        .Y(n1212) );
  AOI21X1 U1683 ( .A(n2508), .B(n2502), .C(n3175), .Y(n1202) );
  OAI21X1 U1684 ( .A(n3124), .B(n3299), .C(n327), .Y(n2224) );
  AOI22X1 U1685 ( .A(n1216), .B(\data_in<8> ), .C(n1217), .D(\data_in<0> ), 
        .Y(n1215) );
  OAI21X1 U1686 ( .A(n3124), .B(n3298), .C(n326), .Y(n2225) );
  AOI22X1 U1687 ( .A(n1216), .B(\data_in<9> ), .C(n1217), .D(\data_in<1> ), 
        .Y(n1218) );
  OAI21X1 U1688 ( .A(n3124), .B(n3297), .C(n325), .Y(n2226) );
  AOI22X1 U1689 ( .A(n1216), .B(\data_in<10> ), .C(n1217), .D(\data_in<2> ), 
        .Y(n1219) );
  OAI21X1 U1690 ( .A(n3124), .B(n3296), .C(n324), .Y(n2227) );
  AOI22X1 U1691 ( .A(n1216), .B(\data_in<11> ), .C(n1217), .D(\data_in<3> ), 
        .Y(n1220) );
  OAI21X1 U1692 ( .A(n3124), .B(n3295), .C(n323), .Y(n2228) );
  AOI22X1 U1693 ( .A(n1216), .B(\data_in<12> ), .C(n1217), .D(\data_in<4> ), 
        .Y(n1221) );
  OAI21X1 U1694 ( .A(n3124), .B(n3294), .C(n322), .Y(n2229) );
  AOI22X1 U1695 ( .A(n1216), .B(\data_in<13> ), .C(n1217), .D(\data_in<5> ), 
        .Y(n1222) );
  OAI21X1 U1696 ( .A(n3124), .B(n3293), .C(n321), .Y(n2230) );
  AOI22X1 U1697 ( .A(n1216), .B(\data_in<14> ), .C(n1217), .D(\data_in<6> ), 
        .Y(n1223) );
  OAI21X1 U1698 ( .A(n3124), .B(n3292), .C(n320), .Y(n2231) );
  AOI22X1 U1699 ( .A(n1216), .B(\data_in<15> ), .C(n1217), .D(\data_in<7> ), 
        .Y(n1224) );
  AOI21X1 U1700 ( .A(n2502), .B(n2504), .C(n3175), .Y(n1214) );
  OAI21X1 U1701 ( .A(n3123), .B(n3291), .C(n319), .Y(n2232) );
  AOI22X1 U1702 ( .A(n1228), .B(\data_in<8> ), .C(n1229), .D(\data_in<0> ), 
        .Y(n1227) );
  OAI21X1 U1703 ( .A(n3123), .B(n3290), .C(n318), .Y(n2233) );
  AOI22X1 U1704 ( .A(n1228), .B(\data_in<9> ), .C(n1229), .D(\data_in<1> ), 
        .Y(n1230) );
  OAI21X1 U1705 ( .A(n3123), .B(n3289), .C(n317), .Y(n2234) );
  AOI22X1 U1706 ( .A(n1228), .B(\data_in<10> ), .C(n1229), .D(\data_in<2> ), 
        .Y(n1231) );
  OAI21X1 U1707 ( .A(n3123), .B(n3288), .C(n316), .Y(n2235) );
  AOI22X1 U1708 ( .A(n1228), .B(\data_in<11> ), .C(n1229), .D(\data_in<3> ), 
        .Y(n1232) );
  OAI21X1 U1709 ( .A(n3123), .B(n3287), .C(n315), .Y(n2236) );
  AOI22X1 U1710 ( .A(n1228), .B(\data_in<12> ), .C(n1229), .D(\data_in<4> ), 
        .Y(n1233) );
  OAI21X1 U1711 ( .A(n3123), .B(n3286), .C(n314), .Y(n2237) );
  AOI22X1 U1712 ( .A(n1228), .B(\data_in<13> ), .C(n1229), .D(\data_in<5> ), 
        .Y(n1234) );
  OAI21X1 U1713 ( .A(n3123), .B(n3285), .C(n313), .Y(n2238) );
  AOI22X1 U1714 ( .A(n1228), .B(\data_in<14> ), .C(n1229), .D(\data_in<6> ), 
        .Y(n1235) );
  OAI21X1 U1715 ( .A(n3123), .B(n3284), .C(n312), .Y(n2239) );
  AOI22X1 U1716 ( .A(n1228), .B(\data_in<15> ), .C(n1229), .D(\data_in<7> ), 
        .Y(n1236) );
  AOI21X1 U1717 ( .A(n2504), .B(n2498), .C(n3175), .Y(n1226) );
  OAI21X1 U1718 ( .A(n3122), .B(n3283), .C(n311), .Y(n2240) );
  AOI22X1 U1719 ( .A(n1240), .B(\data_in<8> ), .C(n1241), .D(\data_in<0> ), 
        .Y(n1239) );
  OAI21X1 U1720 ( .A(n3122), .B(n3282), .C(n310), .Y(n2241) );
  AOI22X1 U1721 ( .A(n1240), .B(\data_in<9> ), .C(n1241), .D(\data_in<1> ), 
        .Y(n1242) );
  OAI21X1 U1722 ( .A(n3122), .B(n3281), .C(n309), .Y(n2242) );
  AOI22X1 U1723 ( .A(n1240), .B(\data_in<10> ), .C(n1241), .D(\data_in<2> ), 
        .Y(n1243) );
  OAI21X1 U1724 ( .A(n3122), .B(n3280), .C(n308), .Y(n2243) );
  AOI22X1 U1725 ( .A(n1240), .B(\data_in<11> ), .C(n1241), .D(\data_in<3> ), 
        .Y(n1244) );
  OAI21X1 U1726 ( .A(n3122), .B(n3279), .C(n307), .Y(n2244) );
  AOI22X1 U1727 ( .A(n1240), .B(\data_in<12> ), .C(n1241), .D(\data_in<4> ), 
        .Y(n1245) );
  OAI21X1 U1728 ( .A(n3122), .B(n3278), .C(n306), .Y(n2245) );
  AOI22X1 U1729 ( .A(n1240), .B(\data_in<13> ), .C(n1241), .D(\data_in<5> ), 
        .Y(n1246) );
  OAI21X1 U1730 ( .A(n3122), .B(n3277), .C(n305), .Y(n2246) );
  AOI22X1 U1731 ( .A(n1240), .B(\data_in<14> ), .C(n1241), .D(\data_in<6> ), 
        .Y(n1247) );
  OAI21X1 U1732 ( .A(n3122), .B(n3276), .C(n304), .Y(n2247) );
  AOI22X1 U1733 ( .A(n1240), .B(\data_in<15> ), .C(n1241), .D(\data_in<7> ), 
        .Y(n1248) );
  AOI21X1 U1734 ( .A(n2498), .B(n2500), .C(n3175), .Y(n1238) );
  OAI21X1 U1735 ( .A(n3121), .B(n3275), .C(n303), .Y(n2248) );
  AOI22X1 U1736 ( .A(n1252), .B(\data_in<8> ), .C(n1253), .D(\data_in<0> ), 
        .Y(n1251) );
  OAI21X1 U1737 ( .A(n3121), .B(n3274), .C(n302), .Y(n2249) );
  AOI22X1 U1738 ( .A(n1252), .B(\data_in<9> ), .C(n1253), .D(\data_in<1> ), 
        .Y(n1254) );
  OAI21X1 U1739 ( .A(n3121), .B(n3273), .C(n301), .Y(n2250) );
  AOI22X1 U1740 ( .A(n1252), .B(\data_in<10> ), .C(n1253), .D(\data_in<2> ), 
        .Y(n1255) );
  OAI21X1 U1741 ( .A(n3121), .B(n3272), .C(n300), .Y(n2251) );
  AOI22X1 U1742 ( .A(n1252), .B(\data_in<11> ), .C(n1253), .D(\data_in<3> ), 
        .Y(n1256) );
  OAI21X1 U1743 ( .A(n3121), .B(n3271), .C(n299), .Y(n2252) );
  AOI22X1 U1744 ( .A(n1252), .B(\data_in<12> ), .C(n1253), .D(\data_in<4> ), 
        .Y(n1257) );
  OAI21X1 U1745 ( .A(n3121), .B(n3270), .C(n298), .Y(n2253) );
  AOI22X1 U1746 ( .A(n1252), .B(\data_in<13> ), .C(n1253), .D(\data_in<5> ), 
        .Y(n1258) );
  OAI21X1 U1747 ( .A(n3121), .B(n3269), .C(n297), .Y(n2254) );
  AOI22X1 U1748 ( .A(n1252), .B(\data_in<14> ), .C(n1253), .D(\data_in<6> ), 
        .Y(n1259) );
  OAI21X1 U1749 ( .A(n3121), .B(n3268), .C(n296), .Y(n2255) );
  AOI22X1 U1750 ( .A(n1252), .B(\data_in<15> ), .C(n1253), .D(\data_in<7> ), 
        .Y(n1260) );
  AOI21X1 U1751 ( .A(n2500), .B(n2494), .C(n3175), .Y(n1250) );
  OAI21X1 U1752 ( .A(n3120), .B(n3267), .C(n295), .Y(n2256) );
  AOI22X1 U1753 ( .A(n1264), .B(\data_in<8> ), .C(n1265), .D(\data_in<0> ), 
        .Y(n1263) );
  OAI21X1 U1754 ( .A(n3120), .B(n3266), .C(n294), .Y(n2257) );
  AOI22X1 U1755 ( .A(n1264), .B(\data_in<9> ), .C(n1265), .D(\data_in<1> ), 
        .Y(n1266) );
  OAI21X1 U1756 ( .A(n3120), .B(n3265), .C(n293), .Y(n2258) );
  AOI22X1 U1757 ( .A(n1264), .B(\data_in<10> ), .C(n1265), .D(\data_in<2> ), 
        .Y(n1267) );
  OAI21X1 U1758 ( .A(n3120), .B(n3264), .C(n292), .Y(n2259) );
  AOI22X1 U1759 ( .A(n1264), .B(\data_in<11> ), .C(n1265), .D(\data_in<3> ), 
        .Y(n1268) );
  OAI21X1 U1760 ( .A(n3120), .B(n3263), .C(n291), .Y(n2260) );
  AOI22X1 U1761 ( .A(n1264), .B(\data_in<12> ), .C(n1265), .D(\data_in<4> ), 
        .Y(n1269) );
  OAI21X1 U1762 ( .A(n3120), .B(n3262), .C(n290), .Y(n2261) );
  AOI22X1 U1763 ( .A(n1264), .B(\data_in<13> ), .C(n1265), .D(\data_in<5> ), 
        .Y(n1270) );
  OAI21X1 U1764 ( .A(n3120), .B(n3261), .C(n289), .Y(n2262) );
  AOI22X1 U1765 ( .A(n1264), .B(\data_in<14> ), .C(n1265), .D(\data_in<6> ), 
        .Y(n1271) );
  OAI21X1 U1766 ( .A(n3120), .B(n3260), .C(n288), .Y(n2263) );
  AOI22X1 U1767 ( .A(n1264), .B(\data_in<15> ), .C(n1265), .D(\data_in<7> ), 
        .Y(n1272) );
  AOI21X1 U1768 ( .A(n2494), .B(n2496), .C(n3175), .Y(n1262) );
  OAI21X1 U1769 ( .A(n3119), .B(n3259), .C(n287), .Y(n2264) );
  AOI22X1 U1770 ( .A(n1276), .B(\data_in<8> ), .C(n1277), .D(\data_in<0> ), 
        .Y(n1275) );
  OAI21X1 U1771 ( .A(n3119), .B(n3258), .C(n286), .Y(n2265) );
  AOI22X1 U1772 ( .A(n1276), .B(\data_in<9> ), .C(n1277), .D(\data_in<1> ), 
        .Y(n1278) );
  OAI21X1 U1773 ( .A(n3119), .B(n3257), .C(n285), .Y(n2266) );
  AOI22X1 U1774 ( .A(n1276), .B(\data_in<10> ), .C(n1277), .D(\data_in<2> ), 
        .Y(n1279) );
  OAI21X1 U1775 ( .A(n3119), .B(n3256), .C(n284), .Y(n2267) );
  AOI22X1 U1776 ( .A(n1276), .B(\data_in<11> ), .C(n1277), .D(\data_in<3> ), 
        .Y(n1280) );
  OAI21X1 U1777 ( .A(n3119), .B(n3255), .C(n283), .Y(n2268) );
  AOI22X1 U1778 ( .A(n1276), .B(\data_in<12> ), .C(n1277), .D(\data_in<4> ), 
        .Y(n1281) );
  OAI21X1 U1779 ( .A(n3119), .B(n3254), .C(n282), .Y(n2269) );
  AOI22X1 U1780 ( .A(n1276), .B(\data_in<13> ), .C(n1277), .D(\data_in<5> ), 
        .Y(n1282) );
  OAI21X1 U1781 ( .A(n3119), .B(n3253), .C(n281), .Y(n2270) );
  AOI22X1 U1782 ( .A(n1276), .B(\data_in<14> ), .C(n1277), .D(\data_in<6> ), 
        .Y(n1283) );
  OAI21X1 U1783 ( .A(n3119), .B(n3252), .C(n280), .Y(n2271) );
  AOI22X1 U1784 ( .A(n1276), .B(\data_in<15> ), .C(n1277), .D(\data_in<7> ), 
        .Y(n1284) );
  AOI21X1 U1785 ( .A(n2496), .B(n2516), .C(n3175), .Y(n1274) );
  OAI21X1 U1786 ( .A(n3118), .B(n3251), .C(n279), .Y(n2272) );
  AOI22X1 U1787 ( .A(n1288), .B(\data_in<8> ), .C(n1289), .D(\data_in<0> ), 
        .Y(n1287) );
  OAI21X1 U1788 ( .A(n3118), .B(n3250), .C(n278), .Y(n2273) );
  AOI22X1 U1789 ( .A(n1288), .B(\data_in<9> ), .C(n1289), .D(\data_in<1> ), 
        .Y(n1290) );
  OAI21X1 U1790 ( .A(n3118), .B(n3249), .C(n277), .Y(n2274) );
  AOI22X1 U1791 ( .A(n1288), .B(\data_in<10> ), .C(n1289), .D(\data_in<2> ), 
        .Y(n1291) );
  OAI21X1 U1792 ( .A(n3118), .B(n3248), .C(n276), .Y(n2275) );
  AOI22X1 U1793 ( .A(n1288), .B(\data_in<11> ), .C(n1289), .D(\data_in<3> ), 
        .Y(n1292) );
  OAI21X1 U1794 ( .A(n3118), .B(n3247), .C(n275), .Y(n2276) );
  AOI22X1 U1795 ( .A(n1288), .B(\data_in<12> ), .C(n1289), .D(\data_in<4> ), 
        .Y(n1293) );
  OAI21X1 U1796 ( .A(n3118), .B(n3246), .C(n274), .Y(n2277) );
  AOI22X1 U1797 ( .A(n1288), .B(\data_in<13> ), .C(n1289), .D(\data_in<5> ), 
        .Y(n1294) );
  OAI21X1 U1798 ( .A(n3118), .B(n3245), .C(n273), .Y(n2278) );
  AOI22X1 U1799 ( .A(n1288), .B(\data_in<14> ), .C(n1289), .D(\data_in<6> ), 
        .Y(n1295) );
  OAI21X1 U1800 ( .A(n3118), .B(n3244), .C(n272), .Y(n2279) );
  AOI22X1 U1801 ( .A(n1288), .B(\data_in<15> ), .C(n1289), .D(\data_in<7> ), 
        .Y(n1296) );
  AOI21X1 U1802 ( .A(n2516), .B(n2518), .C(n3175), .Y(n1286) );
  OAI21X1 U1803 ( .A(n3117), .B(n3243), .C(n271), .Y(n2280) );
  AOI22X1 U1804 ( .A(n1300), .B(\data_in<8> ), .C(n1301), .D(\data_in<0> ), 
        .Y(n1299) );
  OAI21X1 U1805 ( .A(n3117), .B(n3242), .C(n270), .Y(n2281) );
  AOI22X1 U1806 ( .A(n1300), .B(\data_in<9> ), .C(n1301), .D(\data_in<1> ), 
        .Y(n1302) );
  OAI21X1 U1807 ( .A(n3117), .B(n3241), .C(n269), .Y(n2282) );
  AOI22X1 U1808 ( .A(n1300), .B(\data_in<10> ), .C(n1301), .D(\data_in<2> ), 
        .Y(n1303) );
  OAI21X1 U1809 ( .A(n3117), .B(n3240), .C(n268), .Y(n2283) );
  AOI22X1 U1810 ( .A(n1300), .B(\data_in<11> ), .C(n1301), .D(\data_in<3> ), 
        .Y(n1304) );
  OAI21X1 U1811 ( .A(n3117), .B(n3239), .C(n267), .Y(n2284) );
  AOI22X1 U1812 ( .A(n1300), .B(\data_in<12> ), .C(n1301), .D(\data_in<4> ), 
        .Y(n1305) );
  OAI21X1 U1813 ( .A(n3117), .B(n3238), .C(n266), .Y(n2285) );
  AOI22X1 U1814 ( .A(n1300), .B(\data_in<13> ), .C(n1301), .D(\data_in<5> ), 
        .Y(n1306) );
  OAI21X1 U1815 ( .A(n3117), .B(n3237), .C(n265), .Y(n2286) );
  AOI22X1 U1816 ( .A(n1300), .B(\data_in<14> ), .C(n1301), .D(\data_in<6> ), 
        .Y(n1307) );
  OAI21X1 U1817 ( .A(n3117), .B(n3236), .C(n264), .Y(n2287) );
  AOI22X1 U1818 ( .A(n1300), .B(\data_in<15> ), .C(n1301), .D(\data_in<7> ), 
        .Y(n1308) );
  AOI21X1 U1819 ( .A(n2518), .B(n2512), .C(n3175), .Y(n1298) );
  OAI21X1 U1820 ( .A(n3116), .B(n3235), .C(n263), .Y(n2288) );
  AOI22X1 U1821 ( .A(n1312), .B(\data_in<8> ), .C(n1313), .D(\data_in<0> ), 
        .Y(n1311) );
  OAI21X1 U1822 ( .A(n3116), .B(n3234), .C(n262), .Y(n2289) );
  AOI22X1 U1823 ( .A(n1312), .B(\data_in<9> ), .C(n1313), .D(\data_in<1> ), 
        .Y(n1314) );
  OAI21X1 U1824 ( .A(n3116), .B(n3233), .C(n261), .Y(n2290) );
  AOI22X1 U1825 ( .A(n1312), .B(\data_in<10> ), .C(n1313), .D(\data_in<2> ), 
        .Y(n1315) );
  OAI21X1 U1826 ( .A(n3116), .B(n3232), .C(n260), .Y(n2291) );
  AOI22X1 U1827 ( .A(n1312), .B(\data_in<11> ), .C(n1313), .D(\data_in<3> ), 
        .Y(n1316) );
  OAI21X1 U1828 ( .A(n3116), .B(n3231), .C(n259), .Y(n2292) );
  AOI22X1 U1829 ( .A(n1312), .B(\data_in<12> ), .C(n1313), .D(\data_in<4> ), 
        .Y(n1317) );
  OAI21X1 U1830 ( .A(n3116), .B(n3230), .C(n258), .Y(n2293) );
  AOI22X1 U1831 ( .A(n1312), .B(\data_in<13> ), .C(n1313), .D(\data_in<5> ), 
        .Y(n1318) );
  OAI21X1 U1832 ( .A(n3116), .B(n3229), .C(n257), .Y(n2294) );
  AOI22X1 U1833 ( .A(n1312), .B(\data_in<14> ), .C(n1313), .D(\data_in<6> ), 
        .Y(n1319) );
  OAI21X1 U1834 ( .A(n3116), .B(n3228), .C(n256), .Y(n2295) );
  AOI22X1 U1835 ( .A(n1312), .B(\data_in<15> ), .C(n1313), .D(\data_in<7> ), 
        .Y(n1320) );
  AOI21X1 U1836 ( .A(n2512), .B(n2514), .C(n3175), .Y(n1310) );
  OAI21X1 U1837 ( .A(n3115), .B(n3227), .C(n255), .Y(n2296) );
  AOI22X1 U1838 ( .A(n1324), .B(\data_in<8> ), .C(n1325), .D(\data_in<0> ), 
        .Y(n1323) );
  OAI21X1 U1839 ( .A(n3115), .B(n3226), .C(n254), .Y(n2297) );
  AOI22X1 U1840 ( .A(n1324), .B(\data_in<9> ), .C(n1325), .D(\data_in<1> ), 
        .Y(n1326) );
  OAI21X1 U1841 ( .A(n3115), .B(n3225), .C(n253), .Y(n2298) );
  AOI22X1 U1842 ( .A(n1324), .B(\data_in<10> ), .C(n1325), .D(\data_in<2> ), 
        .Y(n1327) );
  OAI21X1 U1843 ( .A(n3115), .B(n3224), .C(n252), .Y(n2299) );
  AOI22X1 U1844 ( .A(n1324), .B(\data_in<11> ), .C(n1325), .D(\data_in<3> ), 
        .Y(n1328) );
  OAI21X1 U1845 ( .A(n3115), .B(n3223), .C(n251), .Y(n2300) );
  AOI22X1 U1846 ( .A(n1324), .B(\data_in<12> ), .C(n1325), .D(\data_in<4> ), 
        .Y(n1329) );
  OAI21X1 U1847 ( .A(n3115), .B(n3222), .C(n250), .Y(n2301) );
  AOI22X1 U1848 ( .A(n1324), .B(\data_in<13> ), .C(n1325), .D(\data_in<5> ), 
        .Y(n1330) );
  OAI21X1 U1849 ( .A(n3115), .B(n3221), .C(n249), .Y(n2302) );
  AOI22X1 U1850 ( .A(n1324), .B(\data_in<14> ), .C(n1325), .D(\data_in<6> ), 
        .Y(n1331) );
  OAI21X1 U1851 ( .A(n3115), .B(n3220), .C(n248), .Y(n2303) );
  AOI22X1 U1852 ( .A(n1324), .B(\data_in<15> ), .C(n1325), .D(\data_in<7> ), 
        .Y(n1332) );
  AOI21X1 U1853 ( .A(n2514), .B(n2510), .C(n3175), .Y(n1322) );
  OAI21X1 U1854 ( .A(n3114), .B(n3219), .C(n247), .Y(n2304) );
  AOI22X1 U1855 ( .A(n1336), .B(\data_in<8> ), .C(n1337), .D(\data_in<0> ), 
        .Y(n1335) );
  OAI21X1 U1856 ( .A(n3114), .B(n3218), .C(n246), .Y(n2305) );
  AOI22X1 U1857 ( .A(n1336), .B(\data_in<9> ), .C(n1337), .D(\data_in<1> ), 
        .Y(n1338) );
  OAI21X1 U1858 ( .A(n3114), .B(n3217), .C(n245), .Y(n2306) );
  AOI22X1 U1859 ( .A(n1336), .B(\data_in<10> ), .C(n1337), .D(\data_in<2> ), 
        .Y(n1339) );
  OAI21X1 U1860 ( .A(n3114), .B(n3216), .C(n244), .Y(n2307) );
  AOI22X1 U1861 ( .A(n1336), .B(\data_in<11> ), .C(n1337), .D(\data_in<3> ), 
        .Y(n1340) );
  OAI21X1 U1862 ( .A(n3114), .B(n3215), .C(n243), .Y(n2308) );
  AOI22X1 U1863 ( .A(n1336), .B(\data_in<12> ), .C(n1337), .D(\data_in<4> ), 
        .Y(n1341) );
  OAI21X1 U1864 ( .A(n3114), .B(n3214), .C(n242), .Y(n2309) );
  AOI22X1 U1865 ( .A(n1336), .B(\data_in<13> ), .C(n1337), .D(\data_in<5> ), 
        .Y(n1342) );
  OAI21X1 U1866 ( .A(n3114), .B(n3213), .C(n241), .Y(n2310) );
  AOI22X1 U1867 ( .A(n1336), .B(\data_in<14> ), .C(n1337), .D(\data_in<6> ), 
        .Y(n1343) );
  OAI21X1 U1868 ( .A(n3114), .B(n3212), .C(n240), .Y(n2311) );
  AOI22X1 U1869 ( .A(n1336), .B(\data_in<15> ), .C(n1337), .D(\data_in<7> ), 
        .Y(n1344) );
  AOI21X1 U1870 ( .A(n2510), .B(n2582), .C(n3175), .Y(n1334) );
  OAI21X1 U1871 ( .A(n3113), .B(n3211), .C(n239), .Y(n2312) );
  AOI22X1 U1872 ( .A(n1348), .B(\data_in<8> ), .C(n1349), .D(\data_in<0> ), 
        .Y(n1347) );
  OAI21X1 U1873 ( .A(n3113), .B(n3210), .C(n238), .Y(n2313) );
  AOI22X1 U1874 ( .A(n1348), .B(\data_in<9> ), .C(n1349), .D(\data_in<1> ), 
        .Y(n1350) );
  OAI21X1 U1875 ( .A(n3113), .B(n3209), .C(n237), .Y(n2314) );
  AOI22X1 U1876 ( .A(n1348), .B(\data_in<10> ), .C(n1349), .D(\data_in<2> ), 
        .Y(n1351) );
  OAI21X1 U1877 ( .A(n3113), .B(n3208), .C(n236), .Y(n2315) );
  AOI22X1 U1878 ( .A(n1348), .B(\data_in<11> ), .C(n1349), .D(\data_in<3> ), 
        .Y(n1352) );
  OAI21X1 U1879 ( .A(n3113), .B(n3207), .C(n235), .Y(n2316) );
  AOI22X1 U1880 ( .A(n1348), .B(\data_in<12> ), .C(n1349), .D(\data_in<4> ), 
        .Y(n1353) );
  OAI21X1 U1881 ( .A(n3113), .B(n3206), .C(n234), .Y(n2317) );
  AOI22X1 U1882 ( .A(n1348), .B(\data_in<13> ), .C(n1349), .D(\data_in<5> ), 
        .Y(n1354) );
  OAI21X1 U1883 ( .A(n3113), .B(n3205), .C(n233), .Y(n2318) );
  AOI22X1 U1884 ( .A(n1348), .B(\data_in<14> ), .C(n1349), .D(\data_in<6> ), 
        .Y(n1355) );
  OAI21X1 U1885 ( .A(n3113), .B(n3204), .C(n232), .Y(n2319) );
  AOI22X1 U1886 ( .A(n1348), .B(\data_in<15> ), .C(n1349), .D(\data_in<7> ), 
        .Y(n1356) );
  OAI21X1 U1887 ( .A(n3175), .B(n2582), .C(n2458), .Y(n1346) );
  OAI21X1 U1888 ( .A(n2457), .B(n3203), .C(n2338), .Y(n2320) );
  OAI21X1 U1890 ( .A(n2457), .B(n3202), .C(n2336), .Y(n2321) );
  OAI21X1 U1892 ( .A(n2457), .B(n3201), .C(n2334), .Y(n2322) );
  OAI21X1 U1894 ( .A(n2457), .B(n3200), .C(n2332), .Y(n2323) );
  OAI21X1 U1896 ( .A(n2457), .B(n3199), .C(n2330), .Y(n2324) );
  OAI21X1 U1898 ( .A(n2457), .B(n3198), .C(n2328), .Y(n2325) );
  OAI21X1 U1900 ( .A(n2457), .B(n3197), .C(n1796), .Y(n2326) );
  OAI21X1 U1902 ( .A(n2457), .B(n3196), .C(n1794), .Y(n2327) );
  NAND3X1 U1905 ( .A(enable), .B(n3186), .C(wr), .Y(n625) );
  AOI21X1 U1906 ( .A(n1367), .B(n1368), .C(n2451), .Y(n3709) );
  NOR3X1 U1907 ( .A(n1370), .B(n180), .C(n188), .Y(n1368) );
  AOI22X1 U1909 ( .A(\mem<55><7> ), .B(n2577), .C(\mem<54><7> ), .D(n2579), 
        .Y(n1377) );
  AOI22X1 U1910 ( .A(\mem<53><7> ), .B(n2573), .C(\mem<52><7> ), .D(n2575), 
        .Y(n1376) );
  AOI22X1 U1911 ( .A(\mem<51><7> ), .B(n2569), .C(\mem<50><7> ), .D(n2571), 
        .Y(n1374) );
  AOI22X1 U1912 ( .A(\mem<49><7> ), .B(n2565), .C(\mem<48><7> ), .D(n2567), 
        .Y(n1373) );
  AOI22X1 U1914 ( .A(\mem<63><7> ), .B(n2459), .C(\mem<62><7> ), .D(n2563), 
        .Y(n1382) );
  AOI22X1 U1915 ( .A(\mem<61><7> ), .B(n2559), .C(\mem<60><7> ), .D(n2561), 
        .Y(n1381) );
  AOI22X1 U1916 ( .A(\mem<59><7> ), .B(n2555), .C(\mem<58><7> ), .D(n2557), 
        .Y(n1379) );
  AOI22X1 U1917 ( .A(\mem<57><7> ), .B(n2551), .C(\mem<56><7> ), .D(n2553), 
        .Y(n1378) );
  AOI22X1 U1919 ( .A(\mem<39><7> ), .B(n2547), .C(\mem<38><7> ), .D(n2549), 
        .Y(n1389) );
  AOI22X1 U1920 ( .A(\mem<37><7> ), .B(n2543), .C(\mem<36><7> ), .D(n2545), 
        .Y(n1388) );
  AOI22X1 U1921 ( .A(\mem<35><7> ), .B(n2539), .C(\mem<34><7> ), .D(n2541), 
        .Y(n1386) );
  AOI22X1 U1922 ( .A(\mem<33><7> ), .B(n2536), .C(\mem<32><7> ), .D(n2537), 
        .Y(n1385) );
  AOI22X1 U1924 ( .A(\mem<47><7> ), .B(n2531), .C(\mem<46><7> ), .D(n2533), 
        .Y(n1394) );
  AOI22X1 U1925 ( .A(\mem<45><7> ), .B(n2527), .C(\mem<44><7> ), .D(n2529), 
        .Y(n1393) );
  AOI22X1 U1926 ( .A(\mem<43><7> ), .B(n2523), .C(\mem<42><7> ), .D(n2525), 
        .Y(n1391) );
  AOI22X1 U1927 ( .A(\mem<41><7> ), .B(n2519), .C(\mem<40><7> ), .D(n2521), 
        .Y(n1390) );
  NOR3X1 U1928 ( .A(n1395), .B(n179), .C(n229), .Y(n1367) );
  AOI22X1 U1930 ( .A(\mem<7><7> ), .B(n2515), .C(\mem<6><7> ), .D(n2517), .Y(
        n1402) );
  AOI22X1 U1931 ( .A(\mem<5><7> ), .B(n2511), .C(\mem<4><7> ), .D(n2513), .Y(
        n1401) );
  AOI22X1 U1932 ( .A(\mem<3><7> ), .B(n2509), .C(\mem<2><7> ), .D(n2581), .Y(
        n1399) );
  AOI22X1 U1933 ( .A(\mem<1><7> ), .B(n2455), .C(n1403), .D(\mem<0><7> ), .Y(
        n1398) );
  AOI22X1 U1935 ( .A(\mem<15><7> ), .B(n2505), .C(\mem<14><7> ), .D(n2507), 
        .Y(n1408) );
  AOI22X1 U1936 ( .A(\mem<13><7> ), .B(n2501), .C(\mem<12><7> ), .D(n2503), 
        .Y(n1407) );
  AOI22X1 U1937 ( .A(\mem<11><7> ), .B(n2497), .C(\mem<10><7> ), .D(n2499), 
        .Y(n1405) );
  AOI22X1 U1938 ( .A(\mem<9><7> ), .B(n2493), .C(\mem<8><7> ), .D(n2495), .Y(
        n1404) );
  AOI22X1 U1940 ( .A(\mem<23><7> ), .B(n2489), .C(\mem<22><7> ), .D(n2491), 
        .Y(n1415) );
  AOI22X1 U1941 ( .A(\mem<21><7> ), .B(n2485), .C(\mem<20><7> ), .D(n2487), 
        .Y(n1414) );
  AOI22X1 U1942 ( .A(\mem<19><7> ), .B(n2481), .C(\mem<18><7> ), .D(n2483), 
        .Y(n1412) );
  AOI22X1 U1943 ( .A(\mem<17><7> ), .B(n2477), .C(\mem<16><7> ), .D(n2479), 
        .Y(n1411) );
  AOI22X1 U1945 ( .A(\mem<31><7> ), .B(n2473), .C(\mem<30><7> ), .D(n2475), 
        .Y(n1420) );
  AOI22X1 U1946 ( .A(\mem<29><7> ), .B(n2469), .C(\mem<28><7> ), .D(n2471), 
        .Y(n1419) );
  AOI22X1 U1947 ( .A(\mem<27><7> ), .B(n2465), .C(\mem<26><7> ), .D(n2467), 
        .Y(n1417) );
  AOI22X1 U1948 ( .A(\mem<25><7> ), .B(n2461), .C(\mem<24><7> ), .D(n2463), 
        .Y(n1416) );
  AOI21X1 U1949 ( .A(n1421), .B(n1422), .C(n2451), .Y(n3710) );
  NOR3X1 U1950 ( .A(n1423), .B(n178), .C(n187), .Y(n1422) );
  AOI22X1 U1952 ( .A(\mem<55><6> ), .B(n2577), .C(\mem<54><6> ), .D(n2579), 
        .Y(n1430) );
  AOI22X1 U1953 ( .A(\mem<53><6> ), .B(n2573), .C(\mem<52><6> ), .D(n2575), 
        .Y(n1429) );
  AOI22X1 U1954 ( .A(\mem<51><6> ), .B(n2569), .C(\mem<50><6> ), .D(n2571), 
        .Y(n1427) );
  AOI22X1 U1955 ( .A(\mem<49><6> ), .B(n2565), .C(\mem<48><6> ), .D(n2567), 
        .Y(n1426) );
  AOI22X1 U1957 ( .A(\mem<63><6> ), .B(n2459), .C(\mem<62><6> ), .D(n2563), 
        .Y(n1435) );
  AOI22X1 U1958 ( .A(\mem<61><6> ), .B(n2559), .C(\mem<60><6> ), .D(n2561), 
        .Y(n1434) );
  AOI22X1 U1959 ( .A(\mem<59><6> ), .B(n2555), .C(\mem<58><6> ), .D(n2557), 
        .Y(n1432) );
  AOI22X1 U1960 ( .A(\mem<57><6> ), .B(n2551), .C(\mem<56><6> ), .D(n2553), 
        .Y(n1431) );
  AOI22X1 U1962 ( .A(\mem<39><6> ), .B(n2547), .C(\mem<38><6> ), .D(n2549), 
        .Y(n1442) );
  AOI22X1 U1963 ( .A(\mem<37><6> ), .B(n2543), .C(\mem<36><6> ), .D(n2545), 
        .Y(n1441) );
  AOI22X1 U1964 ( .A(\mem<35><6> ), .B(n2539), .C(\mem<34><6> ), .D(n2541), 
        .Y(n1439) );
  AOI22X1 U1965 ( .A(\mem<33><6> ), .B(n2536), .C(\mem<32><6> ), .D(n2537), 
        .Y(n1438) );
  AOI22X1 U1967 ( .A(\mem<47><6> ), .B(n2531), .C(\mem<46><6> ), .D(n2533), 
        .Y(n1447) );
  AOI22X1 U1968 ( .A(\mem<45><6> ), .B(n2527), .C(\mem<44><6> ), .D(n2529), 
        .Y(n1446) );
  AOI22X1 U1969 ( .A(\mem<43><6> ), .B(n2523), .C(\mem<42><6> ), .D(n2525), 
        .Y(n1444) );
  AOI22X1 U1970 ( .A(\mem<41><6> ), .B(n2519), .C(\mem<40><6> ), .D(n2521), 
        .Y(n1443) );
  NOR3X1 U1971 ( .A(n1448), .B(n177), .C(n226), .Y(n1421) );
  AOI22X1 U1973 ( .A(\mem<7><6> ), .B(n2515), .C(\mem<6><6> ), .D(n2517), .Y(
        n1455) );
  AOI22X1 U1974 ( .A(\mem<5><6> ), .B(n2511), .C(\mem<4><6> ), .D(n2513), .Y(
        n1454) );
  AOI22X1 U1975 ( .A(\mem<3><6> ), .B(n2509), .C(\mem<2><6> ), .D(n2581), .Y(
        n1452) );
  AOI22X1 U1976 ( .A(\mem<1><6> ), .B(n2455), .C(n1403), .D(\mem<0><6> ), .Y(
        n1451) );
  AOI22X1 U1978 ( .A(\mem<15><6> ), .B(n2505), .C(\mem<14><6> ), .D(n2507), 
        .Y(n1460) );
  AOI22X1 U1979 ( .A(\mem<13><6> ), .B(n2501), .C(\mem<12><6> ), .D(n2503), 
        .Y(n1459) );
  AOI22X1 U1980 ( .A(\mem<11><6> ), .B(n2497), .C(\mem<10><6> ), .D(n2499), 
        .Y(n1457) );
  AOI22X1 U1981 ( .A(\mem<9><6> ), .B(n2493), .C(\mem<8><6> ), .D(n2495), .Y(
        n1456) );
  AOI22X1 U1983 ( .A(\mem<23><6> ), .B(n2489), .C(\mem<22><6> ), .D(n2491), 
        .Y(n1467) );
  AOI22X1 U1984 ( .A(\mem<21><6> ), .B(n2485), .C(\mem<20><6> ), .D(n2487), 
        .Y(n1466) );
  AOI22X1 U1985 ( .A(\mem<19><6> ), .B(n2481), .C(\mem<18><6> ), .D(n2483), 
        .Y(n1464) );
  AOI22X1 U1986 ( .A(\mem<17><6> ), .B(n2477), .C(\mem<16><6> ), .D(n2479), 
        .Y(n1463) );
  AOI22X1 U1988 ( .A(\mem<31><6> ), .B(n2473), .C(\mem<30><6> ), .D(n2475), 
        .Y(n1472) );
  AOI22X1 U1989 ( .A(\mem<29><6> ), .B(n2469), .C(\mem<28><6> ), .D(n2471), 
        .Y(n1471) );
  AOI22X1 U1990 ( .A(\mem<27><6> ), .B(n2465), .C(\mem<26><6> ), .D(n2467), 
        .Y(n1469) );
  AOI22X1 U1991 ( .A(\mem<25><6> ), .B(n2461), .C(\mem<24><6> ), .D(n2463), 
        .Y(n1468) );
  AOI21X1 U1992 ( .A(n1473), .B(n1474), .C(n2451), .Y(n3711) );
  NOR3X1 U1993 ( .A(n1475), .B(n176), .C(n186), .Y(n1474) );
  AOI22X1 U1995 ( .A(\mem<55><5> ), .B(n2577), .C(\mem<54><5> ), .D(n2579), 
        .Y(n1482) );
  AOI22X1 U1996 ( .A(\mem<53><5> ), .B(n2573), .C(\mem<52><5> ), .D(n2575), 
        .Y(n1481) );
  AOI22X1 U1997 ( .A(\mem<51><5> ), .B(n2569), .C(\mem<50><5> ), .D(n2571), 
        .Y(n1479) );
  AOI22X1 U1998 ( .A(\mem<49><5> ), .B(n2565), .C(\mem<48><5> ), .D(n2567), 
        .Y(n1478) );
  AOI22X1 U2000 ( .A(\mem<63><5> ), .B(n2459), .C(\mem<62><5> ), .D(n2563), 
        .Y(n1487) );
  AOI22X1 U2001 ( .A(\mem<61><5> ), .B(n2559), .C(\mem<60><5> ), .D(n2561), 
        .Y(n1486) );
  AOI22X1 U2002 ( .A(\mem<59><5> ), .B(n2555), .C(\mem<58><5> ), .D(n2557), 
        .Y(n1484) );
  AOI22X1 U2003 ( .A(\mem<57><5> ), .B(n2551), .C(\mem<56><5> ), .D(n2553), 
        .Y(n1483) );
  AOI22X1 U2005 ( .A(\mem<39><5> ), .B(n2547), .C(\mem<38><5> ), .D(n2549), 
        .Y(n1494) );
  AOI22X1 U2006 ( .A(\mem<37><5> ), .B(n2543), .C(\mem<36><5> ), .D(n2545), 
        .Y(n1493) );
  AOI22X1 U2007 ( .A(\mem<35><5> ), .B(n2539), .C(\mem<34><5> ), .D(n2541), 
        .Y(n1491) );
  AOI22X1 U2008 ( .A(\mem<33><5> ), .B(n2536), .C(\mem<32><5> ), .D(n2537), 
        .Y(n1490) );
  AOI22X1 U2010 ( .A(\mem<47><5> ), .B(n2531), .C(\mem<46><5> ), .D(n2533), 
        .Y(n1499) );
  AOI22X1 U2011 ( .A(\mem<45><5> ), .B(n2527), .C(\mem<44><5> ), .D(n2529), 
        .Y(n1498) );
  AOI22X1 U2012 ( .A(\mem<43><5> ), .B(n2523), .C(\mem<42><5> ), .D(n2525), 
        .Y(n1496) );
  AOI22X1 U2013 ( .A(\mem<41><5> ), .B(n2519), .C(\mem<40><5> ), .D(n2521), 
        .Y(n1495) );
  NOR3X1 U2014 ( .A(n1500), .B(n175), .C(n223), .Y(n1473) );
  AOI22X1 U2016 ( .A(\mem<7><5> ), .B(n2515), .C(\mem<6><5> ), .D(n2517), .Y(
        n1507) );
  AOI22X1 U2017 ( .A(\mem<5><5> ), .B(n2511), .C(\mem<4><5> ), .D(n2513), .Y(
        n1506) );
  AOI22X1 U2018 ( .A(\mem<3><5> ), .B(n2509), .C(\mem<2><5> ), .D(n2581), .Y(
        n1504) );
  AOI22X1 U2019 ( .A(\mem<1><5> ), .B(n2455), .C(n1403), .D(\mem<0><5> ), .Y(
        n1503) );
  AOI22X1 U2021 ( .A(\mem<15><5> ), .B(n2505), .C(\mem<14><5> ), .D(n2507), 
        .Y(n1512) );
  AOI22X1 U2022 ( .A(\mem<13><5> ), .B(n2501), .C(\mem<12><5> ), .D(n2503), 
        .Y(n1511) );
  AOI22X1 U2023 ( .A(\mem<11><5> ), .B(n2497), .C(\mem<10><5> ), .D(n2499), 
        .Y(n1509) );
  AOI22X1 U2024 ( .A(\mem<9><5> ), .B(n2493), .C(\mem<8><5> ), .D(n2495), .Y(
        n1508) );
  AOI22X1 U2026 ( .A(\mem<23><5> ), .B(n2489), .C(\mem<22><5> ), .D(n2491), 
        .Y(n1519) );
  AOI22X1 U2027 ( .A(\mem<21><5> ), .B(n2485), .C(\mem<20><5> ), .D(n2487), 
        .Y(n1518) );
  AOI22X1 U2028 ( .A(\mem<19><5> ), .B(n2481), .C(\mem<18><5> ), .D(n2483), 
        .Y(n1516) );
  AOI22X1 U2029 ( .A(\mem<17><5> ), .B(n2477), .C(\mem<16><5> ), .D(n2479), 
        .Y(n1515) );
  AOI22X1 U2031 ( .A(\mem<31><5> ), .B(n2473), .C(\mem<30><5> ), .D(n2475), 
        .Y(n1524) );
  AOI22X1 U2032 ( .A(\mem<29><5> ), .B(n2469), .C(\mem<28><5> ), .D(n2471), 
        .Y(n1523) );
  AOI22X1 U2033 ( .A(\mem<27><5> ), .B(n2465), .C(\mem<26><5> ), .D(n2467), 
        .Y(n1521) );
  AOI22X1 U2034 ( .A(\mem<25><5> ), .B(n2461), .C(\mem<24><5> ), .D(n2463), 
        .Y(n1520) );
  AOI21X1 U2035 ( .A(n1525), .B(n1526), .C(n2451), .Y(n3712) );
  NOR3X1 U2036 ( .A(n1527), .B(n174), .C(n185), .Y(n1526) );
  AOI22X1 U2038 ( .A(\mem<55><4> ), .B(n2577), .C(\mem<54><4> ), .D(n2579), 
        .Y(n1534) );
  AOI22X1 U2039 ( .A(\mem<53><4> ), .B(n2573), .C(\mem<52><4> ), .D(n2575), 
        .Y(n1533) );
  AOI22X1 U2040 ( .A(\mem<51><4> ), .B(n2569), .C(\mem<50><4> ), .D(n2571), 
        .Y(n1531) );
  AOI22X1 U2041 ( .A(\mem<49><4> ), .B(n2565), .C(\mem<48><4> ), .D(n2567), 
        .Y(n1530) );
  AOI22X1 U2043 ( .A(\mem<63><4> ), .B(n2459), .C(\mem<62><4> ), .D(n2563), 
        .Y(n1539) );
  AOI22X1 U2044 ( .A(\mem<61><4> ), .B(n2559), .C(\mem<60><4> ), .D(n2561), 
        .Y(n1538) );
  AOI22X1 U2045 ( .A(\mem<59><4> ), .B(n2555), .C(\mem<58><4> ), .D(n2557), 
        .Y(n1536) );
  AOI22X1 U2046 ( .A(\mem<57><4> ), .B(n2551), .C(\mem<56><4> ), .D(n2553), 
        .Y(n1535) );
  AOI22X1 U2048 ( .A(\mem<39><4> ), .B(n2547), .C(\mem<38><4> ), .D(n2549), 
        .Y(n1546) );
  AOI22X1 U2049 ( .A(\mem<37><4> ), .B(n2543), .C(\mem<36><4> ), .D(n2545), 
        .Y(n1545) );
  AOI22X1 U2050 ( .A(\mem<35><4> ), .B(n2539), .C(\mem<34><4> ), .D(n2541), 
        .Y(n1543) );
  AOI22X1 U2051 ( .A(\mem<33><4> ), .B(n2536), .C(\mem<32><4> ), .D(n2537), 
        .Y(n1542) );
  AOI22X1 U2053 ( .A(\mem<47><4> ), .B(n2531), .C(\mem<46><4> ), .D(n2533), 
        .Y(n1551) );
  AOI22X1 U2054 ( .A(\mem<45><4> ), .B(n2527), .C(\mem<44><4> ), .D(n2529), 
        .Y(n1550) );
  AOI22X1 U2055 ( .A(\mem<43><4> ), .B(n2523), .C(\mem<42><4> ), .D(n2525), 
        .Y(n1548) );
  AOI22X1 U2056 ( .A(\mem<41><4> ), .B(n2519), .C(\mem<40><4> ), .D(n2521), 
        .Y(n1547) );
  NOR3X1 U2057 ( .A(n1552), .B(n173), .C(n220), .Y(n1525) );
  AOI22X1 U2059 ( .A(\mem<7><4> ), .B(n2515), .C(\mem<6><4> ), .D(n2517), .Y(
        n1559) );
  AOI22X1 U2060 ( .A(\mem<5><4> ), .B(n2511), .C(\mem<4><4> ), .D(n2513), .Y(
        n1558) );
  AOI22X1 U2061 ( .A(\mem<3><4> ), .B(n2509), .C(\mem<2><4> ), .D(n2581), .Y(
        n1556) );
  AOI22X1 U2062 ( .A(\mem<1><4> ), .B(n2455), .C(n1403), .D(\mem<0><4> ), .Y(
        n1555) );
  AOI22X1 U2064 ( .A(\mem<15><4> ), .B(n2505), .C(\mem<14><4> ), .D(n2507), 
        .Y(n1564) );
  AOI22X1 U2065 ( .A(\mem<13><4> ), .B(n2501), .C(\mem<12><4> ), .D(n2503), 
        .Y(n1563) );
  AOI22X1 U2066 ( .A(\mem<11><4> ), .B(n2497), .C(\mem<10><4> ), .D(n2499), 
        .Y(n1561) );
  AOI22X1 U2067 ( .A(\mem<9><4> ), .B(n2493), .C(\mem<8><4> ), .D(n2495), .Y(
        n1560) );
  AOI22X1 U2069 ( .A(\mem<23><4> ), .B(n2489), .C(\mem<22><4> ), .D(n2491), 
        .Y(n1571) );
  AOI22X1 U2070 ( .A(\mem<21><4> ), .B(n2485), .C(\mem<20><4> ), .D(n2487), 
        .Y(n1570) );
  AOI22X1 U2071 ( .A(\mem<19><4> ), .B(n2481), .C(\mem<18><4> ), .D(n2483), 
        .Y(n1568) );
  AOI22X1 U2072 ( .A(\mem<17><4> ), .B(n2477), .C(\mem<16><4> ), .D(n2479), 
        .Y(n1567) );
  AOI22X1 U2074 ( .A(\mem<31><4> ), .B(n2473), .C(\mem<30><4> ), .D(n2475), 
        .Y(n1576) );
  AOI22X1 U2075 ( .A(\mem<29><4> ), .B(n2469), .C(\mem<28><4> ), .D(n2471), 
        .Y(n1575) );
  AOI22X1 U2076 ( .A(\mem<27><4> ), .B(n2465), .C(\mem<26><4> ), .D(n2467), 
        .Y(n1573) );
  AOI22X1 U2077 ( .A(\mem<25><4> ), .B(n2461), .C(\mem<24><4> ), .D(n2463), 
        .Y(n1572) );
  AOI21X1 U2078 ( .A(n1577), .B(n1578), .C(n2451), .Y(n3713) );
  NOR3X1 U2079 ( .A(n1579), .B(n172), .C(n184), .Y(n1578) );
  AOI22X1 U2081 ( .A(\mem<55><3> ), .B(n2577), .C(\mem<54><3> ), .D(n2579), 
        .Y(n1586) );
  AOI22X1 U2082 ( .A(\mem<53><3> ), .B(n2573), .C(\mem<52><3> ), .D(n2575), 
        .Y(n1585) );
  AOI22X1 U2083 ( .A(\mem<51><3> ), .B(n2569), .C(\mem<50><3> ), .D(n2571), 
        .Y(n1583) );
  AOI22X1 U2084 ( .A(\mem<49><3> ), .B(n2565), .C(\mem<48><3> ), .D(n2567), 
        .Y(n1582) );
  AOI22X1 U2086 ( .A(\mem<63><3> ), .B(n2459), .C(\mem<62><3> ), .D(n2563), 
        .Y(n1591) );
  AOI22X1 U2087 ( .A(\mem<61><3> ), .B(n2559), .C(\mem<60><3> ), .D(n2561), 
        .Y(n1590) );
  AOI22X1 U2088 ( .A(\mem<59><3> ), .B(n2555), .C(\mem<58><3> ), .D(n2557), 
        .Y(n1588) );
  AOI22X1 U2089 ( .A(\mem<57><3> ), .B(n2551), .C(\mem<56><3> ), .D(n2553), 
        .Y(n1587) );
  AOI22X1 U2091 ( .A(\mem<39><3> ), .B(n2547), .C(\mem<38><3> ), .D(n2549), 
        .Y(n1598) );
  AOI22X1 U2092 ( .A(\mem<37><3> ), .B(n2543), .C(\mem<36><3> ), .D(n2545), 
        .Y(n1597) );
  AOI22X1 U2093 ( .A(\mem<35><3> ), .B(n2539), .C(\mem<34><3> ), .D(n2541), 
        .Y(n1595) );
  AOI22X1 U2094 ( .A(\mem<33><3> ), .B(n2536), .C(\mem<32><3> ), .D(n2537), 
        .Y(n1594) );
  AOI22X1 U2096 ( .A(\mem<47><3> ), .B(n2531), .C(\mem<46><3> ), .D(n2533), 
        .Y(n1603) );
  AOI22X1 U2097 ( .A(\mem<45><3> ), .B(n2527), .C(\mem<44><3> ), .D(n2529), 
        .Y(n1602) );
  AOI22X1 U2098 ( .A(\mem<43><3> ), .B(n2523), .C(\mem<42><3> ), .D(n2525), 
        .Y(n1600) );
  AOI22X1 U2099 ( .A(\mem<41><3> ), .B(n2519), .C(\mem<40><3> ), .D(n2521), 
        .Y(n1599) );
  NOR3X1 U2100 ( .A(n1604), .B(n171), .C(n217), .Y(n1577) );
  AOI22X1 U2102 ( .A(\mem<7><3> ), .B(n2515), .C(\mem<6><3> ), .D(n2517), .Y(
        n1611) );
  AOI22X1 U2103 ( .A(\mem<5><3> ), .B(n2511), .C(\mem<4><3> ), .D(n2513), .Y(
        n1610) );
  AOI22X1 U2104 ( .A(\mem<3><3> ), .B(n2509), .C(\mem<2><3> ), .D(n2581), .Y(
        n1608) );
  AOI22X1 U2105 ( .A(\mem<1><3> ), .B(n2455), .C(n1403), .D(\mem<0><3> ), .Y(
        n1607) );
  AOI22X1 U2107 ( .A(\mem<15><3> ), .B(n2505), .C(\mem<14><3> ), .D(n2507), 
        .Y(n1616) );
  AOI22X1 U2108 ( .A(\mem<13><3> ), .B(n2501), .C(\mem<12><3> ), .D(n2503), 
        .Y(n1615) );
  AOI22X1 U2109 ( .A(\mem<11><3> ), .B(n2497), .C(\mem<10><3> ), .D(n2499), 
        .Y(n1613) );
  AOI22X1 U2110 ( .A(\mem<9><3> ), .B(n2493), .C(\mem<8><3> ), .D(n2495), .Y(
        n1612) );
  AOI22X1 U2112 ( .A(\mem<23><3> ), .B(n2489), .C(\mem<22><3> ), .D(n2491), 
        .Y(n1623) );
  AOI22X1 U2113 ( .A(\mem<21><3> ), .B(n2485), .C(\mem<20><3> ), .D(n2487), 
        .Y(n1622) );
  AOI22X1 U2114 ( .A(\mem<19><3> ), .B(n2481), .C(\mem<18><3> ), .D(n2483), 
        .Y(n1620) );
  AOI22X1 U2115 ( .A(\mem<17><3> ), .B(n2477), .C(\mem<16><3> ), .D(n2479), 
        .Y(n1619) );
  AOI22X1 U2117 ( .A(\mem<31><3> ), .B(n2473), .C(\mem<30><3> ), .D(n2475), 
        .Y(n1628) );
  AOI22X1 U2118 ( .A(\mem<29><3> ), .B(n2469), .C(\mem<28><3> ), .D(n2471), 
        .Y(n1627) );
  AOI22X1 U2119 ( .A(\mem<27><3> ), .B(n2465), .C(\mem<26><3> ), .D(n2467), 
        .Y(n1625) );
  AOI22X1 U2120 ( .A(\mem<25><3> ), .B(n2461), .C(\mem<24><3> ), .D(n2463), 
        .Y(n1624) );
  AOI21X1 U2121 ( .A(n1629), .B(n1630), .C(n2451), .Y(n3714) );
  NOR3X1 U2122 ( .A(n1631), .B(n170), .C(n183), .Y(n1630) );
  AOI22X1 U2124 ( .A(\mem<55><2> ), .B(n2577), .C(\mem<54><2> ), .D(n2579), 
        .Y(n1638) );
  AOI22X1 U2125 ( .A(\mem<53><2> ), .B(n2573), .C(\mem<52><2> ), .D(n2575), 
        .Y(n1637) );
  AOI22X1 U2126 ( .A(\mem<51><2> ), .B(n2569), .C(\mem<50><2> ), .D(n2571), 
        .Y(n1635) );
  AOI22X1 U2127 ( .A(\mem<49><2> ), .B(n2565), .C(\mem<48><2> ), .D(n2567), 
        .Y(n1634) );
  AOI22X1 U2129 ( .A(\mem<63><2> ), .B(n2459), .C(\mem<62><2> ), .D(n2563), 
        .Y(n1643) );
  AOI22X1 U2130 ( .A(\mem<61><2> ), .B(n2559), .C(\mem<60><2> ), .D(n2561), 
        .Y(n1642) );
  AOI22X1 U2131 ( .A(\mem<59><2> ), .B(n2555), .C(\mem<58><2> ), .D(n2557), 
        .Y(n1640) );
  AOI22X1 U2132 ( .A(\mem<57><2> ), .B(n2551), .C(\mem<56><2> ), .D(n2553), 
        .Y(n1639) );
  AOI22X1 U2134 ( .A(\mem<39><2> ), .B(n2547), .C(\mem<38><2> ), .D(n2549), 
        .Y(n1650) );
  AOI22X1 U2135 ( .A(\mem<37><2> ), .B(n2543), .C(\mem<36><2> ), .D(n2545), 
        .Y(n1649) );
  AOI22X1 U2136 ( .A(\mem<35><2> ), .B(n2539), .C(\mem<34><2> ), .D(n2541), 
        .Y(n1647) );
  AOI22X1 U2137 ( .A(\mem<33><2> ), .B(n2536), .C(\mem<32><2> ), .D(n2537), 
        .Y(n1646) );
  AOI22X1 U2139 ( .A(\mem<47><2> ), .B(n2531), .C(\mem<46><2> ), .D(n2533), 
        .Y(n1655) );
  AOI22X1 U2140 ( .A(\mem<45><2> ), .B(n2527), .C(\mem<44><2> ), .D(n2529), 
        .Y(n1654) );
  AOI22X1 U2141 ( .A(\mem<43><2> ), .B(n2523), .C(\mem<42><2> ), .D(n2525), 
        .Y(n1652) );
  AOI22X1 U2142 ( .A(\mem<41><2> ), .B(n2519), .C(\mem<40><2> ), .D(n2521), 
        .Y(n1651) );
  NOR3X1 U2143 ( .A(n1656), .B(n169), .C(n214), .Y(n1629) );
  AOI22X1 U2145 ( .A(\mem<7><2> ), .B(n2515), .C(\mem<6><2> ), .D(n2517), .Y(
        n1663) );
  AOI22X1 U2146 ( .A(\mem<5><2> ), .B(n2511), .C(\mem<4><2> ), .D(n2513), .Y(
        n1662) );
  AOI22X1 U2147 ( .A(\mem<3><2> ), .B(n2509), .C(\mem<2><2> ), .D(n2581), .Y(
        n1660) );
  AOI22X1 U2148 ( .A(\mem<1><2> ), .B(n2455), .C(n1403), .D(\mem<0><2> ), .Y(
        n1659) );
  AOI22X1 U2150 ( .A(\mem<15><2> ), .B(n2505), .C(\mem<14><2> ), .D(n2507), 
        .Y(n1668) );
  AOI22X1 U2151 ( .A(\mem<13><2> ), .B(n2501), .C(\mem<12><2> ), .D(n2503), 
        .Y(n1667) );
  AOI22X1 U2152 ( .A(\mem<11><2> ), .B(n2497), .C(\mem<10><2> ), .D(n2499), 
        .Y(n1665) );
  AOI22X1 U2153 ( .A(\mem<9><2> ), .B(n2493), .C(\mem<8><2> ), .D(n2495), .Y(
        n1664) );
  AOI22X1 U2155 ( .A(\mem<23><2> ), .B(n2489), .C(\mem<22><2> ), .D(n2491), 
        .Y(n1675) );
  AOI22X1 U2156 ( .A(\mem<21><2> ), .B(n2485), .C(\mem<20><2> ), .D(n2487), 
        .Y(n1674) );
  AOI22X1 U2157 ( .A(\mem<19><2> ), .B(n2481), .C(\mem<18><2> ), .D(n2483), 
        .Y(n1672) );
  AOI22X1 U2158 ( .A(\mem<17><2> ), .B(n2477), .C(\mem<16><2> ), .D(n2479), 
        .Y(n1671) );
  AOI22X1 U2160 ( .A(\mem<31><2> ), .B(n2473), .C(\mem<30><2> ), .D(n2475), 
        .Y(n1680) );
  AOI22X1 U2161 ( .A(\mem<29><2> ), .B(n2469), .C(\mem<28><2> ), .D(n2471), 
        .Y(n1679) );
  AOI22X1 U2162 ( .A(\mem<27><2> ), .B(n2465), .C(\mem<26><2> ), .D(n2467), 
        .Y(n1677) );
  AOI22X1 U2163 ( .A(\mem<25><2> ), .B(n2461), .C(\mem<24><2> ), .D(n2463), 
        .Y(n1676) );
  AOI21X1 U2164 ( .A(n1681), .B(n1682), .C(n2451), .Y(n3715) );
  NOR3X1 U2165 ( .A(n1683), .B(n168), .C(n182), .Y(n1682) );
  AOI22X1 U2167 ( .A(\mem<55><1> ), .B(n2577), .C(\mem<54><1> ), .D(n2579), 
        .Y(n1690) );
  AOI22X1 U2168 ( .A(\mem<53><1> ), .B(n2573), .C(\mem<52><1> ), .D(n2575), 
        .Y(n1689) );
  AOI22X1 U2169 ( .A(\mem<51><1> ), .B(n2569), .C(\mem<50><1> ), .D(n2571), 
        .Y(n1687) );
  AOI22X1 U2170 ( .A(\mem<49><1> ), .B(n2565), .C(\mem<48><1> ), .D(n2567), 
        .Y(n1686) );
  AOI22X1 U2172 ( .A(\mem<63><1> ), .B(n2459), .C(\mem<62><1> ), .D(n2563), 
        .Y(n1695) );
  AOI22X1 U2173 ( .A(\mem<61><1> ), .B(n2559), .C(\mem<60><1> ), .D(n2561), 
        .Y(n1694) );
  AOI22X1 U2174 ( .A(\mem<59><1> ), .B(n2555), .C(\mem<58><1> ), .D(n2557), 
        .Y(n1692) );
  AOI22X1 U2175 ( .A(\mem<57><1> ), .B(n2551), .C(\mem<56><1> ), .D(n2553), 
        .Y(n1691) );
  AOI22X1 U2177 ( .A(\mem<39><1> ), .B(n2547), .C(\mem<38><1> ), .D(n2549), 
        .Y(n1702) );
  AOI22X1 U2178 ( .A(\mem<37><1> ), .B(n2543), .C(\mem<36><1> ), .D(n2545), 
        .Y(n1701) );
  AOI22X1 U2179 ( .A(\mem<35><1> ), .B(n2539), .C(\mem<34><1> ), .D(n2541), 
        .Y(n1699) );
  AOI22X1 U2180 ( .A(\mem<33><1> ), .B(n2536), .C(\mem<32><1> ), .D(n2537), 
        .Y(n1698) );
  AOI22X1 U2182 ( .A(\mem<47><1> ), .B(n2531), .C(\mem<46><1> ), .D(n2533), 
        .Y(n1707) );
  AOI22X1 U2183 ( .A(\mem<45><1> ), .B(n2527), .C(\mem<44><1> ), .D(n2529), 
        .Y(n1706) );
  AOI22X1 U2184 ( .A(\mem<43><1> ), .B(n2523), .C(\mem<42><1> ), .D(n2525), 
        .Y(n1704) );
  AOI22X1 U2185 ( .A(\mem<41><1> ), .B(n2519), .C(\mem<40><1> ), .D(n2521), 
        .Y(n1703) );
  NOR3X1 U2186 ( .A(n1708), .B(n167), .C(n211), .Y(n1681) );
  AOI22X1 U2188 ( .A(\mem<7><1> ), .B(n2515), .C(\mem<6><1> ), .D(n2517), .Y(
        n1715) );
  AOI22X1 U2189 ( .A(\mem<5><1> ), .B(n2511), .C(\mem<4><1> ), .D(n2513), .Y(
        n1714) );
  AOI22X1 U2190 ( .A(\mem<3><1> ), .B(n2509), .C(\mem<2><1> ), .D(n2581), .Y(
        n1712) );
  AOI22X1 U2191 ( .A(\mem<1><1> ), .B(n2455), .C(n1403), .D(\mem<0><1> ), .Y(
        n1711) );
  AOI22X1 U2193 ( .A(\mem<15><1> ), .B(n2505), .C(\mem<14><1> ), .D(n2507), 
        .Y(n1720) );
  AOI22X1 U2194 ( .A(\mem<13><1> ), .B(n2501), .C(\mem<12><1> ), .D(n2503), 
        .Y(n1719) );
  AOI22X1 U2195 ( .A(\mem<11><1> ), .B(n2497), .C(\mem<10><1> ), .D(n2499), 
        .Y(n1717) );
  AOI22X1 U2196 ( .A(\mem<9><1> ), .B(n2493), .C(\mem<8><1> ), .D(n2495), .Y(
        n1716) );
  AOI22X1 U2198 ( .A(\mem<23><1> ), .B(n2489), .C(\mem<22><1> ), .D(n2491), 
        .Y(n1727) );
  AOI22X1 U2199 ( .A(\mem<21><1> ), .B(n2485), .C(\mem<20><1> ), .D(n2487), 
        .Y(n1726) );
  AOI22X1 U2200 ( .A(\mem<19><1> ), .B(n2481), .C(\mem<18><1> ), .D(n2483), 
        .Y(n1724) );
  AOI22X1 U2201 ( .A(\mem<17><1> ), .B(n2477), .C(\mem<16><1> ), .D(n2479), 
        .Y(n1723) );
  AOI22X1 U2203 ( .A(\mem<31><1> ), .B(n2473), .C(\mem<30><1> ), .D(n2475), 
        .Y(n1732) );
  AOI22X1 U2204 ( .A(\mem<29><1> ), .B(n2469), .C(\mem<28><1> ), .D(n2471), 
        .Y(n1731) );
  AOI22X1 U2205 ( .A(\mem<27><1> ), .B(n2465), .C(\mem<26><1> ), .D(n2467), 
        .Y(n1729) );
  AOI22X1 U2206 ( .A(\mem<25><1> ), .B(n2461), .C(\mem<24><1> ), .D(n2463), 
        .Y(n1728) );
  AOI21X1 U2207 ( .A(n1733), .B(n1734), .C(n2451), .Y(n3716) );
  NOR3X1 U2209 ( .A(n1735), .B(n166), .C(n181), .Y(n1734) );
  AOI22X1 U2211 ( .A(\mem<55><0> ), .B(n2577), .C(\mem<54><0> ), .D(n2579), 
        .Y(n1742) );
  AOI22X1 U2214 ( .A(\mem<53><0> ), .B(n2573), .C(\mem<52><0> ), .D(n2575), 
        .Y(n1741) );
  AOI22X1 U2217 ( .A(\mem<51><0> ), .B(n2569), .C(\mem<50><0> ), .D(n2571), 
        .Y(n1739) );
  AOI22X1 U2220 ( .A(\mem<49><0> ), .B(n2565), .C(\mem<48><0> ), .D(n2567), 
        .Y(n1738) );
  AOI22X1 U2224 ( .A(\mem<63><0> ), .B(n2459), .C(\mem<62><0> ), .D(n2563), 
        .Y(n1754) );
  AOI22X1 U2227 ( .A(\mem<61><0> ), .B(n2559), .C(\mem<60><0> ), .D(n2561), 
        .Y(n1753) );
  AOI22X1 U2230 ( .A(\mem<59><0> ), .B(n2555), .C(\mem<58><0> ), .D(n2557), 
        .Y(n1751) );
  AOI22X1 U2233 ( .A(\mem<57><0> ), .B(n2551), .C(\mem<56><0> ), .D(n2553), 
        .Y(n1750) );
  NAND3X1 U2235 ( .A(n1756), .B(N182), .C(n1757), .Y(n1755) );
  AOI22X1 U2239 ( .A(\mem<39><0> ), .B(n2547), .C(\mem<38><0> ), .D(n2549), 
        .Y(n1764) );
  AOI22X1 U2242 ( .A(\mem<37><0> ), .B(n2543), .C(\mem<36><0> ), .D(n2545), 
        .Y(n1763) );
  AOI22X1 U2245 ( .A(\mem<35><0> ), .B(n2539), .C(\mem<34><0> ), .D(n2541), 
        .Y(n1761) );
  AOI22X1 U2248 ( .A(\mem<33><0> ), .B(n2536), .C(\mem<32><0> ), .D(n2537), 
        .Y(n1760) );
  AOI22X1 U2252 ( .A(\mem<47><0> ), .B(n2531), .C(\mem<46><0> ), .D(n2533), 
        .Y(n1769) );
  AOI22X1 U2255 ( .A(\mem<45><0> ), .B(n2527), .C(\mem<44><0> ), .D(n2529), 
        .Y(n1768) );
  AOI22X1 U2258 ( .A(\mem<43><0> ), .B(n2523), .C(\mem<42><0> ), .D(n2525), 
        .Y(n1766) );
  AOI22X1 U2261 ( .A(\mem<41><0> ), .B(n2519), .C(\mem<40><0> ), .D(n2521), 
        .Y(n1765) );
  NAND3X1 U2263 ( .A(n1756), .B(N182), .C(n2353), .Y(n1770) );
  NAND3X1 U2266 ( .A(n1756), .B(N182), .C(n2351), .Y(n1772) );
  NOR3X1 U2268 ( .A(n1774), .B(n165), .C(n208), .Y(n1733) );
  AOI22X1 U2270 ( .A(\mem<7><0> ), .B(n2515), .C(\mem<6><0> ), .D(n2517), .Y(
        n1781) );
  AOI22X1 U2273 ( .A(\mem<5><0> ), .B(n2511), .C(\mem<4><0> ), .D(n2513), .Y(
        n1780) );
  AOI22X1 U2276 ( .A(\mem<3><0> ), .B(n2509), .C(\mem<2><0> ), .D(n2581), .Y(
        n1778) );
  AOI22X1 U2279 ( .A(\mem<1><0> ), .B(n2455), .C(n1403), .D(\mem<0><0> ), .Y(
        n1777) );
  NOR3X1 U2280 ( .A(n1782), .B(n1783), .C(n1784), .Y(n1403) );
  NAND3X1 U2281 ( .A(\addr<8> ), .B(\addr<7> ), .C(\addr<9> ), .Y(n1786) );
  NAND3X1 U2282 ( .A(\addr<15> ), .B(\addr<14> ), .C(\addr<6> ), .Y(n1785) );
  NAND3X1 U2283 ( .A(\addr<10> ), .B(n3192), .C(n3187), .Y(n1783) );
  NAND3X1 U2284 ( .A(N181), .B(N180), .C(N182), .Y(n1787) );
  NAND3X1 U2285 ( .A(\addr<13> ), .B(\addr<11> ), .C(\addr<12> ), .Y(n1782) );
  AOI22X1 U2288 ( .A(\mem<15><0> ), .B(n2505), .C(\mem<14><0> ), .D(n2507), 
        .Y(n1792) );
  AOI22X1 U2291 ( .A(\mem<13><0> ), .B(n2501), .C(\mem<12><0> ), .D(n2503), 
        .Y(n1791) );
  AOI22X1 U2294 ( .A(\mem<11><0> ), .B(n2497), .C(\mem<10><0> ), .D(n2499), 
        .Y(n1789) );
  AOI22X1 U2297 ( .A(\mem<9><0> ), .B(n2493), .C(\mem<8><0> ), .D(n2495), .Y(
        n1788) );
  AOI22X1 U2302 ( .A(\mem<23><0> ), .B(n2489), .C(\mem<22><0> ), .D(n2491), 
        .Y(n1801) );
  AOI22X1 U2305 ( .A(\mem<21><0> ), .B(n2485), .C(\mem<20><0> ), .D(n2487), 
        .Y(n1800) );
  AOI22X1 U2308 ( .A(\mem<19><0> ), .B(n2481), .C(\mem<18><0> ), .D(n2483), 
        .Y(n1798) );
  AOI22X1 U2311 ( .A(\mem<17><0> ), .B(n2477), .C(\mem<16><0> ), .D(n2479), 
        .Y(n1797) );
  AOI22X1 U2317 ( .A(\mem<31><0> ), .B(n2473), .C(\mem<30><0> ), .D(n2475), 
        .Y(n1807) );
  NOR3X1 U2319 ( .A(n3184), .B(n3182), .C(n3181), .Y(n1743) );
  NOR3X1 U2321 ( .A(n3183), .B(N177), .C(n3184), .Y(n1744) );
  AOI22X1 U2322 ( .A(\mem<29><0> ), .B(n2469), .C(\mem<28><0> ), .D(n2471), 
        .Y(n1806) );
  NOR3X1 U2324 ( .A(n3183), .B(N179), .C(n3181), .Y(n1745) );
  NOR3X1 U2326 ( .A(N177), .B(n3182), .C(n3184), .Y(n1746) );
  AOI22X1 U2327 ( .A(\mem<27><0> ), .B(n2465), .C(\mem<26><0> ), .D(n2467), 
        .Y(n1804) );
  NOR3X1 U2329 ( .A(n3182), .B(N179), .C(n3181), .Y(n1747) );
  NOR3X1 U2331 ( .A(N177), .B(N179), .C(n3183), .Y(n1748) );
  AOI22X1 U2332 ( .A(\mem<25><0> ), .B(n2461), .C(\mem<24><0> ), .D(n2463), 
        .Y(n1803) );
  NAND3X1 U2334 ( .A(N179), .B(n3182), .C(N177), .Y(n612) );
  NAND3X1 U2335 ( .A(n1756), .B(N181), .C(n1809), .Y(n1808) );
  NOR2X1 U2336 ( .A(N182), .B(N180), .Y(n1809) );
  NOR3X1 U2338 ( .A(n3182), .B(N179), .C(N177), .Y(n1749) );
  NAND3X1 U2339 ( .A(n1811), .B(N181), .C(n1756), .Y(n1810) );
  NOR2X1 U2340 ( .A(N182), .B(n3185), .Y(n1811) );
  NOR3X1 U2341 ( .A(n3194), .B(\addr<6> ), .C(\addr<15> ), .Y(n1813) );
  NOR3X1 U2342 ( .A(\addr<8> ), .B(\addr<9> ), .C(\addr<7> ), .Y(n1814) );
  NOR3X1 U2343 ( .A(n3195), .B(\addr<11> ), .C(\addr<10> ), .Y(n1812) );
  NOR3X1 U2344 ( .A(\addr<13> ), .B(\addr<14> ), .C(\addr<12> ), .Y(n1815) );
  INVX1 U3 ( .A(n2452), .Y(n3178) );
  AND2X1 U4 ( .A(n1812), .B(n1813), .Y(n1756) );
  INVX1 U5 ( .A(n1815), .Y(n3195) );
  BUFX2 U6 ( .A(n1346), .Y(n3113) );
  OR2X1 U7 ( .A(n8), .B(n9), .Y(n7) );
  OR2X1 U8 ( .A(n18), .B(n19), .Y(n17) );
  OR2X1 U9 ( .A(n28), .B(n29), .Y(n27) );
  OR2X1 U10 ( .A(n38), .B(n39), .Y(n37) );
  OR2X1 U11 ( .A(n48), .B(n49), .Y(n47) );
  OR2X1 U12 ( .A(n58), .B(n59), .Y(n57) );
  OR2X1 U13 ( .A(n68), .B(n69), .Y(n67) );
  OR2X1 U14 ( .A(n78), .B(n79), .Y(n77) );
  OR2X1 U15 ( .A(n88), .B(n89), .Y(n87) );
  OR2X1 U16 ( .A(n98), .B(n99), .Y(n97) );
  OR2X1 U17 ( .A(n108), .B(n109), .Y(n107) );
  OR2X1 U18 ( .A(n118), .B(n119), .Y(n117) );
  OR2X1 U19 ( .A(n128), .B(n129), .Y(n127) );
  OR2X1 U20 ( .A(n138), .B(n139), .Y(n137) );
  OR2X1 U21 ( .A(n148), .B(n149), .Y(n147) );
  OR2X1 U22 ( .A(n158), .B(n159), .Y(n157) );
  AND2X1 U23 ( .A(N189), .B(n2450), .Y(\data_out<11> ) );
  AND2X1 U24 ( .A(n3178), .B(n610), .Y(n598) );
  AND2X1 U25 ( .A(n598), .B(n2460), .Y(n600) );
  AND2X1 U26 ( .A(n2459), .B(n598), .Y(n601) );
  AND2X1 U27 ( .A(n3174), .B(n2564), .Y(n615) );
  AND2X1 U28 ( .A(n2563), .B(n3174), .Y(n616) );
  AND2X1 U29 ( .A(n3173), .B(n2560), .Y(n628) );
  AND2X1 U30 ( .A(n2559), .B(n3173), .Y(n629) );
  AND2X1 U31 ( .A(n3172), .B(n2562), .Y(n640) );
  AND2X1 U32 ( .A(n2561), .B(n3172), .Y(n641) );
  AND2X1 U33 ( .A(n3171), .B(n2556), .Y(n652) );
  AND2X1 U34 ( .A(n2555), .B(n3171), .Y(n653) );
  AND2X1 U35 ( .A(n3170), .B(n2558), .Y(n664) );
  AND2X1 U36 ( .A(n2557), .B(n3170), .Y(n665) );
  AND2X1 U37 ( .A(n3169), .B(n2552), .Y(n676) );
  AND2X1 U38 ( .A(n2551), .B(n3169), .Y(n677) );
  AND2X1 U39 ( .A(n3168), .B(n2554), .Y(n688) );
  AND2X1 U40 ( .A(n2553), .B(n3168), .Y(n689) );
  AND2X1 U41 ( .A(n3167), .B(n2578), .Y(n700) );
  AND2X1 U42 ( .A(n2577), .B(n3167), .Y(n701) );
  AND2X1 U43 ( .A(n3166), .B(n2580), .Y(n712) );
  AND2X1 U44 ( .A(n2579), .B(n3166), .Y(n713) );
  AND2X1 U45 ( .A(n3165), .B(n2574), .Y(n724) );
  AND2X1 U46 ( .A(n2573), .B(n3165), .Y(n725) );
  AND2X1 U47 ( .A(n3164), .B(n2576), .Y(n736) );
  AND2X1 U48 ( .A(n2575), .B(n3164), .Y(n737) );
  AND2X1 U49 ( .A(n3163), .B(n2570), .Y(n748) );
  AND2X1 U50 ( .A(n2569), .B(n3163), .Y(n749) );
  AND2X1 U51 ( .A(n3162), .B(n2572), .Y(n760) );
  AND2X1 U52 ( .A(n2571), .B(n3162), .Y(n761) );
  AND2X1 U53 ( .A(n3161), .B(n2566), .Y(n772) );
  AND2X1 U54 ( .A(n2565), .B(n3161), .Y(n773) );
  AND2X1 U55 ( .A(n3160), .B(n2568), .Y(n784) );
  AND2X1 U56 ( .A(n2567), .B(n3160), .Y(n785) );
  AND2X1 U57 ( .A(n3159), .B(n2532), .Y(n796) );
  AND2X1 U58 ( .A(n2531), .B(n3159), .Y(n797) );
  AND2X1 U59 ( .A(n3158), .B(n2534), .Y(n808) );
  AND2X1 U60 ( .A(n2533), .B(n3158), .Y(n809) );
  AND2X1 U61 ( .A(n3157), .B(n2528), .Y(n820) );
  AND2X1 U62 ( .A(n2527), .B(n3157), .Y(n821) );
  AND2X1 U63 ( .A(n3156), .B(n2530), .Y(n832) );
  AND2X1 U64 ( .A(n2529), .B(n3156), .Y(n833) );
  AND2X1 U65 ( .A(n3155), .B(n2524), .Y(n844) );
  AND2X1 U66 ( .A(n2523), .B(n3155), .Y(n845) );
  AND2X1 U67 ( .A(n3154), .B(n2526), .Y(n856) );
  AND2X1 U68 ( .A(n2525), .B(n3154), .Y(n857) );
  AND2X1 U69 ( .A(n3153), .B(n2520), .Y(n868) );
  AND2X1 U70 ( .A(n2519), .B(n3153), .Y(n869) );
  AND2X1 U71 ( .A(n3152), .B(n2522), .Y(n880) );
  AND2X1 U72 ( .A(n2521), .B(n3152), .Y(n881) );
  AND2X1 U73 ( .A(n3151), .B(n2548), .Y(n892) );
  AND2X1 U74 ( .A(n2547), .B(n3151), .Y(n893) );
  AND2X1 U75 ( .A(n3150), .B(n2550), .Y(n904) );
  AND2X1 U76 ( .A(n2549), .B(n3150), .Y(n905) );
  AND2X1 U77 ( .A(n3149), .B(n2544), .Y(n916) );
  AND2X1 U78 ( .A(n2543), .B(n3149), .Y(n917) );
  AND2X1 U79 ( .A(n3148), .B(n2546), .Y(n928) );
  AND2X1 U80 ( .A(n2545), .B(n3148), .Y(n929) );
  AND2X1 U81 ( .A(n3147), .B(n2540), .Y(n940) );
  AND2X1 U82 ( .A(n2539), .B(n3147), .Y(n941) );
  AND2X1 U83 ( .A(n3146), .B(n2542), .Y(n952) );
  AND2X1 U84 ( .A(n2541), .B(n3146), .Y(n953) );
  AND2X1 U85 ( .A(n3145), .B(n2535), .Y(n964) );
  AND2X1 U86 ( .A(n2536), .B(n3145), .Y(n965) );
  AND2X1 U87 ( .A(n3144), .B(n2538), .Y(n976) );
  AND2X1 U88 ( .A(n2537), .B(n3144), .Y(n977) );
  AND2X1 U89 ( .A(n3143), .B(n2474), .Y(n988) );
  AND2X1 U90 ( .A(n2473), .B(n3143), .Y(n989) );
  AND2X1 U91 ( .A(n3142), .B(n2476), .Y(n1000) );
  AND2X1 U92 ( .A(n2475), .B(n3142), .Y(n1001) );
  AND2X1 U93 ( .A(n3141), .B(n2470), .Y(n1012) );
  AND2X1 U94 ( .A(n2469), .B(n3141), .Y(n1013) );
  AND2X1 U95 ( .A(n3140), .B(n2472), .Y(n1024) );
  AND2X1 U96 ( .A(n2471), .B(n3140), .Y(n1025) );
  AND2X1 U97 ( .A(n3139), .B(n2466), .Y(n1036) );
  AND2X1 U98 ( .A(n2465), .B(n3139), .Y(n1037) );
  AND2X1 U99 ( .A(n3138), .B(n2468), .Y(n1048) );
  AND2X1 U100 ( .A(n2467), .B(n3138), .Y(n1049) );
  AND2X1 U101 ( .A(n3137), .B(n2462), .Y(n1060) );
  AND2X1 U102 ( .A(n2461), .B(n3137), .Y(n1061) );
  AND2X1 U103 ( .A(n3136), .B(n2464), .Y(n1072) );
  AND2X1 U104 ( .A(n2463), .B(n3136), .Y(n1073) );
  AND2X1 U105 ( .A(n3135), .B(n2490), .Y(n1084) );
  AND2X1 U106 ( .A(n2489), .B(n3135), .Y(n1085) );
  AND2X1 U107 ( .A(n3134), .B(n2492), .Y(n1096) );
  AND2X1 U108 ( .A(n2491), .B(n3134), .Y(n1097) );
  AND2X1 U109 ( .A(n3133), .B(n2486), .Y(n1108) );
  AND2X1 U110 ( .A(n2485), .B(n3133), .Y(n1109) );
  AND2X1 U111 ( .A(n3132), .B(n2488), .Y(n1120) );
  AND2X1 U112 ( .A(n2487), .B(n3132), .Y(n1121) );
  AND2X1 U113 ( .A(n3131), .B(n2482), .Y(n1132) );
  AND2X1 U114 ( .A(n2481), .B(n3131), .Y(n1133) );
  AND2X1 U115 ( .A(n3130), .B(n2484), .Y(n1144) );
  AND2X1 U116 ( .A(n2483), .B(n3130), .Y(n1145) );
  AND2X1 U117 ( .A(n3129), .B(n2478), .Y(n1156) );
  AND2X1 U118 ( .A(n2477), .B(n3129), .Y(n1157) );
  AND2X1 U119 ( .A(n3128), .B(n2480), .Y(n1168) );
  AND2X1 U120 ( .A(n2479), .B(n3128), .Y(n1169) );
  AND2X1 U121 ( .A(n3127), .B(n2506), .Y(n1180) );
  AND2X1 U122 ( .A(n2505), .B(n3127), .Y(n1181) );
  AND2X1 U123 ( .A(n3126), .B(n2508), .Y(n1192) );
  AND2X1 U124 ( .A(n2507), .B(n3126), .Y(n1193) );
  AND2X1 U125 ( .A(n3125), .B(n2502), .Y(n1204) );
  AND2X1 U126 ( .A(n2501), .B(n3125), .Y(n1205) );
  AND2X1 U127 ( .A(n3124), .B(n2504), .Y(n1216) );
  AND2X1 U128 ( .A(n2503), .B(n3124), .Y(n1217) );
  AND2X1 U129 ( .A(n3123), .B(n2498), .Y(n1228) );
  AND2X1 U130 ( .A(n2497), .B(n3123), .Y(n1229) );
  AND2X1 U131 ( .A(n3122), .B(n2500), .Y(n1240) );
  AND2X1 U134 ( .A(n2499), .B(n3122), .Y(n1241) );
  AND2X1 U139 ( .A(n3121), .B(n2494), .Y(n1252) );
  AND2X1 U144 ( .A(n2493), .B(n3121), .Y(n1253) );
  AND2X1 U149 ( .A(n3120), .B(n2496), .Y(n1264) );
  AND2X1 U154 ( .A(n2495), .B(n3120), .Y(n1265) );
  AND2X1 U159 ( .A(n3119), .B(n2516), .Y(n1276) );
  AND2X1 U164 ( .A(n2515), .B(n3119), .Y(n1277) );
  AND2X1 U169 ( .A(n3118), .B(n2518), .Y(n1288) );
  AND2X1 U174 ( .A(n2517), .B(n3118), .Y(n1289) );
  AND2X1 U179 ( .A(n3117), .B(n2512), .Y(n1300) );
  AND2X1 U184 ( .A(n2511), .B(n3117), .Y(n1301) );
  AND2X1 U189 ( .A(n3116), .B(n2514), .Y(n1312) );
  AND2X1 U194 ( .A(n2513), .B(n3116), .Y(n1313) );
  AND2X1 U199 ( .A(n3115), .B(n2510), .Y(n1324) );
  AND2X1 U202 ( .A(n2509), .B(n3115), .Y(n1325) );
  AND2X1 U203 ( .A(n3114), .B(n2582), .Y(n1336) );
  AND2X1 U204 ( .A(n2581), .B(n3114), .Y(n1337) );
  AND2X1 U205 ( .A(n3113), .B(n2456), .Y(n1348) );
  AND2X1 U206 ( .A(n2455), .B(n3113), .Y(n1349) );
  INVX1 U207 ( .A(n3093), .Y(n3101) );
  INVX1 U210 ( .A(n3093), .Y(n3102) );
  INVX1 U211 ( .A(n3092), .Y(n3103) );
  INVX1 U217 ( .A(n3092), .Y(n3104) );
  INVX1 U220 ( .A(n3092), .Y(n3105) );
  INVX1 U221 ( .A(n3091), .Y(n3106) );
  INVX1 U222 ( .A(n3091), .Y(n3107) );
  INVX1 U223 ( .A(n3091), .Y(n3108) );
  INVX1 U224 ( .A(n3090), .Y(n3109) );
  INVX1 U225 ( .A(n3090), .Y(n3111) );
  INVX1 U226 ( .A(n3090), .Y(n3110) );
  INVX1 U227 ( .A(n1814), .Y(n3194) );
  AND2X1 U228 ( .A(n3185), .B(N181), .Y(n1757) );
  OR2X1 U229 ( .A(n2341), .B(n190), .Y(n161) );
  OR2X1 U230 ( .A(n2341), .B(n191), .Y(n163) );
  OR2X1 U231 ( .A(n1), .B(n6), .Y(n1774) );
  OR2X1 U232 ( .A(n11), .B(n16), .Y(n1735) );
  OR2X1 U233 ( .A(n21), .B(n26), .Y(n1708) );
  OR2X1 U234 ( .A(n31), .B(n36), .Y(n1683) );
  OR2X1 U235 ( .A(n41), .B(n46), .Y(n1656) );
  OR2X1 U236 ( .A(n51), .B(n56), .Y(n1631) );
  OR2X1 U237 ( .A(n61), .B(n66), .Y(n1604) );
  OR2X1 U238 ( .A(n71), .B(n76), .Y(n1579) );
  OR2X1 U239 ( .A(n81), .B(n86), .Y(n1552) );
  OR2X1 U240 ( .A(n91), .B(n96), .Y(n1527) );
  OR2X1 U241 ( .A(n101), .B(n106), .Y(n1500) );
  OR2X1 U242 ( .A(n111), .B(n116), .Y(n1475) );
  OR2X1 U243 ( .A(n121), .B(n126), .Y(n1448) );
  OR2X1 U244 ( .A(n131), .B(n136), .Y(n1423) );
  OR2X1 U245 ( .A(n141), .B(n146), .Y(n1395) );
  OR2X1 U246 ( .A(n151), .B(n156), .Y(n1370) );
  INVX1 U247 ( .A(wr), .Y(n3708) );
  INVX1 U248 ( .A(n2452), .Y(n3180) );
  INVX2 U249 ( .A(n2452), .Y(n3179) );
  AND2X1 U250 ( .A(N192), .B(n2450), .Y(\data_out<8> ) );
  AND2X1 U251 ( .A(N191), .B(n2450), .Y(\data_out<9> ) );
  AND2X1 U252 ( .A(N190), .B(n2450), .Y(\data_out<10> ) );
  AND2X1 U253 ( .A(N188), .B(n2450), .Y(\data_out<12> ) );
  AND2X1 U254 ( .A(N187), .B(n2450), .Y(\data_out<13> ) );
  AND2X1 U255 ( .A(N186), .B(n2450), .Y(\data_out<14> ) );
  AND2X1 U256 ( .A(N185), .B(n2450), .Y(\data_out<15> ) );
  INVX1 U257 ( .A(\mem<63><0> ), .Y(n3707) );
  INVX1 U258 ( .A(\mem<63><1> ), .Y(n3706) );
  INVX1 U259 ( .A(\mem<63><2> ), .Y(n3705) );
  INVX1 U260 ( .A(\mem<63><3> ), .Y(n3704) );
  INVX1 U261 ( .A(\mem<63><4> ), .Y(n3703) );
  INVX1 U262 ( .A(\mem<63><5> ), .Y(n3702) );
  INVX1 U263 ( .A(\mem<63><6> ), .Y(n3701) );
  INVX1 U264 ( .A(\mem<63><7> ), .Y(n3700) );
  INVX1 U265 ( .A(\mem<62><0> ), .Y(n3699) );
  INVX1 U266 ( .A(\mem<62><1> ), .Y(n3698) );
  INVX1 U267 ( .A(\mem<62><2> ), .Y(n3697) );
  INVX1 U268 ( .A(\mem<62><3> ), .Y(n3696) );
  INVX1 U269 ( .A(\mem<62><4> ), .Y(n3695) );
  INVX1 U270 ( .A(\mem<62><5> ), .Y(n3694) );
  INVX1 U271 ( .A(\mem<62><6> ), .Y(n3693) );
  INVX1 U272 ( .A(\mem<62><7> ), .Y(n3692) );
  INVX1 U273 ( .A(\mem<61><0> ), .Y(n3691) );
  INVX1 U274 ( .A(\mem<61><1> ), .Y(n3690) );
  INVX1 U275 ( .A(\mem<61><2> ), .Y(n3689) );
  INVX1 U276 ( .A(\mem<61><3> ), .Y(n3688) );
  INVX1 U277 ( .A(\mem<61><4> ), .Y(n3687) );
  INVX1 U278 ( .A(\mem<61><5> ), .Y(n3686) );
  INVX1 U279 ( .A(\mem<61><6> ), .Y(n3685) );
  INVX1 U280 ( .A(\mem<61><7> ), .Y(n3684) );
  INVX1 U281 ( .A(\mem<60><0> ), .Y(n3683) );
  INVX1 U282 ( .A(\mem<60><1> ), .Y(n3682) );
  INVX1 U283 ( .A(\mem<60><2> ), .Y(n3681) );
  INVX1 U284 ( .A(\mem<60><3> ), .Y(n3680) );
  INVX1 U285 ( .A(\mem<60><4> ), .Y(n3679) );
  INVX1 U286 ( .A(\mem<60><5> ), .Y(n3678) );
  INVX1 U287 ( .A(\mem<60><6> ), .Y(n3677) );
  INVX1 U288 ( .A(\mem<60><7> ), .Y(n3676) );
  INVX1 U289 ( .A(\mem<59><0> ), .Y(n3675) );
  INVX1 U290 ( .A(\mem<59><1> ), .Y(n3674) );
  INVX1 U291 ( .A(\mem<59><2> ), .Y(n3673) );
  INVX1 U292 ( .A(\mem<59><3> ), .Y(n3672) );
  INVX1 U293 ( .A(\mem<59><4> ), .Y(n3671) );
  INVX1 U294 ( .A(\mem<59><5> ), .Y(n3670) );
  INVX1 U295 ( .A(\mem<59><6> ), .Y(n3669) );
  INVX1 U296 ( .A(\mem<59><7> ), .Y(n3668) );
  INVX1 U297 ( .A(\mem<58><0> ), .Y(n3667) );
  INVX1 U298 ( .A(\mem<58><1> ), .Y(n3666) );
  INVX1 U299 ( .A(\mem<58><2> ), .Y(n3665) );
  INVX1 U300 ( .A(\mem<58><3> ), .Y(n3664) );
  INVX1 U301 ( .A(\mem<58><4> ), .Y(n3663) );
  INVX1 U302 ( .A(\mem<58><5> ), .Y(n3662) );
  INVX1 U303 ( .A(\mem<58><6> ), .Y(n3661) );
  INVX1 U304 ( .A(\mem<58><7> ), .Y(n3660) );
  INVX1 U305 ( .A(\mem<57><0> ), .Y(n3659) );
  INVX1 U306 ( .A(\mem<57><1> ), .Y(n3658) );
  INVX1 U307 ( .A(\mem<57><2> ), .Y(n3657) );
  INVX1 U308 ( .A(\mem<57><3> ), .Y(n3656) );
  INVX1 U309 ( .A(\mem<57><4> ), .Y(n3655) );
  INVX1 U310 ( .A(\mem<57><5> ), .Y(n3654) );
  INVX1 U311 ( .A(\mem<57><6> ), .Y(n3653) );
  INVX1 U312 ( .A(\mem<57><7> ), .Y(n3652) );
  INVX1 U313 ( .A(\mem<56><0> ), .Y(n3651) );
  INVX1 U314 ( .A(\mem<56><1> ), .Y(n3650) );
  INVX1 U315 ( .A(\mem<56><2> ), .Y(n3649) );
  INVX1 U316 ( .A(\mem<56><3> ), .Y(n3648) );
  INVX1 U317 ( .A(\mem<56><4> ), .Y(n3647) );
  INVX1 U318 ( .A(\mem<56><5> ), .Y(n3646) );
  INVX1 U319 ( .A(\mem<56><6> ), .Y(n3645) );
  INVX1 U320 ( .A(\mem<56><7> ), .Y(n3644) );
  INVX1 U321 ( .A(\mem<55><0> ), .Y(n3643) );
  INVX1 U322 ( .A(\mem<55><1> ), .Y(n3642) );
  INVX1 U323 ( .A(\mem<55><2> ), .Y(n3641) );
  INVX1 U324 ( .A(\mem<55><3> ), .Y(n3640) );
  INVX1 U325 ( .A(\mem<55><4> ), .Y(n3639) );
  INVX1 U326 ( .A(\mem<55><5> ), .Y(n3638) );
  INVX1 U327 ( .A(\mem<55><6> ), .Y(n3637) );
  INVX1 U328 ( .A(\mem<55><7> ), .Y(n3636) );
  INVX1 U329 ( .A(\mem<54><0> ), .Y(n3635) );
  INVX1 U330 ( .A(\mem<54><1> ), .Y(n3634) );
  INVX1 U331 ( .A(\mem<54><2> ), .Y(n3633) );
  INVX1 U332 ( .A(\mem<54><3> ), .Y(n3632) );
  INVX1 U333 ( .A(\mem<54><4> ), .Y(n3631) );
  INVX1 U334 ( .A(\mem<54><5> ), .Y(n3630) );
  INVX1 U335 ( .A(\mem<54><6> ), .Y(n3629) );
  INVX1 U336 ( .A(\mem<54><7> ), .Y(n3628) );
  INVX1 U337 ( .A(\mem<53><0> ), .Y(n3627) );
  INVX1 U338 ( .A(\mem<53><1> ), .Y(n3626) );
  INVX1 U339 ( .A(\mem<53><2> ), .Y(n3625) );
  INVX1 U340 ( .A(\mem<53><3> ), .Y(n3624) );
  INVX1 U341 ( .A(\mem<53><4> ), .Y(n3623) );
  INVX1 U342 ( .A(\mem<53><5> ), .Y(n3622) );
  INVX1 U343 ( .A(\mem<53><6> ), .Y(n3621) );
  INVX1 U344 ( .A(\mem<53><7> ), .Y(n3620) );
  INVX1 U345 ( .A(\mem<52><0> ), .Y(n3619) );
  INVX1 U346 ( .A(\mem<52><1> ), .Y(n3618) );
  INVX1 U347 ( .A(\mem<52><2> ), .Y(n3617) );
  INVX1 U348 ( .A(\mem<52><3> ), .Y(n3616) );
  INVX1 U349 ( .A(\mem<52><4> ), .Y(n3615) );
  INVX1 U350 ( .A(\mem<52><5> ), .Y(n3614) );
  INVX1 U351 ( .A(\mem<52><6> ), .Y(n3613) );
  INVX1 U352 ( .A(\mem<52><7> ), .Y(n3612) );
  INVX1 U353 ( .A(\mem<51><0> ), .Y(n3611) );
  INVX1 U354 ( .A(\mem<51><1> ), .Y(n3610) );
  INVX1 U355 ( .A(\mem<51><2> ), .Y(n3609) );
  INVX1 U356 ( .A(\mem<51><3> ), .Y(n3608) );
  INVX1 U357 ( .A(\mem<51><4> ), .Y(n3607) );
  INVX1 U358 ( .A(\mem<51><5> ), .Y(n3606) );
  INVX1 U359 ( .A(\mem<51><6> ), .Y(n3605) );
  INVX1 U360 ( .A(\mem<51><7> ), .Y(n3604) );
  INVX1 U361 ( .A(\mem<50><0> ), .Y(n3603) );
  INVX1 U362 ( .A(\mem<50><1> ), .Y(n3602) );
  INVX1 U363 ( .A(\mem<50><2> ), .Y(n3601) );
  INVX1 U364 ( .A(\mem<50><3> ), .Y(n3600) );
  INVX1 U365 ( .A(\mem<50><4> ), .Y(n3599) );
  INVX1 U366 ( .A(\mem<50><5> ), .Y(n3598) );
  INVX1 U367 ( .A(\mem<50><6> ), .Y(n3597) );
  INVX1 U368 ( .A(\mem<50><7> ), .Y(n3596) );
  INVX1 U369 ( .A(\mem<49><0> ), .Y(n3595) );
  INVX1 U370 ( .A(\mem<49><1> ), .Y(n3594) );
  INVX1 U371 ( .A(\mem<49><2> ), .Y(n3593) );
  INVX1 U372 ( .A(\mem<49><3> ), .Y(n3592) );
  INVX1 U373 ( .A(\mem<49><4> ), .Y(n3591) );
  INVX1 U374 ( .A(\mem<49><5> ), .Y(n3590) );
  INVX1 U375 ( .A(\mem<49><6> ), .Y(n3589) );
  INVX1 U376 ( .A(\mem<49><7> ), .Y(n3588) );
  INVX1 U377 ( .A(\mem<48><0> ), .Y(n3587) );
  INVX1 U378 ( .A(\mem<48><1> ), .Y(n3586) );
  INVX1 U379 ( .A(\mem<48><2> ), .Y(n3585) );
  INVX1 U380 ( .A(\mem<48><3> ), .Y(n3584) );
  INVX1 U381 ( .A(\mem<48><4> ), .Y(n3583) );
  INVX1 U382 ( .A(\mem<48><5> ), .Y(n3582) );
  INVX1 U383 ( .A(\mem<48><6> ), .Y(n3581) );
  INVX1 U384 ( .A(\mem<48><7> ), .Y(n3580) );
  INVX1 U385 ( .A(\mem<47><0> ), .Y(n3579) );
  INVX1 U386 ( .A(\mem<47><1> ), .Y(n3578) );
  INVX1 U387 ( .A(\mem<47><2> ), .Y(n3577) );
  INVX1 U388 ( .A(\mem<47><3> ), .Y(n3576) );
  INVX1 U389 ( .A(\mem<47><4> ), .Y(n3575) );
  INVX1 U390 ( .A(\mem<47><5> ), .Y(n3574) );
  INVX1 U391 ( .A(\mem<47><6> ), .Y(n3573) );
  INVX1 U392 ( .A(\mem<47><7> ), .Y(n3572) );
  INVX1 U393 ( .A(\mem<46><0> ), .Y(n3571) );
  INVX1 U394 ( .A(\mem<46><1> ), .Y(n3570) );
  INVX1 U395 ( .A(\mem<46><2> ), .Y(n3569) );
  INVX1 U396 ( .A(\mem<46><3> ), .Y(n3568) );
  INVX1 U397 ( .A(\mem<46><4> ), .Y(n3567) );
  INVX1 U398 ( .A(\mem<46><5> ), .Y(n3566) );
  INVX1 U399 ( .A(\mem<46><6> ), .Y(n3565) );
  INVX1 U400 ( .A(\mem<46><7> ), .Y(n3564) );
  INVX1 U401 ( .A(\mem<45><0> ), .Y(n3563) );
  INVX1 U402 ( .A(\mem<45><1> ), .Y(n3562) );
  INVX1 U403 ( .A(\mem<45><2> ), .Y(n3561) );
  INVX1 U404 ( .A(\mem<45><3> ), .Y(n3560) );
  INVX1 U405 ( .A(\mem<45><4> ), .Y(n3559) );
  INVX1 U406 ( .A(\mem<45><5> ), .Y(n3558) );
  INVX1 U407 ( .A(\mem<45><6> ), .Y(n3557) );
  INVX1 U408 ( .A(\mem<45><7> ), .Y(n3556) );
  INVX1 U409 ( .A(\mem<44><0> ), .Y(n3555) );
  INVX1 U410 ( .A(\mem<44><1> ), .Y(n3554) );
  INVX1 U411 ( .A(\mem<44><2> ), .Y(n3553) );
  INVX1 U412 ( .A(\mem<44><3> ), .Y(n3552) );
  INVX1 U413 ( .A(\mem<44><4> ), .Y(n3551) );
  INVX1 U414 ( .A(\mem<44><5> ), .Y(n3550) );
  INVX1 U415 ( .A(\mem<44><6> ), .Y(n3549) );
  INVX1 U416 ( .A(\mem<44><7> ), .Y(n3548) );
  INVX1 U417 ( .A(\mem<43><0> ), .Y(n3547) );
  INVX1 U418 ( .A(\mem<43><1> ), .Y(n3546) );
  INVX1 U419 ( .A(\mem<43><2> ), .Y(n3545) );
  INVX1 U420 ( .A(\mem<43><3> ), .Y(n3544) );
  INVX1 U421 ( .A(\mem<43><4> ), .Y(n3543) );
  INVX1 U422 ( .A(\mem<43><5> ), .Y(n3542) );
  INVX1 U423 ( .A(\mem<43><6> ), .Y(n3541) );
  INVX1 U424 ( .A(\mem<43><7> ), .Y(n3540) );
  INVX1 U425 ( .A(\mem<42><0> ), .Y(n3539) );
  INVX1 U426 ( .A(\mem<42><1> ), .Y(n3538) );
  INVX1 U427 ( .A(\mem<42><2> ), .Y(n3537) );
  INVX1 U428 ( .A(\mem<42><3> ), .Y(n3536) );
  INVX1 U429 ( .A(\mem<42><4> ), .Y(n3535) );
  INVX1 U430 ( .A(\mem<42><5> ), .Y(n3534) );
  INVX1 U431 ( .A(\mem<42><6> ), .Y(n3533) );
  INVX1 U432 ( .A(\mem<42><7> ), .Y(n3532) );
  INVX1 U433 ( .A(\mem<41><0> ), .Y(n3531) );
  INVX1 U434 ( .A(\mem<41><1> ), .Y(n3530) );
  INVX1 U435 ( .A(\mem<41><2> ), .Y(n3529) );
  INVX1 U436 ( .A(\mem<41><3> ), .Y(n3528) );
  INVX1 U437 ( .A(\mem<41><4> ), .Y(n3527) );
  INVX1 U438 ( .A(\mem<41><5> ), .Y(n3526) );
  INVX1 U439 ( .A(\mem<41><6> ), .Y(n3525) );
  INVX1 U440 ( .A(\mem<41><7> ), .Y(n3524) );
  INVX1 U441 ( .A(\mem<40><0> ), .Y(n3523) );
  INVX1 U442 ( .A(\mem<40><1> ), .Y(n3522) );
  INVX1 U443 ( .A(\mem<40><2> ), .Y(n3521) );
  INVX1 U444 ( .A(\mem<40><3> ), .Y(n3520) );
  INVX1 U445 ( .A(\mem<40><4> ), .Y(n3519) );
  INVX1 U446 ( .A(\mem<40><5> ), .Y(n3518) );
  INVX1 U447 ( .A(\mem<40><6> ), .Y(n3517) );
  INVX1 U448 ( .A(\mem<40><7> ), .Y(n3516) );
  INVX1 U449 ( .A(\mem<39><0> ), .Y(n3515) );
  INVX1 U450 ( .A(\mem<39><1> ), .Y(n3514) );
  INVX1 U451 ( .A(\mem<39><2> ), .Y(n3513) );
  INVX1 U452 ( .A(\mem<39><3> ), .Y(n3512) );
  INVX1 U453 ( .A(\mem<39><4> ), .Y(n3511) );
  INVX1 U454 ( .A(\mem<39><5> ), .Y(n3510) );
  INVX1 U455 ( .A(\mem<39><6> ), .Y(n3509) );
  INVX1 U456 ( .A(\mem<39><7> ), .Y(n3508) );
  INVX1 U457 ( .A(\mem<38><0> ), .Y(n3507) );
  INVX1 U458 ( .A(\mem<38><1> ), .Y(n3506) );
  INVX1 U459 ( .A(\mem<38><2> ), .Y(n3505) );
  INVX1 U460 ( .A(\mem<38><3> ), .Y(n3504) );
  INVX1 U461 ( .A(\mem<38><4> ), .Y(n3503) );
  INVX1 U462 ( .A(\mem<38><5> ), .Y(n3502) );
  INVX1 U463 ( .A(\mem<38><6> ), .Y(n3501) );
  INVX1 U464 ( .A(\mem<38><7> ), .Y(n3500) );
  INVX1 U465 ( .A(\mem<37><0> ), .Y(n3499) );
  INVX1 U466 ( .A(\mem<37><1> ), .Y(n3498) );
  INVX1 U467 ( .A(\mem<37><2> ), .Y(n3497) );
  INVX1 U468 ( .A(\mem<37><3> ), .Y(n3496) );
  INVX1 U469 ( .A(\mem<37><4> ), .Y(n3495) );
  INVX1 U470 ( .A(\mem<37><5> ), .Y(n3494) );
  INVX1 U471 ( .A(\mem<37><6> ), .Y(n3493) );
  INVX1 U472 ( .A(\mem<37><7> ), .Y(n3492) );
  INVX1 U473 ( .A(\mem<36><0> ), .Y(n3491) );
  INVX1 U474 ( .A(\mem<36><1> ), .Y(n3490) );
  INVX1 U475 ( .A(\mem<36><2> ), .Y(n3489) );
  INVX1 U476 ( .A(\mem<36><3> ), .Y(n3488) );
  INVX1 U477 ( .A(\mem<36><4> ), .Y(n3487) );
  INVX1 U478 ( .A(\mem<36><5> ), .Y(n3486) );
  INVX1 U479 ( .A(\mem<36><6> ), .Y(n3485) );
  INVX1 U480 ( .A(\mem<36><7> ), .Y(n3484) );
  INVX1 U481 ( .A(\mem<35><0> ), .Y(n3483) );
  INVX1 U482 ( .A(\mem<35><1> ), .Y(n3482) );
  INVX1 U483 ( .A(\mem<35><2> ), .Y(n3481) );
  INVX1 U484 ( .A(\mem<35><3> ), .Y(n3480) );
  INVX1 U485 ( .A(\mem<35><4> ), .Y(n3479) );
  INVX1 U486 ( .A(\mem<35><5> ), .Y(n3478) );
  INVX1 U487 ( .A(\mem<35><6> ), .Y(n3477) );
  INVX1 U488 ( .A(\mem<35><7> ), .Y(n3476) );
  INVX1 U489 ( .A(\mem<34><0> ), .Y(n3475) );
  INVX1 U490 ( .A(\mem<34><1> ), .Y(n3474) );
  INVX1 U491 ( .A(\mem<34><2> ), .Y(n3473) );
  INVX1 U492 ( .A(\mem<34><3> ), .Y(n3472) );
  INVX1 U493 ( .A(\mem<34><4> ), .Y(n3471) );
  INVX1 U494 ( .A(\mem<34><5> ), .Y(n3470) );
  INVX1 U495 ( .A(\mem<34><6> ), .Y(n3469) );
  INVX1 U496 ( .A(\mem<34><7> ), .Y(n3468) );
  INVX1 U497 ( .A(\mem<33><0> ), .Y(n3467) );
  INVX1 U498 ( .A(\mem<33><1> ), .Y(n3466) );
  INVX1 U499 ( .A(\mem<33><2> ), .Y(n3465) );
  INVX1 U500 ( .A(\mem<33><3> ), .Y(n3464) );
  INVX1 U501 ( .A(\mem<33><4> ), .Y(n3463) );
  INVX1 U502 ( .A(\mem<33><5> ), .Y(n3462) );
  INVX1 U503 ( .A(\mem<33><6> ), .Y(n3461) );
  INVX1 U504 ( .A(\mem<33><7> ), .Y(n3460) );
  INVX1 U505 ( .A(\mem<32><0> ), .Y(n3459) );
  INVX1 U506 ( .A(\mem<32><1> ), .Y(n3458) );
  INVX1 U507 ( .A(\mem<32><2> ), .Y(n3457) );
  INVX1 U508 ( .A(\mem<32><3> ), .Y(n3456) );
  INVX1 U509 ( .A(\mem<32><4> ), .Y(n3455) );
  INVX1 U510 ( .A(\mem<32><5> ), .Y(n3454) );
  INVX1 U511 ( .A(\mem<32><6> ), .Y(n3453) );
  INVX1 U512 ( .A(\mem<32><7> ), .Y(n3452) );
  INVX1 U513 ( .A(\mem<31><0> ), .Y(n3451) );
  INVX1 U514 ( .A(\mem<31><1> ), .Y(n3450) );
  INVX1 U515 ( .A(\mem<31><2> ), .Y(n3449) );
  INVX1 U516 ( .A(\mem<31><3> ), .Y(n3448) );
  INVX1 U517 ( .A(\mem<31><4> ), .Y(n3447) );
  INVX1 U518 ( .A(\mem<31><5> ), .Y(n3446) );
  INVX1 U519 ( .A(\mem<31><6> ), .Y(n3445) );
  INVX1 U520 ( .A(\mem<31><7> ), .Y(n3444) );
  INVX1 U521 ( .A(\mem<30><0> ), .Y(n3443) );
  INVX1 U522 ( .A(\mem<30><1> ), .Y(n3442) );
  INVX1 U523 ( .A(\mem<30><2> ), .Y(n3441) );
  INVX1 U524 ( .A(\mem<30><3> ), .Y(n3440) );
  INVX1 U525 ( .A(\mem<30><4> ), .Y(n3439) );
  INVX1 U526 ( .A(\mem<30><5> ), .Y(n3438) );
  INVX1 U527 ( .A(\mem<30><6> ), .Y(n3437) );
  INVX1 U528 ( .A(\mem<30><7> ), .Y(n3436) );
  INVX1 U529 ( .A(\mem<29><0> ), .Y(n3435) );
  INVX1 U530 ( .A(\mem<29><1> ), .Y(n3434) );
  INVX1 U531 ( .A(\mem<29><2> ), .Y(n3433) );
  INVX1 U532 ( .A(\mem<29><3> ), .Y(n3432) );
  INVX1 U533 ( .A(\mem<29><4> ), .Y(n3431) );
  INVX1 U534 ( .A(\mem<29><5> ), .Y(n3430) );
  INVX1 U535 ( .A(\mem<29><6> ), .Y(n3429) );
  INVX1 U536 ( .A(\mem<29><7> ), .Y(n3428) );
  INVX1 U537 ( .A(\mem<28><0> ), .Y(n3427) );
  INVX1 U538 ( .A(\mem<28><1> ), .Y(n3426) );
  INVX1 U539 ( .A(\mem<28><2> ), .Y(n3425) );
  INVX1 U540 ( .A(\mem<28><3> ), .Y(n3424) );
  INVX1 U541 ( .A(\mem<28><4> ), .Y(n3423) );
  INVX1 U542 ( .A(\mem<28><5> ), .Y(n3422) );
  INVX1 U543 ( .A(\mem<28><6> ), .Y(n3421) );
  INVX1 U544 ( .A(\mem<28><7> ), .Y(n3420) );
  INVX1 U545 ( .A(\mem<27><0> ), .Y(n3419) );
  INVX1 U546 ( .A(\mem<27><1> ), .Y(n3418) );
  INVX1 U547 ( .A(\mem<27><2> ), .Y(n3417) );
  INVX1 U548 ( .A(\mem<27><3> ), .Y(n3416) );
  INVX1 U549 ( .A(\mem<27><4> ), .Y(n3415) );
  INVX1 U550 ( .A(\mem<27><5> ), .Y(n3414) );
  INVX1 U551 ( .A(\mem<27><6> ), .Y(n3413) );
  INVX1 U552 ( .A(\mem<27><7> ), .Y(n3412) );
  INVX1 U553 ( .A(\mem<26><0> ), .Y(n3411) );
  INVX1 U554 ( .A(\mem<26><1> ), .Y(n3410) );
  INVX1 U555 ( .A(\mem<26><2> ), .Y(n3409) );
  INVX1 U556 ( .A(\mem<26><3> ), .Y(n3408) );
  INVX1 U557 ( .A(\mem<26><4> ), .Y(n3407) );
  INVX1 U558 ( .A(\mem<26><5> ), .Y(n3406) );
  INVX1 U559 ( .A(\mem<26><6> ), .Y(n3405) );
  INVX1 U560 ( .A(\mem<26><7> ), .Y(n3404) );
  INVX1 U561 ( .A(\mem<25><0> ), .Y(n3403) );
  INVX1 U562 ( .A(\mem<25><1> ), .Y(n3402) );
  INVX1 U563 ( .A(\mem<25><2> ), .Y(n3401) );
  INVX1 U564 ( .A(\mem<25><3> ), .Y(n3400) );
  INVX1 U565 ( .A(\mem<25><4> ), .Y(n3399) );
  INVX1 U566 ( .A(\mem<25><5> ), .Y(n3398) );
  INVX1 U567 ( .A(\mem<25><6> ), .Y(n3397) );
  INVX1 U568 ( .A(\mem<25><7> ), .Y(n3396) );
  INVX1 U569 ( .A(\mem<24><0> ), .Y(n3395) );
  INVX1 U570 ( .A(\mem<24><1> ), .Y(n3394) );
  INVX1 U571 ( .A(\mem<24><2> ), .Y(n3393) );
  INVX1 U572 ( .A(\mem<24><3> ), .Y(n3392) );
  INVX1 U573 ( .A(\mem<24><4> ), .Y(n3391) );
  INVX1 U574 ( .A(\mem<24><5> ), .Y(n3390) );
  INVX1 U575 ( .A(\mem<24><6> ), .Y(n3389) );
  INVX1 U576 ( .A(\mem<24><7> ), .Y(n3388) );
  INVX1 U577 ( .A(\mem<23><0> ), .Y(n3387) );
  INVX1 U578 ( .A(\mem<23><1> ), .Y(n3386) );
  INVX1 U579 ( .A(\mem<23><2> ), .Y(n3385) );
  INVX1 U580 ( .A(\mem<23><3> ), .Y(n3384) );
  INVX1 U581 ( .A(\mem<23><4> ), .Y(n3383) );
  INVX1 U582 ( .A(\mem<23><5> ), .Y(n3382) );
  INVX1 U583 ( .A(\mem<23><6> ), .Y(n3381) );
  INVX1 U584 ( .A(\mem<23><7> ), .Y(n3380) );
  INVX1 U585 ( .A(\mem<22><0> ), .Y(n3379) );
  INVX1 U586 ( .A(\mem<22><1> ), .Y(n3378) );
  INVX1 U587 ( .A(\mem<22><2> ), .Y(n3377) );
  INVX1 U588 ( .A(\mem<22><3> ), .Y(n3376) );
  INVX1 U589 ( .A(\mem<22><4> ), .Y(n3375) );
  INVX1 U590 ( .A(\mem<22><5> ), .Y(n3374) );
  INVX1 U591 ( .A(\mem<22><6> ), .Y(n3373) );
  INVX1 U592 ( .A(\mem<22><7> ), .Y(n3372) );
  INVX1 U593 ( .A(\mem<21><0> ), .Y(n3371) );
  INVX1 U594 ( .A(\mem<21><1> ), .Y(n3370) );
  INVX1 U595 ( .A(\mem<21><2> ), .Y(n3369) );
  INVX1 U596 ( .A(\mem<21><3> ), .Y(n3368) );
  INVX1 U597 ( .A(\mem<21><4> ), .Y(n3367) );
  INVX1 U598 ( .A(\mem<21><5> ), .Y(n3366) );
  INVX1 U599 ( .A(\mem<21><6> ), .Y(n3365) );
  INVX1 U600 ( .A(\mem<21><7> ), .Y(n3364) );
  INVX1 U601 ( .A(\mem<20><0> ), .Y(n3363) );
  INVX1 U602 ( .A(\mem<20><1> ), .Y(n3362) );
  INVX1 U603 ( .A(\mem<20><2> ), .Y(n3361) );
  INVX1 U604 ( .A(\mem<20><3> ), .Y(n3360) );
  INVX1 U605 ( .A(\mem<20><4> ), .Y(n3359) );
  INVX1 U606 ( .A(\mem<20><5> ), .Y(n3358) );
  INVX1 U607 ( .A(\mem<20><6> ), .Y(n3357) );
  INVX1 U608 ( .A(\mem<20><7> ), .Y(n3356) );
  INVX1 U609 ( .A(\mem<19><0> ), .Y(n3355) );
  INVX1 U610 ( .A(\mem<19><1> ), .Y(n3354) );
  INVX1 U611 ( .A(\mem<19><2> ), .Y(n3353) );
  INVX1 U612 ( .A(\mem<19><3> ), .Y(n3352) );
  INVX1 U613 ( .A(\mem<19><4> ), .Y(n3351) );
  INVX1 U614 ( .A(\mem<19><5> ), .Y(n3350) );
  INVX1 U615 ( .A(\mem<19><6> ), .Y(n3349) );
  INVX1 U616 ( .A(\mem<19><7> ), .Y(n3348) );
  INVX1 U617 ( .A(\mem<18><0> ), .Y(n3347) );
  INVX1 U618 ( .A(\mem<18><1> ), .Y(n3346) );
  INVX1 U619 ( .A(\mem<18><2> ), .Y(n3345) );
  INVX1 U620 ( .A(\mem<18><3> ), .Y(n3344) );
  INVX1 U621 ( .A(\mem<18><4> ), .Y(n3343) );
  INVX1 U622 ( .A(\mem<18><5> ), .Y(n3342) );
  INVX1 U623 ( .A(\mem<18><6> ), .Y(n3341) );
  INVX1 U624 ( .A(\mem<18><7> ), .Y(n3340) );
  INVX1 U625 ( .A(\mem<17><0> ), .Y(n3339) );
  INVX1 U626 ( .A(\mem<17><1> ), .Y(n3338) );
  INVX1 U627 ( .A(\mem<17><2> ), .Y(n3337) );
  INVX1 U628 ( .A(\mem<17><3> ), .Y(n3336) );
  INVX1 U629 ( .A(\mem<17><4> ), .Y(n3335) );
  INVX1 U630 ( .A(\mem<17><5> ), .Y(n3334) );
  INVX1 U631 ( .A(\mem<17><6> ), .Y(n3333) );
  INVX1 U632 ( .A(\mem<17><7> ), .Y(n3332) );
  INVX1 U633 ( .A(\mem<16><0> ), .Y(n3331) );
  INVX1 U634 ( .A(\mem<16><1> ), .Y(n3330) );
  INVX1 U635 ( .A(\mem<16><2> ), .Y(n3329) );
  INVX1 U636 ( .A(\mem<16><3> ), .Y(n3328) );
  INVX1 U637 ( .A(\mem<16><4> ), .Y(n3327) );
  INVX1 U638 ( .A(\mem<16><5> ), .Y(n3326) );
  INVX1 U639 ( .A(\mem<16><6> ), .Y(n3325) );
  INVX1 U640 ( .A(\mem<16><7> ), .Y(n3324) );
  INVX1 U641 ( .A(\mem<15><0> ), .Y(n3323) );
  INVX1 U642 ( .A(\mem<15><1> ), .Y(n3322) );
  INVX1 U643 ( .A(\mem<15><2> ), .Y(n3321) );
  INVX1 U644 ( .A(\mem<15><3> ), .Y(n3320) );
  INVX1 U645 ( .A(\mem<15><4> ), .Y(n3319) );
  INVX1 U646 ( .A(\mem<15><5> ), .Y(n3318) );
  INVX1 U647 ( .A(\mem<15><6> ), .Y(n3317) );
  INVX1 U648 ( .A(\mem<15><7> ), .Y(n3316) );
  INVX1 U649 ( .A(\mem<14><0> ), .Y(n3315) );
  INVX1 U650 ( .A(\mem<14><1> ), .Y(n3314) );
  INVX1 U651 ( .A(\mem<14><2> ), .Y(n3313) );
  INVX1 U652 ( .A(\mem<14><3> ), .Y(n3312) );
  INVX1 U653 ( .A(\mem<14><4> ), .Y(n3311) );
  INVX1 U654 ( .A(\mem<14><5> ), .Y(n3310) );
  INVX1 U655 ( .A(\mem<14><6> ), .Y(n3309) );
  INVX1 U656 ( .A(\mem<14><7> ), .Y(n3308) );
  INVX1 U657 ( .A(\mem<13><0> ), .Y(n3307) );
  INVX1 U658 ( .A(\mem<13><1> ), .Y(n3306) );
  INVX1 U659 ( .A(\mem<13><2> ), .Y(n3305) );
  INVX1 U660 ( .A(\mem<13><3> ), .Y(n3304) );
  INVX1 U661 ( .A(\mem<13><4> ), .Y(n3303) );
  INVX1 U662 ( .A(\mem<13><5> ), .Y(n3302) );
  INVX1 U663 ( .A(\mem<13><6> ), .Y(n3301) );
  INVX1 U664 ( .A(\mem<13><7> ), .Y(n3300) );
  INVX1 U665 ( .A(\mem<12><0> ), .Y(n3299) );
  INVX1 U666 ( .A(\mem<12><1> ), .Y(n3298) );
  INVX1 U667 ( .A(\mem<12><2> ), .Y(n3297) );
  INVX1 U668 ( .A(\mem<12><3> ), .Y(n3296) );
  INVX1 U669 ( .A(\mem<12><4> ), .Y(n3295) );
  INVX1 U670 ( .A(\mem<12><5> ), .Y(n3294) );
  INVX1 U671 ( .A(\mem<12><6> ), .Y(n3293) );
  INVX1 U672 ( .A(\mem<12><7> ), .Y(n3292) );
  INVX1 U673 ( .A(\mem<11><0> ), .Y(n3291) );
  INVX1 U674 ( .A(\mem<11><1> ), .Y(n3290) );
  INVX1 U675 ( .A(\mem<11><2> ), .Y(n3289) );
  INVX1 U676 ( .A(\mem<11><3> ), .Y(n3288) );
  INVX1 U677 ( .A(\mem<11><4> ), .Y(n3287) );
  INVX1 U678 ( .A(\mem<11><5> ), .Y(n3286) );
  INVX1 U679 ( .A(\mem<11><6> ), .Y(n3285) );
  INVX1 U680 ( .A(\mem<11><7> ), .Y(n3284) );
  INVX1 U681 ( .A(\mem<10><0> ), .Y(n3283) );
  INVX1 U682 ( .A(\mem<10><1> ), .Y(n3282) );
  INVX1 U683 ( .A(\mem<10><2> ), .Y(n3281) );
  INVX1 U684 ( .A(\mem<10><3> ), .Y(n3280) );
  INVX1 U685 ( .A(\mem<10><4> ), .Y(n3279) );
  INVX1 U686 ( .A(\mem<10><5> ), .Y(n3278) );
  INVX1 U687 ( .A(\mem<10><6> ), .Y(n3277) );
  INVX1 U688 ( .A(\mem<10><7> ), .Y(n3276) );
  INVX1 U689 ( .A(\mem<9><0> ), .Y(n3275) );
  INVX1 U690 ( .A(\mem<9><1> ), .Y(n3274) );
  INVX1 U691 ( .A(\mem<9><2> ), .Y(n3273) );
  INVX1 U692 ( .A(\mem<9><3> ), .Y(n3272) );
  INVX1 U693 ( .A(\mem<9><4> ), .Y(n3271) );
  INVX1 U694 ( .A(\mem<9><5> ), .Y(n3270) );
  INVX1 U695 ( .A(\mem<9><6> ), .Y(n3269) );
  INVX1 U696 ( .A(\mem<9><7> ), .Y(n3268) );
  INVX1 U697 ( .A(\mem<8><0> ), .Y(n3267) );
  INVX1 U698 ( .A(\mem<8><1> ), .Y(n3266) );
  INVX1 U699 ( .A(\mem<8><2> ), .Y(n3265) );
  INVX1 U700 ( .A(\mem<8><3> ), .Y(n3264) );
  INVX1 U701 ( .A(\mem<8><4> ), .Y(n3263) );
  INVX1 U702 ( .A(\mem<8><5> ), .Y(n3262) );
  INVX1 U703 ( .A(\mem<8><6> ), .Y(n3261) );
  INVX1 U704 ( .A(\mem<8><7> ), .Y(n3260) );
  INVX1 U705 ( .A(\mem<7><0> ), .Y(n3259) );
  INVX1 U706 ( .A(\mem<7><1> ), .Y(n3258) );
  INVX1 U707 ( .A(\mem<7><2> ), .Y(n3257) );
  INVX1 U708 ( .A(\mem<7><3> ), .Y(n3256) );
  INVX1 U709 ( .A(\mem<7><4> ), .Y(n3255) );
  INVX1 U710 ( .A(\mem<7><5> ), .Y(n3254) );
  INVX1 U711 ( .A(\mem<7><6> ), .Y(n3253) );
  INVX1 U712 ( .A(\mem<7><7> ), .Y(n3252) );
  INVX1 U713 ( .A(\mem<6><0> ), .Y(n3251) );
  INVX1 U714 ( .A(\mem<6><1> ), .Y(n3250) );
  INVX1 U715 ( .A(\mem<6><2> ), .Y(n3249) );
  INVX1 U716 ( .A(\mem<6><3> ), .Y(n3248) );
  INVX1 U717 ( .A(\mem<6><4> ), .Y(n3247) );
  INVX1 U718 ( .A(\mem<6><5> ), .Y(n3246) );
  INVX1 U719 ( .A(\mem<6><6> ), .Y(n3245) );
  INVX1 U720 ( .A(\mem<6><7> ), .Y(n3244) );
  INVX1 U721 ( .A(\mem<5><0> ), .Y(n3243) );
  INVX1 U722 ( .A(\mem<5><1> ), .Y(n3242) );
  INVX1 U723 ( .A(\mem<5><2> ), .Y(n3241) );
  INVX1 U724 ( .A(\mem<5><3> ), .Y(n3240) );
  INVX1 U725 ( .A(\mem<5><4> ), .Y(n3239) );
  INVX1 U726 ( .A(\mem<5><5> ), .Y(n3238) );
  INVX1 U727 ( .A(\mem<5><6> ), .Y(n3237) );
  INVX1 U728 ( .A(\mem<5><7> ), .Y(n3236) );
  INVX1 U729 ( .A(\mem<4><0> ), .Y(n3235) );
  INVX1 U730 ( .A(\mem<4><1> ), .Y(n3234) );
  INVX1 U731 ( .A(\mem<4><2> ), .Y(n3233) );
  INVX1 U732 ( .A(\mem<4><3> ), .Y(n3232) );
  INVX1 U733 ( .A(\mem<4><4> ), .Y(n3231) );
  INVX1 U734 ( .A(\mem<4><5> ), .Y(n3230) );
  INVX1 U735 ( .A(\mem<4><6> ), .Y(n3229) );
  INVX1 U736 ( .A(\mem<4><7> ), .Y(n3228) );
  INVX1 U737 ( .A(\mem<3><0> ), .Y(n3227) );
  INVX1 U738 ( .A(\mem<3><1> ), .Y(n3226) );
  INVX1 U739 ( .A(\mem<3><2> ), .Y(n3225) );
  INVX1 U740 ( .A(\mem<3><3> ), .Y(n3224) );
  INVX1 U741 ( .A(\mem<3><4> ), .Y(n3223) );
  INVX1 U742 ( .A(\mem<3><5> ), .Y(n3222) );
  INVX1 U743 ( .A(\mem<3><6> ), .Y(n3221) );
  INVX1 U744 ( .A(\mem<3><7> ), .Y(n3220) );
  INVX1 U745 ( .A(\mem<2><0> ), .Y(n3219) );
  INVX1 U746 ( .A(\mem<2><1> ), .Y(n3218) );
  INVX1 U747 ( .A(\mem<2><2> ), .Y(n3217) );
  INVX1 U748 ( .A(\mem<2><3> ), .Y(n3216) );
  INVX1 U749 ( .A(\mem<2><4> ), .Y(n3215) );
  INVX1 U750 ( .A(\mem<2><5> ), .Y(n3214) );
  INVX1 U751 ( .A(\mem<2><6> ), .Y(n3213) );
  INVX1 U752 ( .A(\mem<2><7> ), .Y(n3212) );
  INVX1 U753 ( .A(\mem<1><0> ), .Y(n3211) );
  INVX1 U754 ( .A(\mem<1><1> ), .Y(n3210) );
  INVX1 U755 ( .A(\mem<1><2> ), .Y(n3209) );
  INVX1 U756 ( .A(\mem<1><3> ), .Y(n3208) );
  INVX1 U757 ( .A(\mem<1><4> ), .Y(n3207) );
  INVX1 U758 ( .A(\mem<1><5> ), .Y(n3206) );
  INVX1 U759 ( .A(\mem<1><6> ), .Y(n3205) );
  INVX1 U760 ( .A(\mem<1><7> ), .Y(n3204) );
  INVX1 U761 ( .A(\mem<0><0> ), .Y(n3203) );
  INVX1 U762 ( .A(\mem<0><1> ), .Y(n3202) );
  INVX1 U763 ( .A(\mem<0><2> ), .Y(n3201) );
  INVX1 U764 ( .A(\mem<0><3> ), .Y(n3200) );
  INVX1 U765 ( .A(\mem<0><4> ), .Y(n3199) );
  INVX1 U766 ( .A(\mem<0><5> ), .Y(n3198) );
  INVX1 U767 ( .A(\mem<0><6> ), .Y(n3197) );
  INVX1 U768 ( .A(\mem<0><7> ), .Y(n3196) );
  INVX1 U769 ( .A(n3112), .Y(n3092) );
  INVX1 U770 ( .A(n3112), .Y(n3090) );
  INVX1 U771 ( .A(n3112), .Y(n3091) );
  INVX1 U772 ( .A(n3112), .Y(n3093) );
  INVX1 U773 ( .A(n3181), .Y(n3098) );
  INVX1 U774 ( .A(n3181), .Y(n3096) );
  INVX1 U775 ( .A(n3183), .Y(n3087) );
  INVX1 U776 ( .A(n3183), .Y(n3088) );
  INVX1 U777 ( .A(n3183), .Y(n3086) );
  INVX1 U778 ( .A(n3181), .Y(n3094) );
  INVX1 U779 ( .A(n3181), .Y(n3095) );
  INVX1 U780 ( .A(n3183), .Y(n3083) );
  INVX1 U781 ( .A(n3183), .Y(n3089) );
  INVX1 U782 ( .A(n3092), .Y(n3099) );
  INVX1 U783 ( .A(n3090), .Y(n3100) );
  INVX1 U784 ( .A(n3091), .Y(n3097) );
  INVX1 U785 ( .A(n3184), .Y(n3082) );
  INVX1 U786 ( .A(n3184), .Y(n3081) );
  INVX1 U787 ( .A(N178), .Y(n3183) );
  INVX1 U788 ( .A(n3183), .Y(n3084) );
  INVX1 U789 ( .A(n3183), .Y(n3085) );
  OR2X1 U790 ( .A(n2407), .B(n210), .Y(n181) );
  OR2X1 U791 ( .A(n2413), .B(n213), .Y(n182) );
  OR2X1 U792 ( .A(n2419), .B(n216), .Y(n183) );
  OR2X1 U793 ( .A(n2425), .B(n219), .Y(n184) );
  OR2X1 U794 ( .A(n2431), .B(n222), .Y(n185) );
  OR2X1 U795 ( .A(n2437), .B(n225), .Y(n186) );
  OR2X1 U796 ( .A(n2443), .B(n228), .Y(n187) );
  OR2X1 U797 ( .A(n2449), .B(n231), .Y(n188) );
  INVX1 U798 ( .A(N180), .Y(n3185) );
  INVX1 U799 ( .A(N177), .Y(n3181) );
  OR2X1 U800 ( .A(n2356), .B(n192), .Y(n165) );
  OR2X1 U801 ( .A(n2359), .B(n193), .Y(n166) );
  OR2X1 U802 ( .A(n2362), .B(n194), .Y(n167) );
  OR2X1 U803 ( .A(n2365), .B(n195), .Y(n168) );
  OR2X1 U804 ( .A(n2368), .B(n196), .Y(n169) );
  OR2X1 U805 ( .A(n2371), .B(n197), .Y(n170) );
  OR2X1 U806 ( .A(n2374), .B(n198), .Y(n171) );
  OR2X1 U807 ( .A(n2377), .B(n199), .Y(n172) );
  OR2X1 U808 ( .A(n2380), .B(n200), .Y(n173) );
  OR2X1 U809 ( .A(n2383), .B(n201), .Y(n174) );
  OR2X1 U810 ( .A(n2386), .B(n202), .Y(n175) );
  OR2X1 U811 ( .A(n2389), .B(n203), .Y(n176) );
  OR2X1 U812 ( .A(n2392), .B(n204), .Y(n177) );
  OR2X1 U813 ( .A(n2395), .B(n205), .Y(n178) );
  OR2X1 U814 ( .A(n2398), .B(n206), .Y(n179) );
  OR2X1 U815 ( .A(n2401), .B(n207), .Y(n180) );
  OR2X1 U816 ( .A(n189), .B(n3185), .Y(n190) );
  OR2X1 U1889 ( .A(n10), .B(n7), .Y(n6) );
  OR2X1 U1891 ( .A(n20), .B(n17), .Y(n16) );
  OR2X1 U1893 ( .A(n30), .B(n27), .Y(n26) );
  OR2X1 U1895 ( .A(n40), .B(n37), .Y(n36) );
  OR2X1 U1897 ( .A(n50), .B(n47), .Y(n46) );
  OR2X1 U1899 ( .A(n60), .B(n57), .Y(n56) );
  OR2X1 U1901 ( .A(n70), .B(n67), .Y(n66) );
  OR2X1 U1903 ( .A(n80), .B(n77), .Y(n76) );
  OR2X1 U1904 ( .A(n90), .B(n87), .Y(n86) );
  OR2X1 U1908 ( .A(n100), .B(n97), .Y(n96) );
  OR2X1 U1913 ( .A(n110), .B(n107), .Y(n106) );
  OR2X1 U1918 ( .A(n120), .B(n117), .Y(n116) );
  OR2X1 U1923 ( .A(n130), .B(n127), .Y(n126) );
  OR2X1 U1929 ( .A(n140), .B(n137), .Y(n136) );
  OR2X1 U1934 ( .A(n150), .B(n147), .Y(n146) );
  OR2X1 U1939 ( .A(n160), .B(n157), .Y(n156) );
  INVX1 U1944 ( .A(n3181), .Y(n3112) );
  INVX1 U1951 ( .A(N179), .Y(n3184) );
  INVX1 U1956 ( .A(n3183), .Y(n3182) );
  OR2X1 U1961 ( .A(n3), .B(n4), .Y(n2) );
  OR2X1 U1966 ( .A(n13), .B(n14), .Y(n12) );
  OR2X1 U1972 ( .A(n23), .B(n24), .Y(n22) );
  OR2X1 U1977 ( .A(n33), .B(n34), .Y(n32) );
  OR2X1 U1982 ( .A(n43), .B(n44), .Y(n42) );
  OR2X1 U1987 ( .A(n53), .B(n54), .Y(n52) );
  OR2X1 U1994 ( .A(n63), .B(n64), .Y(n62) );
  OR2X1 U1999 ( .A(n73), .B(n74), .Y(n72) );
  OR2X1 U2004 ( .A(n83), .B(n84), .Y(n82) );
  OR2X1 U2009 ( .A(n93), .B(n94), .Y(n92) );
  OR2X1 U2015 ( .A(n103), .B(n104), .Y(n102) );
  OR2X1 U2020 ( .A(n113), .B(n114), .Y(n112) );
  OR2X1 U2025 ( .A(n123), .B(n124), .Y(n122) );
  OR2X1 U2030 ( .A(n133), .B(n134), .Y(n132) );
  OR2X1 U2037 ( .A(n143), .B(n144), .Y(n142) );
  OR2X1 U2042 ( .A(n153), .B(n154), .Y(n152) );
  OR2X1 U2047 ( .A(n5), .B(n2), .Y(n1) );
  OR2X1 U2052 ( .A(n15), .B(n12), .Y(n11) );
  OR2X1 U2058 ( .A(n25), .B(n22), .Y(n21) );
  OR2X1 U2063 ( .A(n35), .B(n32), .Y(n31) );
  OR2X1 U2068 ( .A(n45), .B(n42), .Y(n41) );
  OR2X1 U2073 ( .A(n55), .B(n52), .Y(n51) );
  OR2X1 U2080 ( .A(n65), .B(n62), .Y(n61) );
  OR2X1 U2085 ( .A(n75), .B(n72), .Y(n71) );
  OR2X1 U2090 ( .A(n85), .B(n82), .Y(n81) );
  OR2X1 U2095 ( .A(n95), .B(n92), .Y(n91) );
  OR2X1 U2101 ( .A(n105), .B(n102), .Y(n101) );
  OR2X1 U2106 ( .A(n115), .B(n112), .Y(n111) );
  OR2X1 U2111 ( .A(n125), .B(n122), .Y(n121) );
  OR2X1 U2116 ( .A(n135), .B(n132), .Y(n131) );
  OR2X1 U2123 ( .A(n145), .B(n142), .Y(n141) );
  OR2X1 U2128 ( .A(n155), .B(n152), .Y(n151) );
  INVX1 U2133 ( .A(n3184), .Y(n3080) );
  INVX1 U2138 ( .A(n3184), .Y(n3079) );
  INVX1 U2144 ( .A(n3180), .Y(n3177) );
  INVX1 U2149 ( .A(n1805), .Y(n3) );
  INVX1 U2154 ( .A(n1804), .Y(n4) );
  INVX1 U2159 ( .A(n1803), .Y(n5) );
  INVX1 U2166 ( .A(n1799), .Y(n8) );
  INVX1 U2171 ( .A(n1798), .Y(n9) );
  INVX1 U2176 ( .A(n1797), .Y(n10) );
  INVX1 U2181 ( .A(n1767), .Y(n13) );
  INVX1 U2187 ( .A(n1766), .Y(n14) );
  INVX1 U2192 ( .A(n1765), .Y(n15) );
  INVX1 U2197 ( .A(n1762), .Y(n18) );
  INVX1 U2202 ( .A(n1761), .Y(n19) );
  INVX1 U2208 ( .A(n1760), .Y(n20) );
  INVX1 U2210 ( .A(n1730), .Y(n23) );
  INVX1 U2212 ( .A(n1729), .Y(n24) );
  INVX1 U2213 ( .A(n1728), .Y(n25) );
  INVX1 U2215 ( .A(n1725), .Y(n28) );
  INVX1 U2216 ( .A(n1724), .Y(n29) );
  INVX1 U2218 ( .A(n1723), .Y(n30) );
  INVX1 U2219 ( .A(n1705), .Y(n33) );
  INVX1 U2221 ( .A(n1704), .Y(n34) );
  INVX1 U2222 ( .A(n1703), .Y(n35) );
  INVX1 U2223 ( .A(n1700), .Y(n38) );
  INVX1 U2225 ( .A(n1699), .Y(n39) );
  INVX1 U2226 ( .A(n1698), .Y(n40) );
  INVX1 U2228 ( .A(n1678), .Y(n43) );
  INVX1 U2229 ( .A(n1677), .Y(n44) );
  INVX1 U2231 ( .A(n1676), .Y(n45) );
  INVX1 U2232 ( .A(n1673), .Y(n48) );
  INVX1 U2234 ( .A(n1672), .Y(n49) );
  INVX1 U2236 ( .A(n1671), .Y(n50) );
  INVX1 U2237 ( .A(n1653), .Y(n53) );
  INVX1 U2238 ( .A(n1652), .Y(n54) );
  INVX1 U2240 ( .A(n1651), .Y(n55) );
  INVX1 U2241 ( .A(n1648), .Y(n58) );
  INVX1 U2243 ( .A(n1647), .Y(n59) );
  INVX1 U2244 ( .A(n1646), .Y(n60) );
  INVX1 U2246 ( .A(n1626), .Y(n63) );
  INVX1 U2247 ( .A(n1625), .Y(n64) );
  INVX1 U2249 ( .A(n1624), .Y(n65) );
  INVX1 U2250 ( .A(n1621), .Y(n68) );
  INVX1 U2251 ( .A(n1620), .Y(n69) );
  INVX1 U2253 ( .A(n1619), .Y(n70) );
  INVX1 U2254 ( .A(n1601), .Y(n73) );
  INVX1 U2256 ( .A(n1600), .Y(n74) );
  INVX1 U2257 ( .A(n1599), .Y(n75) );
  INVX1 U2259 ( .A(n1596), .Y(n78) );
  INVX1 U2260 ( .A(n1595), .Y(n79) );
  INVX1 U2262 ( .A(n1594), .Y(n80) );
  INVX1 U2264 ( .A(n1574), .Y(n83) );
  INVX1 U2265 ( .A(n1573), .Y(n84) );
  INVX1 U2267 ( .A(n1572), .Y(n85) );
  INVX1 U2269 ( .A(n1569), .Y(n88) );
  INVX1 U2271 ( .A(n1568), .Y(n89) );
  INVX1 U2272 ( .A(n1567), .Y(n90) );
  INVX1 U2274 ( .A(n1549), .Y(n93) );
  INVX1 U2275 ( .A(n1548), .Y(n94) );
  INVX1 U2277 ( .A(n1547), .Y(n95) );
  INVX1 U2278 ( .A(n1544), .Y(n98) );
  INVX1 U2286 ( .A(n1543), .Y(n99) );
  INVX1 U2287 ( .A(n1542), .Y(n100) );
  INVX1 U2289 ( .A(n1522), .Y(n103) );
  INVX1 U2290 ( .A(n1521), .Y(n104) );
  INVX1 U2292 ( .A(n1520), .Y(n105) );
  INVX1 U2293 ( .A(n1517), .Y(n108) );
  INVX1 U2295 ( .A(n1516), .Y(n109) );
  INVX1 U2296 ( .A(n1515), .Y(n110) );
  INVX1 U2298 ( .A(n1497), .Y(n113) );
  INVX1 U2299 ( .A(n1496), .Y(n114) );
  INVX1 U2300 ( .A(n1495), .Y(n115) );
  INVX1 U2301 ( .A(n1492), .Y(n118) );
  INVX1 U2303 ( .A(n1491), .Y(n119) );
  INVX1 U2304 ( .A(n1490), .Y(n120) );
  INVX1 U2306 ( .A(n1470), .Y(n123) );
  INVX1 U2307 ( .A(n1469), .Y(n124) );
  INVX1 U2309 ( .A(n1468), .Y(n125) );
  INVX1 U2310 ( .A(n1465), .Y(n128) );
  INVX1 U2312 ( .A(n1464), .Y(n129) );
  INVX1 U2313 ( .A(n1463), .Y(n130) );
  INVX1 U2314 ( .A(n1445), .Y(n133) );
  INVX1 U2315 ( .A(n1444), .Y(n134) );
  INVX1 U2316 ( .A(n1443), .Y(n135) );
  INVX1 U2318 ( .A(n1440), .Y(n138) );
  INVX1 U2320 ( .A(n1439), .Y(n139) );
  INVX1 U2323 ( .A(n1438), .Y(n140) );
  INVX1 U2325 ( .A(n1418), .Y(n143) );
  INVX1 U2328 ( .A(n1417), .Y(n144) );
  INVX1 U2330 ( .A(n1416), .Y(n145) );
  INVX1 U2333 ( .A(n1413), .Y(n148) );
  INVX1 U2337 ( .A(n1412), .Y(n149) );
  INVX1 U2345 ( .A(n1411), .Y(n150) );
  INVX1 U2346 ( .A(n1392), .Y(n153) );
  INVX1 U2347 ( .A(n1391), .Y(n154) );
  INVX1 U2348 ( .A(n1390), .Y(n155) );
  INVX1 U2349 ( .A(n1387), .Y(n158) );
  INVX1 U2350 ( .A(n1386), .Y(n159) );
  INVX1 U2351 ( .A(n1385), .Y(n160) );
  INVX1 U2352 ( .A(n161), .Y(n162) );
  INVX1 U2353 ( .A(n163), .Y(n164) );
  OR2X1 U2354 ( .A(N182), .B(N181), .Y(n189) );
  INVX1 U2355 ( .A(n3178), .Y(n3175) );
  INVX1 U2356 ( .A(n3179), .Y(n3176) );
  INVX1 U2357 ( .A(rst), .Y(n3186) );
  OR2X1 U2358 ( .A(n189), .B(N180), .Y(n191) );
  OR2X1 U2359 ( .A(n2354), .B(n2355), .Y(n192) );
  OR2X1 U2360 ( .A(n2357), .B(n2358), .Y(n193) );
  OR2X1 U2361 ( .A(n2360), .B(n2361), .Y(n194) );
  OR2X1 U2362 ( .A(n2363), .B(n2364), .Y(n195) );
  OR2X1 U2363 ( .A(n2366), .B(n2367), .Y(n196) );
  OR2X1 U2364 ( .A(n2369), .B(n2370), .Y(n197) );
  OR2X1 U2365 ( .A(n2372), .B(n2373), .Y(n198) );
  OR2X1 U2366 ( .A(n2375), .B(n2376), .Y(n199) );
  OR2X1 U2367 ( .A(n2378), .B(n2379), .Y(n200) );
  OR2X1 U2368 ( .A(n2381), .B(n2382), .Y(n201) );
  OR2X1 U2369 ( .A(n2384), .B(n2385), .Y(n202) );
  OR2X1 U2370 ( .A(n2387), .B(n2388), .Y(n203) );
  OR2X1 U2371 ( .A(n2390), .B(n2391), .Y(n204) );
  OR2X1 U2372 ( .A(n2393), .B(n2394), .Y(n205) );
  OR2X1 U2373 ( .A(n2396), .B(n2397), .Y(n206) );
  OR2X1 U2374 ( .A(n2399), .B(n2400), .Y(n207) );
  OR2X1 U2375 ( .A(n2404), .B(n209), .Y(n208) );
  OR2X1 U2376 ( .A(n2402), .B(n2403), .Y(n209) );
  OR2X1 U2377 ( .A(n2405), .B(n2406), .Y(n210) );
  OR2X1 U2378 ( .A(n2410), .B(n212), .Y(n211) );
  OR2X1 U2379 ( .A(n2408), .B(n2409), .Y(n212) );
  OR2X1 U2380 ( .A(n2411), .B(n2412), .Y(n213) );
  OR2X1 U2381 ( .A(n2416), .B(n215), .Y(n214) );
  OR2X1 U2382 ( .A(n2414), .B(n2415), .Y(n215) );
  OR2X1 U2383 ( .A(n2417), .B(n2418), .Y(n216) );
  OR2X1 U2384 ( .A(n2422), .B(n218), .Y(n217) );
  OR2X1 U2385 ( .A(n2420), .B(n2421), .Y(n218) );
  OR2X1 U2386 ( .A(n2423), .B(n2424), .Y(n219) );
  OR2X1 U2387 ( .A(n2428), .B(n221), .Y(n220) );
  OR2X1 U2388 ( .A(n2426), .B(n2427), .Y(n221) );
  OR2X1 U2389 ( .A(n2429), .B(n2430), .Y(n222) );
  OR2X1 U2390 ( .A(n2434), .B(n224), .Y(n223) );
  OR2X1 U2391 ( .A(n2432), .B(n2433), .Y(n224) );
  OR2X1 U2392 ( .A(n2435), .B(n2436), .Y(n225) );
  OR2X1 U2393 ( .A(n2440), .B(n227), .Y(n226) );
  OR2X1 U2394 ( .A(n2438), .B(n2439), .Y(n227) );
  OR2X1 U2395 ( .A(n2441), .B(n2442), .Y(n228) );
  OR2X1 U2396 ( .A(n2446), .B(n230), .Y(n229) );
  OR2X1 U2397 ( .A(n2444), .B(n2445), .Y(n230) );
  OR2X1 U2398 ( .A(n2447), .B(n2448), .Y(n231) );
  BUFX2 U2399 ( .A(n1356), .Y(n232) );
  BUFX2 U2400 ( .A(n1355), .Y(n233) );
  BUFX2 U2401 ( .A(n1354), .Y(n234) );
  BUFX2 U2402 ( .A(n1353), .Y(n235) );
  BUFX2 U2403 ( .A(n1352), .Y(n236) );
  BUFX2 U2404 ( .A(n1351), .Y(n237) );
  BUFX2 U2405 ( .A(n1350), .Y(n238) );
  BUFX2 U2406 ( .A(n1347), .Y(n239) );
  BUFX2 U2407 ( .A(n1344), .Y(n240) );
  BUFX2 U2408 ( .A(n1343), .Y(n241) );
  BUFX2 U2409 ( .A(n1342), .Y(n242) );
  BUFX2 U2410 ( .A(n1341), .Y(n243) );
  BUFX2 U2411 ( .A(n1340), .Y(n244) );
  BUFX2 U2412 ( .A(n1339), .Y(n245) );
  BUFX2 U2413 ( .A(n1338), .Y(n246) );
  BUFX2 U2414 ( .A(n1335), .Y(n247) );
  BUFX2 U2415 ( .A(n1332), .Y(n248) );
  BUFX2 U2416 ( .A(n1331), .Y(n249) );
  BUFX2 U2417 ( .A(n1330), .Y(n250) );
  BUFX2 U2418 ( .A(n1329), .Y(n251) );
  BUFX2 U2419 ( .A(n1328), .Y(n252) );
  BUFX2 U2420 ( .A(n1327), .Y(n253) );
  BUFX2 U2421 ( .A(n1326), .Y(n254) );
  BUFX2 U2422 ( .A(n1323), .Y(n255) );
  BUFX2 U2423 ( .A(n1320), .Y(n256) );
  BUFX2 U2424 ( .A(n1319), .Y(n257) );
  BUFX2 U2425 ( .A(n1318), .Y(n258) );
  BUFX2 U2426 ( .A(n1317), .Y(n259) );
  BUFX2 U2427 ( .A(n1316), .Y(n260) );
  BUFX2 U2428 ( .A(n1315), .Y(n261) );
  BUFX2 U2429 ( .A(n1314), .Y(n262) );
  BUFX2 U2430 ( .A(n1311), .Y(n263) );
  BUFX2 U2431 ( .A(n1308), .Y(n264) );
  BUFX2 U2432 ( .A(n1307), .Y(n265) );
  BUFX2 U2433 ( .A(n1306), .Y(n266) );
  BUFX2 U2434 ( .A(n1305), .Y(n267) );
  BUFX2 U2435 ( .A(n1304), .Y(n268) );
  BUFX2 U2436 ( .A(n1303), .Y(n269) );
  BUFX2 U2437 ( .A(n1302), .Y(n270) );
  BUFX2 U2438 ( .A(n1299), .Y(n271) );
  BUFX2 U2439 ( .A(n1296), .Y(n272) );
  BUFX2 U2440 ( .A(n1295), .Y(n273) );
  BUFX2 U2441 ( .A(n1294), .Y(n274) );
  BUFX2 U2442 ( .A(n1293), .Y(n275) );
  BUFX2 U2443 ( .A(n1292), .Y(n276) );
  BUFX2 U2444 ( .A(n1291), .Y(n277) );
  BUFX2 U2445 ( .A(n1290), .Y(n278) );
  BUFX2 U2446 ( .A(n1287), .Y(n279) );
  BUFX2 U2447 ( .A(n1284), .Y(n280) );
  BUFX2 U2448 ( .A(n1283), .Y(n281) );
  BUFX2 U2449 ( .A(n1282), .Y(n282) );
  BUFX2 U2450 ( .A(n1281), .Y(n283) );
  BUFX2 U2451 ( .A(n1280), .Y(n284) );
  BUFX2 U2452 ( .A(n1279), .Y(n285) );
  BUFX2 U2453 ( .A(n1278), .Y(n286) );
  BUFX2 U2454 ( .A(n1275), .Y(n287) );
  BUFX2 U2455 ( .A(n1272), .Y(n288) );
  BUFX2 U2456 ( .A(n1271), .Y(n289) );
  BUFX2 U2457 ( .A(n1270), .Y(n290) );
  BUFX2 U2458 ( .A(n1269), .Y(n291) );
  BUFX2 U2459 ( .A(n1268), .Y(n292) );
  BUFX2 U2460 ( .A(n1267), .Y(n293) );
  BUFX2 U2461 ( .A(n1266), .Y(n294) );
  BUFX2 U2462 ( .A(n1263), .Y(n295) );
  BUFX2 U2463 ( .A(n1260), .Y(n296) );
  BUFX2 U2464 ( .A(n1259), .Y(n297) );
  BUFX2 U2465 ( .A(n1258), .Y(n298) );
  BUFX2 U2466 ( .A(n1257), .Y(n299) );
  BUFX2 U2467 ( .A(n1256), .Y(n300) );
  BUFX2 U2468 ( .A(n1255), .Y(n301) );
  BUFX2 U2469 ( .A(n1254), .Y(n302) );
  BUFX2 U2470 ( .A(n1251), .Y(n303) );
  BUFX2 U2471 ( .A(n1248), .Y(n304) );
  BUFX2 U2472 ( .A(n1247), .Y(n305) );
  BUFX2 U2473 ( .A(n1246), .Y(n306) );
  BUFX2 U2474 ( .A(n1245), .Y(n307) );
  BUFX2 U2475 ( .A(n1244), .Y(n308) );
  BUFX2 U2476 ( .A(n1243), .Y(n309) );
  BUFX2 U2477 ( .A(n1242), .Y(n310) );
  BUFX2 U2478 ( .A(n1239), .Y(n311) );
  BUFX2 U2479 ( .A(n1236), .Y(n312) );
  BUFX2 U2480 ( .A(n1235), .Y(n313) );
  BUFX2 U2481 ( .A(n1234), .Y(n314) );
  BUFX2 U2482 ( .A(n1233), .Y(n315) );
  BUFX2 U2483 ( .A(n1232), .Y(n316) );
  BUFX2 U2484 ( .A(n1231), .Y(n317) );
  BUFX2 U2485 ( .A(n1230), .Y(n318) );
  BUFX2 U2486 ( .A(n1227), .Y(n319) );
  BUFX2 U2487 ( .A(n1224), .Y(n320) );
  BUFX2 U2488 ( .A(n1223), .Y(n321) );
  BUFX2 U2489 ( .A(n1222), .Y(n322) );
  BUFX2 U2490 ( .A(n1221), .Y(n323) );
  BUFX2 U2491 ( .A(n1220), .Y(n324) );
  BUFX2 U2492 ( .A(n1219), .Y(n325) );
  BUFX2 U2493 ( .A(n1218), .Y(n326) );
  BUFX2 U2494 ( .A(n1215), .Y(n327) );
  BUFX2 U2495 ( .A(n1212), .Y(n328) );
  BUFX2 U2496 ( .A(n1211), .Y(n329) );
  BUFX2 U2497 ( .A(n1210), .Y(n330) );
  BUFX2 U2498 ( .A(n1209), .Y(n331) );
  BUFX2 U2499 ( .A(n1208), .Y(n332) );
  BUFX2 U2500 ( .A(n1207), .Y(n333) );
  BUFX2 U2501 ( .A(n1206), .Y(n334) );
  BUFX2 U2502 ( .A(n1203), .Y(n335) );
  BUFX2 U2503 ( .A(n1200), .Y(n336) );
  BUFX2 U2504 ( .A(n1199), .Y(n337) );
  BUFX2 U2505 ( .A(n1198), .Y(n338) );
  BUFX2 U2506 ( .A(n1197), .Y(n339) );
  BUFX2 U2507 ( .A(n1196), .Y(n340) );
  BUFX2 U2508 ( .A(n1195), .Y(n341) );
  BUFX2 U2509 ( .A(n1194), .Y(n342) );
  BUFX2 U2510 ( .A(n1191), .Y(n343) );
  BUFX2 U2511 ( .A(n1188), .Y(n344) );
  BUFX2 U2512 ( .A(n1187), .Y(n345) );
  BUFX2 U2513 ( .A(n1186), .Y(n346) );
  BUFX2 U2514 ( .A(n1185), .Y(n347) );
  BUFX2 U2515 ( .A(n1184), .Y(n348) );
  BUFX2 U2516 ( .A(n1183), .Y(n349) );
  BUFX2 U2517 ( .A(n1182), .Y(n350) );
  BUFX2 U2518 ( .A(n1179), .Y(n351) );
  BUFX2 U2519 ( .A(n1176), .Y(n352) );
  BUFX2 U2520 ( .A(n1175), .Y(n353) );
  BUFX2 U2521 ( .A(n1174), .Y(n354) );
  BUFX2 U2522 ( .A(n1173), .Y(n355) );
  BUFX2 U2523 ( .A(n1172), .Y(n356) );
  BUFX2 U2524 ( .A(n1171), .Y(n357) );
  BUFX2 U2525 ( .A(n1170), .Y(n358) );
  BUFX2 U2526 ( .A(n1167), .Y(n359) );
  BUFX2 U2527 ( .A(n1164), .Y(n360) );
  BUFX2 U2528 ( .A(n1163), .Y(n361) );
  BUFX2 U2529 ( .A(n1162), .Y(n362) );
  BUFX2 U2530 ( .A(n1161), .Y(n363) );
  BUFX2 U2531 ( .A(n1160), .Y(n364) );
  BUFX2 U2532 ( .A(n1159), .Y(n365) );
  BUFX2 U2533 ( .A(n1158), .Y(n366) );
  BUFX2 U2534 ( .A(n1155), .Y(n367) );
  BUFX2 U2535 ( .A(n1152), .Y(n368) );
  BUFX2 U2536 ( .A(n1151), .Y(n369) );
  BUFX2 U2537 ( .A(n1150), .Y(n370) );
  BUFX2 U2538 ( .A(n1149), .Y(n371) );
  BUFX2 U2539 ( .A(n1148), .Y(n372) );
  BUFX2 U2540 ( .A(n1147), .Y(n373) );
  BUFX2 U2541 ( .A(n1146), .Y(n374) );
  BUFX2 U2542 ( .A(n1143), .Y(n375) );
  BUFX2 U2543 ( .A(n1140), .Y(n376) );
  BUFX2 U2544 ( .A(n1139), .Y(n377) );
  BUFX2 U2545 ( .A(n1138), .Y(n378) );
  BUFX2 U2546 ( .A(n1137), .Y(n379) );
  BUFX2 U2547 ( .A(n1136), .Y(n380) );
  BUFX2 U2548 ( .A(n1135), .Y(n381) );
  BUFX2 U2549 ( .A(n1134), .Y(n382) );
  BUFX2 U2550 ( .A(n1131), .Y(n383) );
  BUFX2 U2551 ( .A(n1128), .Y(n384) );
  BUFX2 U2552 ( .A(n1127), .Y(n385) );
  BUFX2 U2553 ( .A(n1126), .Y(n386) );
  BUFX2 U2554 ( .A(n1125), .Y(n387) );
  BUFX2 U2555 ( .A(n1124), .Y(n388) );
  BUFX2 U2556 ( .A(n1123), .Y(n389) );
  BUFX2 U2557 ( .A(n1122), .Y(n390) );
  BUFX2 U2558 ( .A(n1119), .Y(n391) );
  BUFX2 U2559 ( .A(n1116), .Y(n392) );
  BUFX2 U2560 ( .A(n1115), .Y(n393) );
  BUFX2 U2561 ( .A(n1114), .Y(n394) );
  BUFX2 U2562 ( .A(n1113), .Y(n395) );
  BUFX2 U2563 ( .A(n1112), .Y(n396) );
  BUFX2 U2564 ( .A(n1111), .Y(n397) );
  BUFX2 U2565 ( .A(n1110), .Y(n398) );
  BUFX2 U2566 ( .A(n1107), .Y(n399) );
  BUFX2 U2567 ( .A(n1104), .Y(n400) );
  BUFX2 U2568 ( .A(n1103), .Y(n401) );
  BUFX2 U2569 ( .A(n1102), .Y(n402) );
  BUFX2 U2570 ( .A(n1101), .Y(n403) );
  BUFX2 U2571 ( .A(n1100), .Y(n404) );
  BUFX2 U2572 ( .A(n1099), .Y(n405) );
  BUFX2 U2573 ( .A(n1098), .Y(n406) );
  BUFX2 U2574 ( .A(n1095), .Y(n407) );
  BUFX2 U2575 ( .A(n1092), .Y(n408) );
  BUFX2 U2576 ( .A(n1091), .Y(n409) );
  BUFX2 U2577 ( .A(n1090), .Y(n410) );
  BUFX2 U2578 ( .A(n1089), .Y(n411) );
  BUFX2 U2579 ( .A(n1088), .Y(n412) );
  BUFX2 U2580 ( .A(n1087), .Y(n413) );
  BUFX2 U2581 ( .A(n1086), .Y(n414) );
  BUFX2 U2582 ( .A(n1083), .Y(n415) );
  BUFX2 U2583 ( .A(n1080), .Y(n416) );
  BUFX2 U2584 ( .A(n1079), .Y(n417) );
  BUFX2 U2585 ( .A(n1078), .Y(n418) );
  BUFX2 U2586 ( .A(n1077), .Y(n419) );
  BUFX2 U2587 ( .A(n1076), .Y(n420) );
  BUFX2 U2588 ( .A(n1075), .Y(n421) );
  BUFX2 U2589 ( .A(n1074), .Y(n422) );
  BUFX2 U2590 ( .A(n1071), .Y(n423) );
  BUFX2 U2591 ( .A(n1068), .Y(n424) );
  BUFX2 U2592 ( .A(n1067), .Y(n425) );
  BUFX2 U2593 ( .A(n1066), .Y(n426) );
  BUFX2 U2594 ( .A(n1065), .Y(n427) );
  BUFX2 U2595 ( .A(n1064), .Y(n428) );
  BUFX2 U2596 ( .A(n1063), .Y(n429) );
  BUFX2 U2597 ( .A(n1062), .Y(n430) );
  BUFX2 U2598 ( .A(n1059), .Y(n431) );
  BUFX2 U2599 ( .A(n1056), .Y(n432) );
  BUFX2 U2600 ( .A(n1055), .Y(n433) );
  BUFX2 U2601 ( .A(n1054), .Y(n434) );
  BUFX2 U2602 ( .A(n1053), .Y(n435) );
  BUFX2 U2603 ( .A(n1052), .Y(n436) );
  BUFX2 U2604 ( .A(n1051), .Y(n437) );
  BUFX2 U2605 ( .A(n1050), .Y(n438) );
  BUFX2 U2606 ( .A(n1047), .Y(n439) );
  BUFX2 U2607 ( .A(n1044), .Y(n440) );
  BUFX2 U2608 ( .A(n1043), .Y(n441) );
  BUFX2 U2609 ( .A(n1042), .Y(n442) );
  BUFX2 U2610 ( .A(n1041), .Y(n443) );
  BUFX2 U2611 ( .A(n1040), .Y(n444) );
  BUFX2 U2612 ( .A(n1039), .Y(n445) );
  BUFX2 U2613 ( .A(n1038), .Y(n446) );
  BUFX2 U2614 ( .A(n1035), .Y(n447) );
  BUFX2 U2615 ( .A(n1032), .Y(n448) );
  BUFX2 U2616 ( .A(n1031), .Y(n449) );
  BUFX2 U2617 ( .A(n1030), .Y(n450) );
  BUFX2 U2618 ( .A(n1029), .Y(n451) );
  BUFX2 U2619 ( .A(n1028), .Y(n452) );
  BUFX2 U2620 ( .A(n1027), .Y(n453) );
  BUFX2 U2621 ( .A(n1026), .Y(n454) );
  BUFX2 U2622 ( .A(n1023), .Y(n455) );
  BUFX2 U2623 ( .A(n1020), .Y(n456) );
  BUFX2 U2624 ( .A(n1019), .Y(n457) );
  BUFX2 U2625 ( .A(n1018), .Y(n458) );
  BUFX2 U2626 ( .A(n1017), .Y(n459) );
  BUFX2 U2627 ( .A(n1016), .Y(n460) );
  BUFX2 U2628 ( .A(n1015), .Y(n461) );
  BUFX2 U2629 ( .A(n1014), .Y(n462) );
  BUFX2 U2630 ( .A(n1011), .Y(n463) );
  BUFX2 U2631 ( .A(n1008), .Y(n464) );
  BUFX2 U2632 ( .A(n1007), .Y(n465) );
  BUFX2 U2633 ( .A(n1006), .Y(n466) );
  BUFX2 U2634 ( .A(n1005), .Y(n467) );
  BUFX2 U2635 ( .A(n1004), .Y(n468) );
  BUFX2 U2636 ( .A(n1003), .Y(n469) );
  BUFX2 U2637 ( .A(n1002), .Y(n470) );
  BUFX2 U2638 ( .A(n999), .Y(n471) );
  BUFX2 U2639 ( .A(n996), .Y(n472) );
  BUFX2 U2640 ( .A(n995), .Y(n473) );
  BUFX2 U2641 ( .A(n994), .Y(n474) );
  BUFX2 U2642 ( .A(n993), .Y(n475) );
  BUFX2 U2643 ( .A(n992), .Y(n476) );
  BUFX2 U2644 ( .A(n991), .Y(n477) );
  BUFX2 U2645 ( .A(n990), .Y(n478) );
  BUFX2 U2646 ( .A(n987), .Y(n479) );
  BUFX2 U2647 ( .A(n984), .Y(n480) );
  BUFX2 U2648 ( .A(n983), .Y(n481) );
  BUFX2 U2649 ( .A(n982), .Y(n482) );
  BUFX2 U2650 ( .A(n981), .Y(n483) );
  BUFX2 U2651 ( .A(n980), .Y(n484) );
  BUFX2 U2652 ( .A(n979), .Y(n485) );
  BUFX2 U2653 ( .A(n978), .Y(n486) );
  BUFX2 U2654 ( .A(n975), .Y(n487) );
  BUFX2 U2655 ( .A(n972), .Y(n488) );
  BUFX2 U2656 ( .A(n971), .Y(n489) );
  BUFX2 U2657 ( .A(n970), .Y(n490) );
  BUFX2 U2658 ( .A(n969), .Y(n491) );
  BUFX2 U2659 ( .A(n968), .Y(n492) );
  BUFX2 U2660 ( .A(n967), .Y(n493) );
  BUFX2 U2661 ( .A(n966), .Y(n494) );
  BUFX2 U2662 ( .A(n963), .Y(n495) );
  BUFX2 U2663 ( .A(n960), .Y(n496) );
  BUFX2 U2664 ( .A(n959), .Y(n497) );
  BUFX2 U2665 ( .A(n958), .Y(n498) );
  BUFX2 U2666 ( .A(n957), .Y(n499) );
  BUFX2 U2667 ( .A(n956), .Y(n500) );
  BUFX2 U2668 ( .A(n955), .Y(n501) );
  BUFX2 U2669 ( .A(n954), .Y(n502) );
  BUFX2 U2670 ( .A(n951), .Y(n503) );
  BUFX2 U2671 ( .A(n948), .Y(n504) );
  BUFX2 U2672 ( .A(n947), .Y(n505) );
  BUFX2 U2673 ( .A(n946), .Y(n506) );
  BUFX2 U2674 ( .A(n945), .Y(n507) );
  BUFX2 U2675 ( .A(n944), .Y(n508) );
  BUFX2 U2676 ( .A(n943), .Y(n509) );
  BUFX2 U2677 ( .A(n942), .Y(n510) );
  BUFX2 U2678 ( .A(n939), .Y(n511) );
  BUFX2 U2679 ( .A(n936), .Y(n512) );
  BUFX2 U2680 ( .A(n935), .Y(n513) );
  BUFX2 U2681 ( .A(n934), .Y(n514) );
  BUFX2 U2682 ( .A(n933), .Y(n515) );
  BUFX2 U2683 ( .A(n932), .Y(n516) );
  BUFX2 U2684 ( .A(n931), .Y(n517) );
  BUFX2 U2685 ( .A(n930), .Y(n518) );
  BUFX2 U2686 ( .A(n927), .Y(n519) );
  BUFX2 U2687 ( .A(n924), .Y(n520) );
  BUFX2 U2688 ( .A(n923), .Y(n521) );
  BUFX2 U2689 ( .A(n922), .Y(n522) );
  BUFX2 U2690 ( .A(n921), .Y(n523) );
  BUFX2 U2691 ( .A(n920), .Y(n524) );
  BUFX2 U2692 ( .A(n919), .Y(n525) );
  BUFX2 U2693 ( .A(n918), .Y(n526) );
  BUFX2 U2694 ( .A(n915), .Y(n527) );
  BUFX2 U2695 ( .A(n912), .Y(n528) );
  BUFX2 U2696 ( .A(n911), .Y(n529) );
  BUFX2 U2697 ( .A(n910), .Y(n530) );
  BUFX2 U2698 ( .A(n909), .Y(n531) );
  BUFX2 U2699 ( .A(n908), .Y(n532) );
  BUFX2 U2700 ( .A(n907), .Y(n533) );
  BUFX2 U2701 ( .A(n906), .Y(n534) );
  BUFX2 U2702 ( .A(n903), .Y(n535) );
  BUFX2 U2703 ( .A(n900), .Y(n536) );
  BUFX2 U2704 ( .A(n899), .Y(n537) );
  BUFX2 U2705 ( .A(n898), .Y(n538) );
  BUFX2 U2706 ( .A(n897), .Y(n539) );
  BUFX2 U2707 ( .A(n896), .Y(n540) );
  BUFX2 U2708 ( .A(n895), .Y(n541) );
  BUFX2 U2709 ( .A(n894), .Y(n542) );
  BUFX2 U2710 ( .A(n891), .Y(n543) );
  BUFX2 U2711 ( .A(n888), .Y(n544) );
  BUFX2 U2712 ( .A(n887), .Y(n545) );
  BUFX2 U2713 ( .A(n886), .Y(n546) );
  BUFX2 U2714 ( .A(n885), .Y(n547) );
  BUFX2 U2715 ( .A(n884), .Y(n548) );
  BUFX2 U2716 ( .A(n883), .Y(n549) );
  BUFX2 U2717 ( .A(n882), .Y(n550) );
  BUFX2 U2718 ( .A(n879), .Y(n551) );
  BUFX2 U2719 ( .A(n876), .Y(n552) );
  BUFX2 U2720 ( .A(n875), .Y(n553) );
  BUFX2 U2721 ( .A(n874), .Y(n554) );
  BUFX2 U2722 ( .A(n873), .Y(n555) );
  BUFX2 U2723 ( .A(n872), .Y(n556) );
  BUFX2 U2724 ( .A(n871), .Y(n557) );
  BUFX2 U2725 ( .A(n870), .Y(n558) );
  BUFX2 U2726 ( .A(n867), .Y(n559) );
  BUFX2 U2727 ( .A(n864), .Y(n560) );
  BUFX2 U2728 ( .A(n863), .Y(n561) );
  BUFX2 U2729 ( .A(n862), .Y(n562) );
  BUFX2 U2730 ( .A(n861), .Y(n563) );
  BUFX2 U2731 ( .A(n860), .Y(n564) );
  BUFX2 U2732 ( .A(n859), .Y(n565) );
  BUFX2 U2733 ( .A(n858), .Y(n566) );
  BUFX2 U2734 ( .A(n855), .Y(n567) );
  BUFX2 U2735 ( .A(n852), .Y(n568) );
  BUFX2 U2736 ( .A(n851), .Y(n569) );
  BUFX2 U2737 ( .A(n850), .Y(n570) );
  BUFX2 U2738 ( .A(n849), .Y(n571) );
  BUFX2 U2739 ( .A(n848), .Y(n572) );
  BUFX2 U2740 ( .A(n847), .Y(n573) );
  BUFX2 U2741 ( .A(n846), .Y(n574) );
  BUFX2 U2742 ( .A(n843), .Y(n575) );
  BUFX2 U2743 ( .A(n840), .Y(n576) );
  BUFX2 U2744 ( .A(n839), .Y(n577) );
  BUFX2 U2745 ( .A(n838), .Y(n578) );
  BUFX2 U2746 ( .A(n837), .Y(n579) );
  BUFX2 U2747 ( .A(n836), .Y(n580) );
  BUFX2 U2748 ( .A(n835), .Y(n581) );
  BUFX2 U2749 ( .A(n834), .Y(n582) );
  BUFX2 U2750 ( .A(n831), .Y(n583) );
  BUFX2 U2751 ( .A(n828), .Y(n584) );
  BUFX2 U2752 ( .A(n827), .Y(n585) );
  BUFX2 U2753 ( .A(n826), .Y(n586) );
  BUFX2 U2754 ( .A(n825), .Y(n587) );
  BUFX2 U2755 ( .A(n824), .Y(n588) );
  BUFX2 U2756 ( .A(n823), .Y(n589) );
  BUFX2 U2757 ( .A(n822), .Y(n590) );
  BUFX2 U2758 ( .A(n819), .Y(n591) );
  BUFX2 U2759 ( .A(n816), .Y(n592) );
  BUFX2 U2760 ( .A(n815), .Y(n593) );
  BUFX2 U2761 ( .A(n814), .Y(n594) );
  BUFX2 U2762 ( .A(n813), .Y(n595) );
  BUFX2 U2763 ( .A(n812), .Y(n596) );
  BUFX2 U2764 ( .A(n811), .Y(n597) );
  BUFX2 U2765 ( .A(n810), .Y(n609) );
  BUFX2 U2766 ( .A(n807), .Y(n611) );
  BUFX2 U2767 ( .A(n804), .Y(n624) );
  BUFX2 U2768 ( .A(n803), .Y(n637) );
  BUFX2 U2769 ( .A(n802), .Y(n649) );
  BUFX2 U2770 ( .A(n801), .Y(n661) );
  BUFX2 U2771 ( .A(n800), .Y(n673) );
  BUFX2 U2772 ( .A(n799), .Y(n685) );
  BUFX2 U2773 ( .A(n798), .Y(n697) );
  BUFX2 U2774 ( .A(n795), .Y(n709) );
  BUFX2 U2775 ( .A(n792), .Y(n721) );
  BUFX2 U2776 ( .A(n791), .Y(n733) );
  BUFX2 U2777 ( .A(n790), .Y(n745) );
  BUFX2 U2778 ( .A(n789), .Y(n757) );
  BUFX2 U2779 ( .A(n788), .Y(n769) );
  BUFX2 U2780 ( .A(n787), .Y(n781) );
  BUFX2 U2781 ( .A(n786), .Y(n793) );
  BUFX2 U2782 ( .A(n783), .Y(n805) );
  BUFX2 U2783 ( .A(n780), .Y(n817) );
  BUFX2 U2784 ( .A(n779), .Y(n829) );
  BUFX2 U2785 ( .A(n778), .Y(n841) );
  BUFX2 U2786 ( .A(n777), .Y(n853) );
  BUFX2 U2787 ( .A(n776), .Y(n865) );
  BUFX2 U2788 ( .A(n775), .Y(n877) );
  BUFX2 U2789 ( .A(n774), .Y(n889) );
  BUFX2 U2790 ( .A(n771), .Y(n901) );
  BUFX2 U2791 ( .A(n768), .Y(n913) );
  BUFX2 U2792 ( .A(n767), .Y(n925) );
  BUFX2 U2793 ( .A(n766), .Y(n937) );
  BUFX2 U2794 ( .A(n765), .Y(n949) );
  BUFX2 U2795 ( .A(n764), .Y(n961) );
  BUFX2 U2796 ( .A(n763), .Y(n973) );
  BUFX2 U2797 ( .A(n762), .Y(n985) );
  BUFX2 U2798 ( .A(n759), .Y(n997) );
  BUFX2 U2799 ( .A(n756), .Y(n1009) );
  BUFX2 U2800 ( .A(n755), .Y(n1021) );
  BUFX2 U2801 ( .A(n754), .Y(n1033) );
  BUFX2 U2802 ( .A(n753), .Y(n1045) );
  BUFX2 U2803 ( .A(n752), .Y(n1057) );
  BUFX2 U2804 ( .A(n751), .Y(n1069) );
  BUFX2 U2805 ( .A(n750), .Y(n1081) );
  BUFX2 U2806 ( .A(n747), .Y(n1093) );
  BUFX2 U2807 ( .A(n744), .Y(n1105) );
  BUFX2 U2808 ( .A(n743), .Y(n1117) );
  BUFX2 U2809 ( .A(n742), .Y(n1129) );
  BUFX2 U2810 ( .A(n741), .Y(n1141) );
  BUFX2 U2811 ( .A(n740), .Y(n1153) );
  BUFX2 U2812 ( .A(n739), .Y(n1165) );
  BUFX2 U2813 ( .A(n738), .Y(n1177) );
  BUFX2 U2814 ( .A(n735), .Y(n1189) );
  BUFX2 U2815 ( .A(n732), .Y(n1201) );
  BUFX2 U2816 ( .A(n731), .Y(n1213) );
  BUFX2 U2817 ( .A(n730), .Y(n1225) );
  BUFX2 U2818 ( .A(n729), .Y(n1237) );
  BUFX2 U2819 ( .A(n728), .Y(n1249) );
  BUFX2 U2820 ( .A(n727), .Y(n1261) );
  BUFX2 U2821 ( .A(n726), .Y(n1273) );
  BUFX2 U2822 ( .A(n723), .Y(n1285) );
  BUFX2 U2823 ( .A(n720), .Y(n1297) );
  BUFX2 U2824 ( .A(n719), .Y(n1309) );
  BUFX2 U2825 ( .A(n718), .Y(n1321) );
  BUFX2 U2826 ( .A(n717), .Y(n1333) );
  BUFX2 U2827 ( .A(n716), .Y(n1345) );
  BUFX2 U2828 ( .A(n715), .Y(n1357) );
  BUFX2 U2829 ( .A(n714), .Y(n1358) );
  BUFX2 U2830 ( .A(n711), .Y(n1359) );
  BUFX2 U2831 ( .A(n708), .Y(n1360) );
  BUFX2 U2832 ( .A(n707), .Y(n1361) );
  BUFX2 U2833 ( .A(n706), .Y(n1362) );
  BUFX2 U2834 ( .A(n705), .Y(n1363) );
  BUFX2 U2835 ( .A(n704), .Y(n1364) );
  BUFX2 U2836 ( .A(n703), .Y(n1365) );
  BUFX2 U2837 ( .A(n702), .Y(n1366) );
  BUFX2 U2838 ( .A(n699), .Y(n1369) );
  BUFX2 U2839 ( .A(n696), .Y(n1371) );
  BUFX2 U2840 ( .A(n695), .Y(n1372) );
  BUFX2 U2841 ( .A(n694), .Y(n1383) );
  BUFX2 U2842 ( .A(n693), .Y(n1384) );
  BUFX2 U2843 ( .A(n692), .Y(n1396) );
  BUFX2 U2844 ( .A(n691), .Y(n1397) );
  BUFX2 U2845 ( .A(n690), .Y(n1409) );
  BUFX2 U2846 ( .A(n687), .Y(n1410) );
  BUFX2 U2847 ( .A(n684), .Y(n1424) );
  BUFX2 U2848 ( .A(n683), .Y(n1425) );
  BUFX2 U2849 ( .A(n682), .Y(n1436) );
  BUFX2 U2850 ( .A(n681), .Y(n1437) );
  BUFX2 U2851 ( .A(n680), .Y(n1449) );
  BUFX2 U2852 ( .A(n679), .Y(n1450) );
  BUFX2 U2853 ( .A(n678), .Y(n1461) );
  BUFX2 U2854 ( .A(n675), .Y(n1462) );
  BUFX2 U2855 ( .A(n672), .Y(n1476) );
  BUFX2 U2856 ( .A(n671), .Y(n1477) );
  BUFX2 U2857 ( .A(n670), .Y(n1488) );
  BUFX2 U2858 ( .A(n669), .Y(n1489) );
  BUFX2 U2859 ( .A(n668), .Y(n1501) );
  BUFX2 U2860 ( .A(n667), .Y(n1502) );
  BUFX2 U2861 ( .A(n666), .Y(n1513) );
  BUFX2 U2862 ( .A(n663), .Y(n1514) );
  BUFX2 U2863 ( .A(n660), .Y(n1528) );
  BUFX2 U2864 ( .A(n659), .Y(n1529) );
  BUFX2 U2865 ( .A(n658), .Y(n1540) );
  BUFX2 U2866 ( .A(n657), .Y(n1541) );
  BUFX2 U2867 ( .A(n656), .Y(n1553) );
  BUFX2 U2868 ( .A(n655), .Y(n1554) );
  BUFX2 U2869 ( .A(n654), .Y(n1565) );
  BUFX2 U2870 ( .A(n651), .Y(n1566) );
  BUFX2 U2871 ( .A(n648), .Y(n1580) );
  BUFX2 U2872 ( .A(n647), .Y(n1581) );
  BUFX2 U2873 ( .A(n646), .Y(n1592) );
  BUFX2 U2874 ( .A(n645), .Y(n1593) );
  BUFX2 U2875 ( .A(n644), .Y(n1605) );
  BUFX2 U2876 ( .A(n643), .Y(n1606) );
  BUFX2 U2877 ( .A(n642), .Y(n1617) );
  BUFX2 U2878 ( .A(n639), .Y(n1618) );
  BUFX2 U2879 ( .A(n636), .Y(n1632) );
  BUFX2 U2880 ( .A(n635), .Y(n1633) );
  BUFX2 U2881 ( .A(n634), .Y(n1644) );
  BUFX2 U2882 ( .A(n633), .Y(n1645) );
  BUFX2 U2883 ( .A(n632), .Y(n1657) );
  BUFX2 U2884 ( .A(n631), .Y(n1658) );
  BUFX2 U2885 ( .A(n630), .Y(n1669) );
  BUFX2 U2886 ( .A(n627), .Y(n1670) );
  BUFX2 U2887 ( .A(n623), .Y(n1684) );
  BUFX2 U2888 ( .A(n622), .Y(n1685) );
  BUFX2 U2889 ( .A(n621), .Y(n1696) );
  BUFX2 U2890 ( .A(n620), .Y(n1697) );
  BUFX2 U2891 ( .A(n619), .Y(n1709) );
  BUFX2 U2892 ( .A(n618), .Y(n1710) );
  BUFX2 U2893 ( .A(n617), .Y(n1721) );
  BUFX2 U2894 ( .A(n614), .Y(n1722) );
  BUFX2 U2895 ( .A(n608), .Y(n1736) );
  BUFX2 U2896 ( .A(n607), .Y(n1737) );
  BUFX2 U2897 ( .A(n606), .Y(n1758) );
  BUFX2 U2898 ( .A(n605), .Y(n1759) );
  BUFX2 U2899 ( .A(n604), .Y(n1771) );
  BUFX2 U2900 ( .A(n603), .Y(n1773) );
  BUFX2 U2901 ( .A(n602), .Y(n1775) );
  BUFX2 U2902 ( .A(n599), .Y(n1776) );
  AND2X1 U2903 ( .A(n2457), .B(\data_in<15> ), .Y(n1793) );
  INVX1 U2904 ( .A(n1793), .Y(n1794) );
  AND2X1 U2905 ( .A(n2457), .B(\data_in<14> ), .Y(n1795) );
  INVX1 U2906 ( .A(n1795), .Y(n1796) );
  AND2X1 U2907 ( .A(n2457), .B(\data_in<13> ), .Y(n1802) );
  INVX1 U2908 ( .A(n1802), .Y(n2328) );
  AND2X1 U2909 ( .A(n2457), .B(\data_in<12> ), .Y(n2329) );
  INVX1 U2910 ( .A(n2329), .Y(n2330) );
  AND2X1 U2911 ( .A(n2457), .B(\data_in<11> ), .Y(n2331) );
  INVX1 U2912 ( .A(n2331), .Y(n2332) );
  AND2X1 U2913 ( .A(n2457), .B(\data_in<10> ), .Y(n2333) );
  INVX1 U2914 ( .A(n2333), .Y(n2334) );
  AND2X1 U2915 ( .A(n2457), .B(\data_in<9> ), .Y(n2335) );
  INVX1 U2916 ( .A(n2335), .Y(n2336) );
  AND2X1 U2917 ( .A(n2457), .B(\data_in<8> ), .Y(n2337) );
  INVX1 U2918 ( .A(n2337), .Y(n2338) );
  BUFX2 U2919 ( .A(n1810), .Y(n2339) );
  INVX1 U2920 ( .A(n2339), .Y(n3188) );
  BUFX2 U2921 ( .A(n1808), .Y(n2340) );
  INVX1 U2922 ( .A(n2340), .Y(n3193) );
  INVX1 U2923 ( .A(n1756), .Y(n2341) );
  INVX1 U2924 ( .A(n1787), .Y(n3192) );
  INVX1 U2925 ( .A(n1772), .Y(n3189) );
  INVX1 U2926 ( .A(n1770), .Y(n3191) );
  INVX1 U2927 ( .A(n1755), .Y(n3190) );
  BUFX2 U2928 ( .A(n3716), .Y(\data_out<0> ) );
  BUFX2 U2929 ( .A(n3715), .Y(\data_out<1> ) );
  BUFX2 U2930 ( .A(n3714), .Y(\data_out<2> ) );
  BUFX2 U2931 ( .A(n3713), .Y(\data_out<3> ) );
  BUFX2 U2932 ( .A(n3712), .Y(\data_out<4> ) );
  BUFX2 U2933 ( .A(n3711), .Y(\data_out<5> ) );
  BUFX2 U2934 ( .A(n3710), .Y(\data_out<6> ) );
  BUFX2 U2935 ( .A(n3709), .Y(\data_out<7> ) );
  OR2X1 U2936 ( .A(N181), .B(n3185), .Y(n2350) );
  INVX1 U2937 ( .A(n2350), .Y(n2351) );
  OR2X1 U2938 ( .A(N181), .B(N180), .Y(n2352) );
  INVX1 U2939 ( .A(n2352), .Y(n2353) );
  INVX1 U2940 ( .A(n1790), .Y(n2354) );
  INVX1 U2941 ( .A(n1789), .Y(n2355) );
  INVX1 U2942 ( .A(n1788), .Y(n2356) );
  INVX1 U2943 ( .A(n612), .Y(n3187) );
  INVX1 U2944 ( .A(n1752), .Y(n2357) );
  INVX1 U2945 ( .A(n1751), .Y(n2358) );
  INVX1 U2946 ( .A(n1750), .Y(n2359) );
  INVX1 U2947 ( .A(n1718), .Y(n2360) );
  INVX1 U2948 ( .A(n1717), .Y(n2361) );
  INVX1 U2949 ( .A(n1716), .Y(n2362) );
  INVX1 U2950 ( .A(n1693), .Y(n2363) );
  INVX1 U2951 ( .A(n1692), .Y(n2364) );
  INVX1 U2952 ( .A(n1691), .Y(n2365) );
  INVX1 U2953 ( .A(n1666), .Y(n2366) );
  INVX1 U2954 ( .A(n1665), .Y(n2367) );
  INVX1 U2955 ( .A(n1664), .Y(n2368) );
  INVX1 U2956 ( .A(n1641), .Y(n2369) );
  INVX1 U2957 ( .A(n1640), .Y(n2370) );
  INVX1 U2958 ( .A(n1639), .Y(n2371) );
  INVX1 U2959 ( .A(n1614), .Y(n2372) );
  INVX1 U2960 ( .A(n1613), .Y(n2373) );
  INVX1 U2961 ( .A(n1612), .Y(n2374) );
  INVX1 U2962 ( .A(n1589), .Y(n2375) );
  INVX1 U2963 ( .A(n1588), .Y(n2376) );
  INVX1 U2964 ( .A(n1587), .Y(n2377) );
  INVX1 U2965 ( .A(n1562), .Y(n2378) );
  INVX1 U2966 ( .A(n1561), .Y(n2379) );
  INVX1 U2967 ( .A(n1560), .Y(n2380) );
  INVX1 U2968 ( .A(n1537), .Y(n2381) );
  INVX1 U2969 ( .A(n1536), .Y(n2382) );
  INVX1 U2970 ( .A(n1535), .Y(n2383) );
  INVX1 U2971 ( .A(n1510), .Y(n2384) );
  INVX1 U2972 ( .A(n1509), .Y(n2385) );
  INVX1 U2973 ( .A(n1508), .Y(n2386) );
  INVX1 U2974 ( .A(n1485), .Y(n2387) );
  INVX1 U2975 ( .A(n1484), .Y(n2388) );
  INVX1 U2976 ( .A(n1483), .Y(n2389) );
  INVX1 U2977 ( .A(n1458), .Y(n2390) );
  INVX1 U2978 ( .A(n1457), .Y(n2391) );
  INVX1 U2979 ( .A(n1456), .Y(n2392) );
  INVX1 U2980 ( .A(n1433), .Y(n2393) );
  INVX1 U2981 ( .A(n1432), .Y(n2394) );
  INVX1 U2982 ( .A(n1431), .Y(n2395) );
  INVX1 U2983 ( .A(n1406), .Y(n2396) );
  INVX1 U2984 ( .A(n1405), .Y(n2397) );
  INVX1 U2985 ( .A(n1404), .Y(n2398) );
  INVX1 U2986 ( .A(n1380), .Y(n2399) );
  INVX1 U2987 ( .A(n1379), .Y(n2400) );
  INVX1 U2988 ( .A(n1378), .Y(n2401) );
  INVX1 U2989 ( .A(n1779), .Y(n2402) );
  INVX1 U2990 ( .A(n1778), .Y(n2403) );
  INVX1 U2991 ( .A(n1777), .Y(n2404) );
  INVX1 U2992 ( .A(n1740), .Y(n2405) );
  INVX1 U2993 ( .A(n1739), .Y(n2406) );
  INVX1 U2994 ( .A(n1738), .Y(n2407) );
  INVX1 U2995 ( .A(n1713), .Y(n2408) );
  INVX1 U2996 ( .A(n1712), .Y(n2409) );
  INVX1 U2997 ( .A(n1711), .Y(n2410) );
  INVX1 U2998 ( .A(n1688), .Y(n2411) );
  INVX1 U2999 ( .A(n1687), .Y(n2412) );
  INVX1 U3000 ( .A(n1686), .Y(n2413) );
  INVX1 U3001 ( .A(n1661), .Y(n2414) );
  INVX1 U3002 ( .A(n1660), .Y(n2415) );
  INVX1 U3003 ( .A(n1659), .Y(n2416) );
  INVX1 U3004 ( .A(n1636), .Y(n2417) );
  INVX1 U3005 ( .A(n1635), .Y(n2418) );
  INVX1 U3006 ( .A(n1634), .Y(n2419) );
  INVX1 U3007 ( .A(n1609), .Y(n2420) );
  INVX1 U3008 ( .A(n1608), .Y(n2421) );
  INVX1 U3009 ( .A(n1607), .Y(n2422) );
  INVX1 U3010 ( .A(n1584), .Y(n2423) );
  INVX1 U3011 ( .A(n1583), .Y(n2424) );
  INVX1 U3012 ( .A(n1582), .Y(n2425) );
  INVX1 U3013 ( .A(n1557), .Y(n2426) );
  INVX1 U3014 ( .A(n1556), .Y(n2427) );
  INVX1 U3015 ( .A(n1555), .Y(n2428) );
  INVX1 U3016 ( .A(n1532), .Y(n2429) );
  INVX1 U3017 ( .A(n1531), .Y(n2430) );
  INVX1 U3018 ( .A(n1530), .Y(n2431) );
  INVX1 U3019 ( .A(n1505), .Y(n2432) );
  INVX1 U3020 ( .A(n1504), .Y(n2433) );
  INVX1 U3021 ( .A(n1503), .Y(n2434) );
  INVX1 U3022 ( .A(n1480), .Y(n2435) );
  INVX1 U3023 ( .A(n1479), .Y(n2436) );
  INVX1 U3024 ( .A(n1478), .Y(n2437) );
  INVX1 U3025 ( .A(n1453), .Y(n2438) );
  INVX1 U3026 ( .A(n1452), .Y(n2439) );
  INVX1 U3027 ( .A(n1451), .Y(n2440) );
  INVX1 U3028 ( .A(n1428), .Y(n2441) );
  INVX1 U3029 ( .A(n1427), .Y(n2442) );
  INVX1 U3030 ( .A(n1426), .Y(n2443) );
  INVX1 U3031 ( .A(n1400), .Y(n2444) );
  INVX1 U3032 ( .A(n1399), .Y(n2445) );
  INVX1 U3033 ( .A(n1398), .Y(n2446) );
  INVX1 U3034 ( .A(n1375), .Y(n2447) );
  INVX1 U3035 ( .A(n1374), .Y(n2448) );
  INVX1 U3036 ( .A(n1373), .Y(n2449) );
  BUFX2 U3037 ( .A(n1334), .Y(n3114) );
  BUFX2 U3038 ( .A(n1322), .Y(n3115) );
  BUFX2 U3039 ( .A(n1310), .Y(n3116) );
  BUFX2 U3040 ( .A(n1298), .Y(n3117) );
  BUFX2 U3041 ( .A(n1286), .Y(n3118) );
  BUFX2 U3042 ( .A(n1274), .Y(n3119) );
  BUFX2 U3043 ( .A(n1262), .Y(n3120) );
  BUFX2 U3044 ( .A(n1250), .Y(n3121) );
  BUFX2 U3045 ( .A(n1238), .Y(n3122) );
  BUFX2 U3046 ( .A(n1226), .Y(n3123) );
  BUFX2 U3047 ( .A(n1214), .Y(n3124) );
  BUFX2 U3048 ( .A(n1202), .Y(n3125) );
  BUFX2 U3049 ( .A(n1190), .Y(n3126) );
  BUFX2 U3050 ( .A(n1178), .Y(n3127) );
  BUFX2 U3051 ( .A(n1166), .Y(n3128) );
  BUFX2 U3052 ( .A(n1154), .Y(n3129) );
  BUFX2 U3053 ( .A(n1142), .Y(n3130) );
  BUFX2 U3054 ( .A(n1130), .Y(n3131) );
  BUFX2 U3055 ( .A(n1118), .Y(n3132) );
  BUFX2 U3056 ( .A(n1106), .Y(n3133) );
  BUFX2 U3057 ( .A(n1094), .Y(n3134) );
  BUFX2 U3058 ( .A(n1082), .Y(n3135) );
  BUFX2 U3059 ( .A(n1070), .Y(n3136) );
  BUFX2 U3060 ( .A(n1058), .Y(n3137) );
  BUFX2 U3061 ( .A(n1046), .Y(n3138) );
  BUFX2 U3062 ( .A(n1034), .Y(n3139) );
  BUFX2 U3063 ( .A(n1022), .Y(n3140) );
  BUFX2 U3064 ( .A(n1010), .Y(n3141) );
  BUFX2 U3065 ( .A(n998), .Y(n3142) );
  BUFX2 U3066 ( .A(n986), .Y(n3143) );
  BUFX2 U3067 ( .A(n974), .Y(n3144) );
  BUFX2 U3068 ( .A(n962), .Y(n3145) );
  BUFX2 U3069 ( .A(n950), .Y(n3146) );
  BUFX2 U3070 ( .A(n938), .Y(n3147) );
  BUFX2 U3071 ( .A(n926), .Y(n3148) );
  BUFX2 U3072 ( .A(n914), .Y(n3149) );
  BUFX2 U3073 ( .A(n902), .Y(n3150) );
  BUFX2 U3074 ( .A(n890), .Y(n3151) );
  BUFX2 U3075 ( .A(n878), .Y(n3152) );
  BUFX2 U3076 ( .A(n866), .Y(n3153) );
  BUFX2 U3077 ( .A(n854), .Y(n3154) );
  BUFX2 U3078 ( .A(n842), .Y(n3155) );
  BUFX2 U3079 ( .A(n830), .Y(n3156) );
  BUFX2 U3080 ( .A(n818), .Y(n3157) );
  BUFX2 U3081 ( .A(n806), .Y(n3158) );
  BUFX2 U3082 ( .A(n794), .Y(n3159) );
  BUFX2 U3083 ( .A(n782), .Y(n3160) );
  BUFX2 U3084 ( .A(n770), .Y(n3161) );
  BUFX2 U3085 ( .A(n758), .Y(n3162) );
  BUFX2 U3086 ( .A(n746), .Y(n3163) );
  BUFX2 U3087 ( .A(n734), .Y(n3164) );
  BUFX2 U3088 ( .A(n722), .Y(n3165) );
  BUFX2 U3089 ( .A(n710), .Y(n3166) );
  BUFX2 U3090 ( .A(n698), .Y(n3167) );
  BUFX2 U3091 ( .A(n686), .Y(n3168) );
  BUFX2 U3092 ( .A(n674), .Y(n3169) );
  BUFX2 U3093 ( .A(n662), .Y(n3170) );
  BUFX2 U3094 ( .A(n650), .Y(n3171) );
  BUFX2 U3095 ( .A(n638), .Y(n3172) );
  BUFX2 U3096 ( .A(n626), .Y(n3173) );
  BUFX2 U3097 ( .A(n613), .Y(n3174) );
  AND2X1 U3098 ( .A(enable), .B(n3708), .Y(n2450) );
  INVX1 U3099 ( .A(n2450), .Y(n2451) );
  BUFX2 U3100 ( .A(n625), .Y(n2452) );
  AND2X1 U3101 ( .A(n1756), .B(n3192), .Y(n2453) );
  INVX1 U3102 ( .A(n2453), .Y(n2454) );
  AND2X1 U3103 ( .A(n164), .B(n1749), .Y(n2455) );
  INVX1 U3104 ( .A(n2455), .Y(n2456) );
  AND2X1 U3105 ( .A(n2455), .B(n3178), .Y(n2457) );
  INVX1 U3106 ( .A(n2457), .Y(n2458) );
  AND2X1 U3107 ( .A(n1744), .B(n2453), .Y(n2459) );
  INVX1 U3108 ( .A(n2459), .Y(n2460) );
  AND2X1 U3109 ( .A(n3188), .B(n1749), .Y(n2461) );
  INVX1 U3110 ( .A(n2461), .Y(n2462) );
  AND2X1 U3111 ( .A(n3193), .B(n3187), .Y(n2463) );
  INVX1 U3112 ( .A(n2463), .Y(n2464) );
  AND2X1 U3113 ( .A(n3188), .B(n1748), .Y(n2465) );
  INVX1 U3114 ( .A(n2465), .Y(n2466) );
  AND2X1 U3115 ( .A(n3188), .B(n1747), .Y(n2467) );
  INVX1 U3116 ( .A(n2467), .Y(n2468) );
  AND2X1 U3117 ( .A(n3188), .B(n1746), .Y(n2469) );
  INVX1 U3118 ( .A(n2469), .Y(n2470) );
  AND2X1 U3119 ( .A(n3188), .B(n1745), .Y(n2471) );
  INVX1 U3120 ( .A(n2471), .Y(n2472) );
  AND2X1 U3121 ( .A(n3188), .B(n1744), .Y(n2473) );
  INVX1 U3122 ( .A(n2473), .Y(n2474) );
  AND2X1 U3123 ( .A(n3188), .B(n1743), .Y(n2475) );
  INVX1 U3124 ( .A(n2475), .Y(n2476) );
  AND2X1 U3125 ( .A(n3193), .B(n1749), .Y(n2477) );
  INVX1 U3126 ( .A(n2477), .Y(n2478) );
  AND2X1 U3127 ( .A(n162), .B(n3187), .Y(n2479) );
  INVX1 U3128 ( .A(n2479), .Y(n2480) );
  AND2X1 U3129 ( .A(n3193), .B(n1748), .Y(n2481) );
  INVX1 U3130 ( .A(n2481), .Y(n2482) );
  AND2X1 U3131 ( .A(n3193), .B(n1747), .Y(n2483) );
  INVX1 U3132 ( .A(n2483), .Y(n2484) );
  AND2X1 U3133 ( .A(n3193), .B(n1746), .Y(n2485) );
  INVX1 U3134 ( .A(n2485), .Y(n2486) );
  AND2X1 U3135 ( .A(n3193), .B(n1745), .Y(n2487) );
  INVX1 U3136 ( .A(n2487), .Y(n2488) );
  AND2X1 U3137 ( .A(n3193), .B(n1744), .Y(n2489) );
  INVX1 U3138 ( .A(n2489), .Y(n2490) );
  AND2X1 U3139 ( .A(n3193), .B(n1743), .Y(n2491) );
  INVX1 U3140 ( .A(n2491), .Y(n2492) );
  AND2X1 U3141 ( .A(n162), .B(n1749), .Y(n2493) );
  INVX1 U3142 ( .A(n2493), .Y(n2494) );
  AND2X1 U3143 ( .A(n164), .B(n3187), .Y(n2495) );
  INVX1 U3144 ( .A(n2495), .Y(n2496) );
  AND2X1 U3145 ( .A(n162), .B(n1748), .Y(n2497) );
  INVX1 U3146 ( .A(n2497), .Y(n2498) );
  AND2X1 U3147 ( .A(n162), .B(n1747), .Y(n2499) );
  INVX1 U3148 ( .A(n2499), .Y(n2500) );
  AND2X1 U3149 ( .A(n162), .B(n1746), .Y(n2501) );
  INVX1 U3150 ( .A(n2501), .Y(n2502) );
  AND2X1 U3151 ( .A(n162), .B(n1745), .Y(n2503) );
  INVX1 U3152 ( .A(n2503), .Y(n2504) );
  AND2X1 U3153 ( .A(n162), .B(n1744), .Y(n2505) );
  INVX1 U3154 ( .A(n2505), .Y(n2506) );
  AND2X1 U3155 ( .A(n162), .B(n1743), .Y(n2507) );
  INVX1 U3156 ( .A(n2507), .Y(n2508) );
  AND2X1 U3157 ( .A(n164), .B(n1748), .Y(n2509) );
  INVX1 U3158 ( .A(n2509), .Y(n2510) );
  AND2X1 U3159 ( .A(n164), .B(n1746), .Y(n2511) );
  INVX1 U3160 ( .A(n2511), .Y(n2512) );
  AND2X1 U3161 ( .A(n164), .B(n1745), .Y(n2513) );
  INVX1 U3162 ( .A(n2513), .Y(n2514) );
  AND2X1 U3163 ( .A(n164), .B(n1744), .Y(n2515) );
  INVX1 U3164 ( .A(n2515), .Y(n2516) );
  AND2X1 U3165 ( .A(n164), .B(n1743), .Y(n2517) );
  INVX1 U3166 ( .A(n2517), .Y(n2518) );
  AND2X1 U3167 ( .A(n3189), .B(n1749), .Y(n2519) );
  INVX1 U3168 ( .A(n2519), .Y(n2520) );
  AND2X1 U3169 ( .A(n3191), .B(n3187), .Y(n2521) );
  INVX1 U3170 ( .A(n2521), .Y(n2522) );
  AND2X1 U3171 ( .A(n3189), .B(n1748), .Y(n2523) );
  INVX1 U3172 ( .A(n2523), .Y(n2524) );
  AND2X1 U3173 ( .A(n3189), .B(n1747), .Y(n2525) );
  INVX1 U3174 ( .A(n2525), .Y(n2526) );
  AND2X1 U3175 ( .A(n3189), .B(n1746), .Y(n2527) );
  INVX1 U3176 ( .A(n2527), .Y(n2528) );
  AND2X1 U3177 ( .A(n3189), .B(n1745), .Y(n2529) );
  INVX1 U3178 ( .A(n2529), .Y(n2530) );
  AND2X1 U3179 ( .A(n3189), .B(n1744), .Y(n2531) );
  INVX1 U3180 ( .A(n2531), .Y(n2532) );
  AND2X1 U3181 ( .A(n3189), .B(n1743), .Y(n2533) );
  INVX1 U3182 ( .A(n2533), .Y(n2534) );
  INVX1 U3183 ( .A(n2536), .Y(n2535) );
  AND2X1 U3184 ( .A(n3191), .B(n1749), .Y(n2536) );
  AND2X1 U3185 ( .A(n3188), .B(n3187), .Y(n2537) );
  INVX1 U3186 ( .A(n2537), .Y(n2538) );
  AND2X1 U3187 ( .A(n3191), .B(n1748), .Y(n2539) );
  INVX1 U3188 ( .A(n2539), .Y(n2540) );
  AND2X1 U3189 ( .A(n3191), .B(n1747), .Y(n2541) );
  INVX1 U3190 ( .A(n2541), .Y(n2542) );
  AND2X1 U3191 ( .A(n3191), .B(n1746), .Y(n2543) );
  INVX1 U3192 ( .A(n2543), .Y(n2544) );
  AND2X1 U3193 ( .A(n3191), .B(n1745), .Y(n2545) );
  INVX1 U3194 ( .A(n2545), .Y(n2546) );
  AND2X1 U3195 ( .A(n3191), .B(n1744), .Y(n2547) );
  INVX1 U3196 ( .A(n2547), .Y(n2548) );
  AND2X1 U3197 ( .A(n3191), .B(n1743), .Y(n2549) );
  INVX1 U3198 ( .A(n2549), .Y(n2550) );
  AND2X1 U3199 ( .A(n1749), .B(n2453), .Y(n2551) );
  INVX1 U3200 ( .A(n2551), .Y(n2552) );
  AND2X1 U3201 ( .A(n3190), .B(n3187), .Y(n2553) );
  INVX1 U3202 ( .A(n2553), .Y(n2554) );
  AND2X1 U3203 ( .A(n1748), .B(n2453), .Y(n2555) );
  INVX1 U3204 ( .A(n2555), .Y(n2556) );
  AND2X1 U3205 ( .A(n1747), .B(n2453), .Y(n2557) );
  INVX1 U3206 ( .A(n2557), .Y(n2558) );
  AND2X1 U3207 ( .A(n1746), .B(n2453), .Y(n2559) );
  INVX1 U3208 ( .A(n2559), .Y(n2560) );
  AND2X1 U3209 ( .A(n1745), .B(n2453), .Y(n2561) );
  INVX1 U3210 ( .A(n2561), .Y(n2562) );
  AND2X1 U3211 ( .A(n1743), .B(n2453), .Y(n2563) );
  INVX1 U3212 ( .A(n2563), .Y(n2564) );
  AND2X1 U3213 ( .A(n3190), .B(n1749), .Y(n2565) );
  INVX1 U3214 ( .A(n2565), .Y(n2566) );
  AND2X1 U3215 ( .A(n3189), .B(n3187), .Y(n2567) );
  INVX1 U3216 ( .A(n2567), .Y(n2568) );
  AND2X1 U3217 ( .A(n3190), .B(n1748), .Y(n2569) );
  INVX1 U3218 ( .A(n2569), .Y(n2570) );
  AND2X1 U3219 ( .A(n3190), .B(n1747), .Y(n2571) );
  INVX1 U3220 ( .A(n2571), .Y(n2572) );
  AND2X1 U3221 ( .A(n3190), .B(n1746), .Y(n2573) );
  INVX1 U3222 ( .A(n2573), .Y(n2574) );
  AND2X1 U3223 ( .A(n3190), .B(n1745), .Y(n2575) );
  INVX1 U3224 ( .A(n2575), .Y(n2576) );
  AND2X1 U3225 ( .A(n3190), .B(n1744), .Y(n2577) );
  INVX1 U3226 ( .A(n2577), .Y(n2578) );
  AND2X1 U3227 ( .A(n3190), .B(n1743), .Y(n2579) );
  INVX1 U3228 ( .A(n2579), .Y(n2580) );
  AND2X1 U3229 ( .A(n164), .B(n1747), .Y(n2581) );
  INVX1 U3230 ( .A(n2581), .Y(n2582) );
  MUX2X1 U3231 ( .B(n2584), .A(n2585), .S(n3083), .Y(n2583) );
  MUX2X1 U3232 ( .B(n2587), .A(n2588), .S(n3088), .Y(n2586) );
  MUX2X1 U3233 ( .B(n2590), .A(n2591), .S(n3089), .Y(n2589) );
  MUX2X1 U3234 ( .B(n2593), .A(n2594), .S(n3089), .Y(n2592) );
  MUX2X1 U3235 ( .B(n2596), .A(n2597), .S(N180), .Y(n2595) );
  MUX2X1 U3236 ( .B(n2599), .A(n2600), .S(n3083), .Y(n2598) );
  MUX2X1 U3237 ( .B(n2602), .A(n2603), .S(n3083), .Y(n2601) );
  MUX2X1 U3238 ( .B(n2605), .A(n2606), .S(n3083), .Y(n2604) );
  MUX2X1 U3239 ( .B(n2608), .A(n2609), .S(n3089), .Y(n2607) );
  MUX2X1 U3240 ( .B(n2611), .A(n2612), .S(N180), .Y(n2610) );
  MUX2X1 U3241 ( .B(n2614), .A(n2615), .S(n3083), .Y(n2613) );
  MUX2X1 U3242 ( .B(n2617), .A(n2618), .S(n3083), .Y(n2616) );
  MUX2X1 U3243 ( .B(n2620), .A(n2621), .S(n3083), .Y(n2619) );
  MUX2X1 U3244 ( .B(n2623), .A(n2624), .S(n3083), .Y(n2622) );
  MUX2X1 U3245 ( .B(n2626), .A(n2627), .S(N180), .Y(n2625) );
  MUX2X1 U3246 ( .B(n2629), .A(n2630), .S(n3083), .Y(n2628) );
  MUX2X1 U3247 ( .B(n2632), .A(n2633), .S(n3083), .Y(n2631) );
  MUX2X1 U3248 ( .B(n2635), .A(n2636), .S(n3083), .Y(n2634) );
  MUX2X1 U3249 ( .B(n2638), .A(n2639), .S(n3083), .Y(n2637) );
  MUX2X1 U3250 ( .B(n2641), .A(n2642), .S(N180), .Y(n2640) );
  MUX2X1 U3251 ( .B(n2643), .A(n2644), .S(N182), .Y(N192) );
  MUX2X1 U3252 ( .B(n2646), .A(n2647), .S(n3083), .Y(n2645) );
  MUX2X1 U3253 ( .B(n2649), .A(n2650), .S(n3083), .Y(n2648) );
  MUX2X1 U3254 ( .B(n2652), .A(n2653), .S(n3083), .Y(n2651) );
  MUX2X1 U3255 ( .B(n2655), .A(n2656), .S(n3083), .Y(n2654) );
  MUX2X1 U3256 ( .B(n2658), .A(n2659), .S(N180), .Y(n2657) );
  MUX2X1 U3257 ( .B(n2661), .A(n2662), .S(n3087), .Y(n2660) );
  MUX2X1 U3258 ( .B(n2664), .A(n2665), .S(n3089), .Y(n2663) );
  MUX2X1 U3259 ( .B(n2667), .A(n2668), .S(n3087), .Y(n2666) );
  MUX2X1 U3260 ( .B(n2670), .A(n2671), .S(n3089), .Y(n2669) );
  MUX2X1 U3261 ( .B(n2673), .A(n2674), .S(N180), .Y(n2672) );
  MUX2X1 U3262 ( .B(n2676), .A(n2677), .S(n3089), .Y(n2675) );
  MUX2X1 U3263 ( .B(n2679), .A(n2680), .S(n3089), .Y(n2678) );
  MUX2X1 U3264 ( .B(n2682), .A(n2683), .S(n3083), .Y(n2681) );
  MUX2X1 U3265 ( .B(n2685), .A(n2686), .S(n3086), .Y(n2684) );
  MUX2X1 U3266 ( .B(n2688), .A(n2689), .S(N180), .Y(n2687) );
  MUX2X1 U3267 ( .B(n2691), .A(n2692), .S(n3086), .Y(n2690) );
  MUX2X1 U3268 ( .B(n2694), .A(n2695), .S(n3083), .Y(n2693) );
  MUX2X1 U3269 ( .B(n2697), .A(n2698), .S(n3088), .Y(n2696) );
  MUX2X1 U3270 ( .B(n2700), .A(n2701), .S(n3083), .Y(n2699) );
  MUX2X1 U3271 ( .B(n2703), .A(n2704), .S(N180), .Y(n2702) );
  MUX2X1 U3272 ( .B(n2705), .A(n2706), .S(N182), .Y(N191) );
  MUX2X1 U3273 ( .B(n2708), .A(n2709), .S(n3084), .Y(n2707) );
  MUX2X1 U3274 ( .B(n2711), .A(n2712), .S(n3084), .Y(n2710) );
  MUX2X1 U3275 ( .B(n2714), .A(n2715), .S(n3084), .Y(n2713) );
  MUX2X1 U3276 ( .B(n2717), .A(n2718), .S(n3084), .Y(n2716) );
  MUX2X1 U3277 ( .B(n2720), .A(n2721), .S(N180), .Y(n2719) );
  MUX2X1 U3278 ( .B(n2723), .A(n2724), .S(n3084), .Y(n2722) );
  MUX2X1 U3279 ( .B(n2726), .A(n2727), .S(n3084), .Y(n2725) );
  MUX2X1 U3280 ( .B(n2729), .A(n2730), .S(n3084), .Y(n2728) );
  MUX2X1 U3281 ( .B(n2732), .A(n2733), .S(n3084), .Y(n2731) );
  MUX2X1 U3282 ( .B(n2735), .A(n2736), .S(N180), .Y(n2734) );
  MUX2X1 U3283 ( .B(n2738), .A(n2739), .S(n3084), .Y(n2737) );
  MUX2X1 U3284 ( .B(n2741), .A(n2742), .S(n3084), .Y(n2740) );
  MUX2X1 U3285 ( .B(n2744), .A(n2745), .S(n3084), .Y(n2743) );
  MUX2X1 U3286 ( .B(n2747), .A(n2748), .S(n3084), .Y(n2746) );
  MUX2X1 U3287 ( .B(n2750), .A(n2751), .S(N180), .Y(n2749) );
  MUX2X1 U3288 ( .B(n2753), .A(n2754), .S(n3085), .Y(n2752) );
  MUX2X1 U3289 ( .B(n2756), .A(n2757), .S(n3085), .Y(n2755) );
  MUX2X1 U3290 ( .B(n2759), .A(n2760), .S(n3085), .Y(n2758) );
  MUX2X1 U3291 ( .B(n2762), .A(n2763), .S(n3085), .Y(n2761) );
  MUX2X1 U3292 ( .B(n2765), .A(n2766), .S(N180), .Y(n2764) );
  MUX2X1 U3293 ( .B(n2767), .A(n2768), .S(N182), .Y(N190) );
  MUX2X1 U3294 ( .B(n2770), .A(n2771), .S(n3085), .Y(n2769) );
  MUX2X1 U3295 ( .B(n2773), .A(n2774), .S(n3085), .Y(n2772) );
  MUX2X1 U3296 ( .B(n2776), .A(n2777), .S(n3085), .Y(n2775) );
  MUX2X1 U3297 ( .B(n2779), .A(n2780), .S(n3085), .Y(n2778) );
  MUX2X1 U3298 ( .B(n2782), .A(n2783), .S(N180), .Y(n2781) );
  MUX2X1 U3299 ( .B(n2785), .A(n2786), .S(n3085), .Y(n2784) );
  MUX2X1 U3300 ( .B(n2788), .A(n2789), .S(n3085), .Y(n2787) );
  MUX2X1 U3301 ( .B(n2791), .A(n2792), .S(n3085), .Y(n2790) );
  MUX2X1 U3302 ( .B(n2794), .A(n2795), .S(n3085), .Y(n2793) );
  MUX2X1 U3303 ( .B(n2797), .A(n2798), .S(N180), .Y(n2796) );
  MUX2X1 U3304 ( .B(n2800), .A(n2801), .S(n3084), .Y(n2799) );
  MUX2X1 U3305 ( .B(n2803), .A(n2804), .S(n3085), .Y(n2802) );
  MUX2X1 U3306 ( .B(n2806), .A(n2807), .S(n3085), .Y(n2805) );
  MUX2X1 U3307 ( .B(n2809), .A(n2810), .S(n3084), .Y(n2808) );
  MUX2X1 U3308 ( .B(n2812), .A(n2813), .S(N180), .Y(n2811) );
  MUX2X1 U3309 ( .B(n2815), .A(n2816), .S(n3084), .Y(n2814) );
  MUX2X1 U3310 ( .B(n2818), .A(n2819), .S(n3084), .Y(n2817) );
  MUX2X1 U3311 ( .B(n2821), .A(n2822), .S(n3085), .Y(n2820) );
  MUX2X1 U3312 ( .B(n2824), .A(n2825), .S(n3084), .Y(n2823) );
  MUX2X1 U3313 ( .B(n2827), .A(n2828), .S(N180), .Y(n2826) );
  MUX2X1 U3314 ( .B(n2829), .A(n2830), .S(N182), .Y(N189) );
  MUX2X1 U3315 ( .B(n2832), .A(n2833), .S(n3084), .Y(n2831) );
  MUX2X1 U3316 ( .B(n2835), .A(n2836), .S(n3084), .Y(n2834) );
  MUX2X1 U3317 ( .B(n2838), .A(n2839), .S(n3085), .Y(n2837) );
  MUX2X1 U3318 ( .B(n2841), .A(n2842), .S(n3085), .Y(n2840) );
  MUX2X1 U3319 ( .B(n2844), .A(n2845), .S(N180), .Y(n2843) );
  MUX2X1 U3320 ( .B(n2847), .A(n2848), .S(n3086), .Y(n2846) );
  MUX2X1 U3321 ( .B(n2850), .A(n2851), .S(n3086), .Y(n2849) );
  MUX2X1 U3322 ( .B(n2853), .A(n2854), .S(n3086), .Y(n2852) );
  MUX2X1 U3323 ( .B(n2856), .A(n2857), .S(n3086), .Y(n2855) );
  MUX2X1 U3324 ( .B(n2859), .A(n2860), .S(N180), .Y(n2858) );
  MUX2X1 U3325 ( .B(n2862), .A(n2863), .S(n3086), .Y(n2861) );
  MUX2X1 U3326 ( .B(n2865), .A(n2866), .S(n3086), .Y(n2864) );
  MUX2X1 U3327 ( .B(n2868), .A(n2869), .S(n3086), .Y(n2867) );
  MUX2X1 U3328 ( .B(n2871), .A(n2872), .S(n3086), .Y(n2870) );
  MUX2X1 U3329 ( .B(n2874), .A(n2875), .S(N180), .Y(n2873) );
  MUX2X1 U3330 ( .B(n2877), .A(n2878), .S(n3086), .Y(n2876) );
  MUX2X1 U3331 ( .B(n2880), .A(n2881), .S(n3086), .Y(n2879) );
  MUX2X1 U3332 ( .B(n2883), .A(n2884), .S(n3086), .Y(n2882) );
  MUX2X1 U3333 ( .B(n2886), .A(n2887), .S(n3086), .Y(n2885) );
  MUX2X1 U3334 ( .B(n2889), .A(n2890), .S(N180), .Y(n2888) );
  MUX2X1 U3335 ( .B(n2891), .A(n2892), .S(N182), .Y(N188) );
  MUX2X1 U3336 ( .B(n2894), .A(n2895), .S(n3087), .Y(n2893) );
  MUX2X1 U3337 ( .B(n2897), .A(n2898), .S(n3087), .Y(n2896) );
  MUX2X1 U3338 ( .B(n2900), .A(n2901), .S(n3087), .Y(n2899) );
  MUX2X1 U3339 ( .B(n2903), .A(n2904), .S(n3087), .Y(n2902) );
  MUX2X1 U3340 ( .B(n2906), .A(n2907), .S(N180), .Y(n2905) );
  MUX2X1 U3341 ( .B(n2909), .A(n2910), .S(n3087), .Y(n2908) );
  MUX2X1 U3342 ( .B(n2912), .A(n2913), .S(n3087), .Y(n2911) );
  MUX2X1 U3343 ( .B(n2915), .A(n2916), .S(n3087), .Y(n2914) );
  MUX2X1 U3344 ( .B(n2918), .A(n2919), .S(n3087), .Y(n2917) );
  MUX2X1 U3345 ( .B(n2921), .A(n2922), .S(N180), .Y(n2920) );
  MUX2X1 U3346 ( .B(n2924), .A(n2925), .S(n3087), .Y(n2923) );
  MUX2X1 U3347 ( .B(n2927), .A(n2928), .S(n3087), .Y(n2926) );
  MUX2X1 U3348 ( .B(n2930), .A(n2931), .S(n3087), .Y(n2929) );
  MUX2X1 U3349 ( .B(n2933), .A(n2934), .S(n3087), .Y(n2932) );
  MUX2X1 U3350 ( .B(n2936), .A(n2937), .S(N180), .Y(n2935) );
  MUX2X1 U3351 ( .B(n2939), .A(n2940), .S(n3088), .Y(n2938) );
  MUX2X1 U3352 ( .B(n2942), .A(n2943), .S(n3088), .Y(n2941) );
  MUX2X1 U3353 ( .B(n2945), .A(n2946), .S(n3088), .Y(n2944) );
  MUX2X1 U3354 ( .B(n2948), .A(n2949), .S(n3088), .Y(n2947) );
  MUX2X1 U3355 ( .B(n2951), .A(n2952), .S(N180), .Y(n2950) );
  MUX2X1 U3356 ( .B(n2953), .A(n2954), .S(N182), .Y(N187) );
  MUX2X1 U3357 ( .B(n2956), .A(n2957), .S(n3088), .Y(n2955) );
  MUX2X1 U3358 ( .B(n2959), .A(n2960), .S(n3088), .Y(n2958) );
  MUX2X1 U3359 ( .B(n2962), .A(n2963), .S(n3088), .Y(n2961) );
  MUX2X1 U3360 ( .B(n2965), .A(n2966), .S(n3088), .Y(n2964) );
  MUX2X1 U3361 ( .B(n2968), .A(n2969), .S(N180), .Y(n2967) );
  MUX2X1 U3362 ( .B(n2971), .A(n2972), .S(n3088), .Y(n2970) );
  MUX2X1 U3363 ( .B(n2974), .A(n2975), .S(n3088), .Y(n2973) );
  MUX2X1 U3364 ( .B(n2977), .A(n2978), .S(n3088), .Y(n2976) );
  MUX2X1 U3365 ( .B(n2980), .A(n2981), .S(n3088), .Y(n2979) );
  MUX2X1 U3366 ( .B(n2983), .A(n2984), .S(N180), .Y(n2982) );
  MUX2X1 U3367 ( .B(n2986), .A(n2987), .S(n3087), .Y(n2985) );
  MUX2X1 U3368 ( .B(n2989), .A(n2990), .S(n3087), .Y(n2988) );
  MUX2X1 U3369 ( .B(n2992), .A(n2993), .S(n3086), .Y(n2991) );
  MUX2X1 U3370 ( .B(n2995), .A(n2996), .S(n3087), .Y(n2994) );
  MUX2X1 U3371 ( .B(n2998), .A(n2999), .S(N180), .Y(n2997) );
  MUX2X1 U3372 ( .B(n3001), .A(n3002), .S(n3086), .Y(n3000) );
  MUX2X1 U3373 ( .B(n3004), .A(n3005), .S(n3087), .Y(n3003) );
  MUX2X1 U3374 ( .B(n3007), .A(n3008), .S(n3088), .Y(n3006) );
  MUX2X1 U3375 ( .B(n3010), .A(n3011), .S(n3088), .Y(n3009) );
  MUX2X1 U3376 ( .B(n3013), .A(n3014), .S(N180), .Y(n3012) );
  MUX2X1 U3377 ( .B(n3015), .A(n3016), .S(N182), .Y(N186) );
  MUX2X1 U3378 ( .B(n3018), .A(n3019), .S(n3086), .Y(n3017) );
  MUX2X1 U3379 ( .B(n3021), .A(n3022), .S(n3086), .Y(n3020) );
  MUX2X1 U3380 ( .B(n3024), .A(n3025), .S(n3088), .Y(n3023) );
  MUX2X1 U3381 ( .B(n3027), .A(n3028), .S(n3088), .Y(n3026) );
  MUX2X1 U3382 ( .B(n3030), .A(n3031), .S(N180), .Y(n3029) );
  MUX2X1 U3383 ( .B(n3033), .A(n3034), .S(n3089), .Y(n3032) );
  MUX2X1 U3384 ( .B(n3036), .A(n3037), .S(n3089), .Y(n3035) );
  MUX2X1 U3385 ( .B(n3039), .A(n3040), .S(n3089), .Y(n3038) );
  MUX2X1 U3386 ( .B(n3042), .A(n3043), .S(n3089), .Y(n3041) );
  MUX2X1 U3387 ( .B(n3045), .A(n3046), .S(N180), .Y(n3044) );
  MUX2X1 U3388 ( .B(n3048), .A(n3049), .S(n3089), .Y(n3047) );
  MUX2X1 U3389 ( .B(n3051), .A(n3052), .S(n3089), .Y(n3050) );
  MUX2X1 U3390 ( .B(n3054), .A(n3055), .S(n3089), .Y(n3053) );
  MUX2X1 U3391 ( .B(n3057), .A(n3058), .S(n3089), .Y(n3056) );
  MUX2X1 U3392 ( .B(n3060), .A(n3061), .S(N180), .Y(n3059) );
  MUX2X1 U3393 ( .B(n3063), .A(n3064), .S(n3089), .Y(n3062) );
  MUX2X1 U3394 ( .B(n3066), .A(n3067), .S(n3089), .Y(n3065) );
  MUX2X1 U3395 ( .B(n3069), .A(n3070), .S(n3089), .Y(n3068) );
  MUX2X1 U3396 ( .B(n3072), .A(n3073), .S(n3089), .Y(n3071) );
  MUX2X1 U3397 ( .B(n3075), .A(n3076), .S(N180), .Y(n3074) );
  MUX2X1 U3398 ( .B(n3077), .A(n3078), .S(N182), .Y(N185) );
  MUX2X1 U3399 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n3095), .Y(n2585) );
  MUX2X1 U3400 ( .B(\mem<60><0> ), .A(\mem<61><0> ), .S(n3094), .Y(n2584) );
  MUX2X1 U3401 ( .B(\mem<58><0> ), .A(\mem<59><0> ), .S(n3095), .Y(n2588) );
  MUX2X1 U3402 ( .B(\mem<56><0> ), .A(\mem<57><0> ), .S(n3094), .Y(n2587) );
  MUX2X1 U3403 ( .B(n2586), .A(n2583), .S(n3082), .Y(n2597) );
  MUX2X1 U3404 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n3094), .Y(n2591) );
  MUX2X1 U3405 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n3094), .Y(n2590) );
  MUX2X1 U3406 ( .B(\mem<50><0> ), .A(\mem<51><0> ), .S(n3094), .Y(n2594) );
  MUX2X1 U3407 ( .B(\mem<48><0> ), .A(\mem<49><0> ), .S(n3094), .Y(n2593) );
  MUX2X1 U3408 ( .B(n2592), .A(n2589), .S(n3082), .Y(n2596) );
  MUX2X1 U3409 ( .B(\mem<46><0> ), .A(\mem<47><0> ), .S(n3094), .Y(n2600) );
  MUX2X1 U3410 ( .B(\mem<44><0> ), .A(\mem<45><0> ), .S(n3094), .Y(n2599) );
  MUX2X1 U3411 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n3094), .Y(n2603) );
  MUX2X1 U3412 ( .B(\mem<40><0> ), .A(\mem<41><0> ), .S(n3094), .Y(n2602) );
  MUX2X1 U3413 ( .B(n2601), .A(n2598), .S(n3082), .Y(n2612) );
  MUX2X1 U3414 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n3094), .Y(n2606) );
  MUX2X1 U3415 ( .B(\mem<36><0> ), .A(\mem<37><0> ), .S(n3094), .Y(n2605) );
  MUX2X1 U3416 ( .B(\mem<34><0> ), .A(\mem<35><0> ), .S(n3094), .Y(n2609) );
  MUX2X1 U3417 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n3094), .Y(n2608) );
  MUX2X1 U3418 ( .B(n2607), .A(n2604), .S(n3082), .Y(n2611) );
  MUX2X1 U3419 ( .B(n2610), .A(n2595), .S(N181), .Y(n2644) );
  MUX2X1 U3420 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n3095), .Y(n2615) );
  MUX2X1 U3421 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n3095), .Y(n2614) );
  MUX2X1 U3422 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n3095), .Y(n2618) );
  MUX2X1 U3423 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n3095), .Y(n2617) );
  MUX2X1 U3424 ( .B(n2616), .A(n2613), .S(n3082), .Y(n2627) );
  MUX2X1 U3425 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n3095), .Y(n2621) );
  MUX2X1 U3426 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n3095), .Y(n2620) );
  MUX2X1 U3427 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n3095), .Y(n2624) );
  MUX2X1 U3428 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n3095), .Y(n2623) );
  MUX2X1 U3429 ( .B(n2622), .A(n2619), .S(n3082), .Y(n2626) );
  MUX2X1 U3430 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n3095), .Y(n2630) );
  MUX2X1 U3431 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n3095), .Y(n2629) );
  MUX2X1 U3432 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n3095), .Y(n2633) );
  MUX2X1 U3433 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n3095), .Y(n2632) );
  MUX2X1 U3434 ( .B(n2631), .A(n2628), .S(n3082), .Y(n2642) );
  MUX2X1 U3435 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n3096), .Y(n2636) );
  MUX2X1 U3436 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n3096), .Y(n2635) );
  MUX2X1 U3437 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n3096), .Y(n2639) );
  MUX2X1 U3438 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n3096), .Y(n2638) );
  MUX2X1 U3439 ( .B(n2637), .A(n2634), .S(n3082), .Y(n2641) );
  MUX2X1 U3440 ( .B(n2640), .A(n2625), .S(N181), .Y(n2643) );
  MUX2X1 U3441 ( .B(\mem<62><1> ), .A(\mem<63><1> ), .S(n3096), .Y(n2647) );
  MUX2X1 U3442 ( .B(\mem<60><1> ), .A(\mem<61><1> ), .S(n3096), .Y(n2646) );
  MUX2X1 U3443 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n3096), .Y(n2650) );
  MUX2X1 U3444 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n3096), .Y(n2649) );
  MUX2X1 U3445 ( .B(n2648), .A(n2645), .S(n3082), .Y(n2659) );
  MUX2X1 U3446 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n3096), .Y(n2653) );
  MUX2X1 U3447 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n3096), .Y(n2652) );
  MUX2X1 U3448 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n3096), .Y(n2656) );
  MUX2X1 U3449 ( .B(\mem<48><1> ), .A(\mem<49><1> ), .S(n3096), .Y(n2655) );
  MUX2X1 U3450 ( .B(n2654), .A(n2651), .S(n3082), .Y(n2658) );
  MUX2X1 U3451 ( .B(\mem<46><1> ), .A(\mem<47><1> ), .S(n3097), .Y(n2662) );
  MUX2X1 U3452 ( .B(\mem<44><1> ), .A(\mem<45><1> ), .S(n3097), .Y(n2661) );
  MUX2X1 U3453 ( .B(\mem<42><1> ), .A(\mem<43><1> ), .S(n3097), .Y(n2665) );
  MUX2X1 U3454 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n3097), .Y(n2664) );
  MUX2X1 U3455 ( .B(n2663), .A(n2660), .S(n3082), .Y(n2674) );
  MUX2X1 U3456 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n3097), .Y(n2668) );
  MUX2X1 U3457 ( .B(\mem<36><1> ), .A(\mem<37><1> ), .S(n3097), .Y(n2667) );
  MUX2X1 U3458 ( .B(\mem<34><1> ), .A(\mem<35><1> ), .S(n3097), .Y(n2671) );
  MUX2X1 U3459 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n3097), .Y(n2670) );
  MUX2X1 U3460 ( .B(n2669), .A(n2666), .S(n3082), .Y(n2673) );
  MUX2X1 U3461 ( .B(n2672), .A(n2657), .S(N181), .Y(n2706) );
  MUX2X1 U3462 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n3097), .Y(n2677) );
  MUX2X1 U3463 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n3097), .Y(n2676) );
  MUX2X1 U3464 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n3097), .Y(n2680) );
  MUX2X1 U3465 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n3097), .Y(n2679) );
  MUX2X1 U3466 ( .B(n2678), .A(n2675), .S(n3081), .Y(n2689) );
  MUX2X1 U3467 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n3098), .Y(n2683) );
  MUX2X1 U3468 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n3098), .Y(n2682) );
  MUX2X1 U3469 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n3098), .Y(n2686) );
  MUX2X1 U3470 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n3098), .Y(n2685) );
  MUX2X1 U3471 ( .B(n2684), .A(n2681), .S(n3081), .Y(n2688) );
  MUX2X1 U3472 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n3098), .Y(n2692) );
  MUX2X1 U3473 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n3098), .Y(n2691) );
  MUX2X1 U3474 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n3098), .Y(n2695) );
  MUX2X1 U3475 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n3098), .Y(n2694) );
  MUX2X1 U3476 ( .B(n2693), .A(n2690), .S(n3081), .Y(n2704) );
  MUX2X1 U3477 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n3098), .Y(n2698) );
  MUX2X1 U3478 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n3098), .Y(n2697) );
  MUX2X1 U3479 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n3098), .Y(n2701) );
  MUX2X1 U3480 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n3098), .Y(n2700) );
  MUX2X1 U3481 ( .B(n2699), .A(n2696), .S(n3081), .Y(n2703) );
  MUX2X1 U3482 ( .B(n2702), .A(n2687), .S(N181), .Y(n2705) );
  MUX2X1 U3483 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n3099), .Y(n2709) );
  MUX2X1 U3484 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n3099), .Y(n2708) );
  MUX2X1 U3485 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n3099), .Y(n2712) );
  MUX2X1 U3486 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n3099), .Y(n2711) );
  MUX2X1 U3487 ( .B(n2710), .A(n2707), .S(n3081), .Y(n2721) );
  MUX2X1 U3488 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n3099), .Y(n2715) );
  MUX2X1 U3489 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n3099), .Y(n2714) );
  MUX2X1 U3490 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n3099), .Y(n2718) );
  MUX2X1 U3491 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n3099), .Y(n2717) );
  MUX2X1 U3492 ( .B(n2716), .A(n2713), .S(n3081), .Y(n2720) );
  MUX2X1 U3493 ( .B(\mem<46><2> ), .A(\mem<47><2> ), .S(n3099), .Y(n2724) );
  MUX2X1 U3494 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n3099), .Y(n2723) );
  MUX2X1 U3495 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n3099), .Y(n2727) );
  MUX2X1 U3496 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n3099), .Y(n2726) );
  MUX2X1 U3497 ( .B(n2725), .A(n2722), .S(n3081), .Y(n2736) );
  MUX2X1 U3498 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n3100), .Y(n2730) );
  MUX2X1 U3499 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n3100), .Y(n2729) );
  MUX2X1 U3500 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n3100), .Y(n2733) );
  MUX2X1 U3501 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n3100), .Y(n2732) );
  MUX2X1 U3502 ( .B(n2731), .A(n2728), .S(n3081), .Y(n2735) );
  MUX2X1 U3503 ( .B(n2734), .A(n2719), .S(N181), .Y(n2768) );
  MUX2X1 U3504 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n3100), .Y(n2739) );
  MUX2X1 U3505 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n3100), .Y(n2738) );
  MUX2X1 U3506 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n3100), .Y(n2742) );
  MUX2X1 U3507 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n3100), .Y(n2741) );
  MUX2X1 U3508 ( .B(n2740), .A(n2737), .S(n3081), .Y(n2751) );
  MUX2X1 U3509 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n3100), .Y(n2745) );
  MUX2X1 U3510 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n3100), .Y(n2744) );
  MUX2X1 U3511 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n3100), .Y(n2748) );
  MUX2X1 U3512 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n3100), .Y(n2747) );
  MUX2X1 U3513 ( .B(n2746), .A(n2743), .S(n3081), .Y(n2750) );
  MUX2X1 U3514 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n3096), .Y(n2754) );
  MUX2X1 U3515 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n3096), .Y(n2753) );
  MUX2X1 U3516 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n3096), .Y(n2757) );
  MUX2X1 U3517 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n3096), .Y(n2756) );
  MUX2X1 U3518 ( .B(n2755), .A(n2752), .S(n3081), .Y(n2766) );
  MUX2X1 U3519 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n3098), .Y(n2760) );
  MUX2X1 U3520 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n3098), .Y(n2759) );
  MUX2X1 U3521 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n3096), .Y(n2763) );
  MUX2X1 U3522 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n3096), .Y(n2762) );
  MUX2X1 U3523 ( .B(n2761), .A(n2758), .S(n3081), .Y(n2765) );
  MUX2X1 U3524 ( .B(n2764), .A(n2749), .S(N181), .Y(n2767) );
  MUX2X1 U3525 ( .B(\mem<62><3> ), .A(\mem<63><3> ), .S(n3097), .Y(n2771) );
  MUX2X1 U3526 ( .B(\mem<60><3> ), .A(\mem<61><3> ), .S(n3098), .Y(n2770) );
  MUX2X1 U3527 ( .B(\mem<58><3> ), .A(\mem<59><3> ), .S(n3099), .Y(n2774) );
  MUX2X1 U3528 ( .B(\mem<56><3> ), .A(\mem<57><3> ), .S(n3100), .Y(n2773) );
  MUX2X1 U3529 ( .B(n2772), .A(n2769), .S(n3081), .Y(n2783) );
  MUX2X1 U3530 ( .B(\mem<54><3> ), .A(\mem<55><3> ), .S(n3101), .Y(n2777) );
  MUX2X1 U3531 ( .B(\mem<52><3> ), .A(\mem<53><3> ), .S(n3101), .Y(n2776) );
  MUX2X1 U3532 ( .B(\mem<50><3> ), .A(\mem<51><3> ), .S(n3101), .Y(n2780) );
  MUX2X1 U3533 ( .B(\mem<48><3> ), .A(\mem<49><3> ), .S(n3101), .Y(n2779) );
  MUX2X1 U3534 ( .B(n2778), .A(n2775), .S(n3082), .Y(n2782) );
  MUX2X1 U3535 ( .B(\mem<46><3> ), .A(\mem<47><3> ), .S(n3101), .Y(n2786) );
  MUX2X1 U3536 ( .B(\mem<44><3> ), .A(\mem<45><3> ), .S(n3101), .Y(n2785) );
  MUX2X1 U3537 ( .B(\mem<42><3> ), .A(\mem<43><3> ), .S(n3101), .Y(n2789) );
  MUX2X1 U3538 ( .B(\mem<40><3> ), .A(\mem<41><3> ), .S(n3101), .Y(n2788) );
  MUX2X1 U3539 ( .B(n2787), .A(n2784), .S(n3082), .Y(n2798) );
  MUX2X1 U3540 ( .B(\mem<38><3> ), .A(\mem<39><3> ), .S(n3101), .Y(n2792) );
  MUX2X1 U3541 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n3101), .Y(n2791) );
  MUX2X1 U3542 ( .B(\mem<34><3> ), .A(\mem<35><3> ), .S(n3101), .Y(n2795) );
  MUX2X1 U3543 ( .B(\mem<32><3> ), .A(\mem<33><3> ), .S(n3101), .Y(n2794) );
  MUX2X1 U3544 ( .B(n2793), .A(n2790), .S(n3081), .Y(n2797) );
  MUX2X1 U3545 ( .B(n2796), .A(n2781), .S(N181), .Y(n2830) );
  MUX2X1 U3546 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n3102), .Y(n2801) );
  MUX2X1 U3547 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n3102), .Y(n2800) );
  MUX2X1 U3548 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n3102), .Y(n2804) );
  MUX2X1 U3549 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n3102), .Y(n2803) );
  MUX2X1 U3550 ( .B(n2802), .A(n2799), .S(n3081), .Y(n2813) );
  MUX2X1 U3551 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n3102), .Y(n2807) );
  MUX2X1 U3552 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n3102), .Y(n2806) );
  MUX2X1 U3553 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n3102), .Y(n2810) );
  MUX2X1 U3554 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n3102), .Y(n2809) );
  MUX2X1 U3555 ( .B(n2808), .A(n2805), .S(n3082), .Y(n2812) );
  MUX2X1 U3556 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n3102), .Y(n2816) );
  MUX2X1 U3557 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n3102), .Y(n2815) );
  MUX2X1 U3558 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n3102), .Y(n2819) );
  MUX2X1 U3559 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n3102), .Y(n2818) );
  MUX2X1 U3560 ( .B(n2817), .A(n2814), .S(n3081), .Y(n2828) );
  MUX2X1 U3561 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n3098), .Y(n2822) );
  MUX2X1 U3562 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n3096), .Y(n2821) );
  MUX2X1 U3563 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n3098), .Y(n2825) );
  MUX2X1 U3564 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n3096), .Y(n2824) );
  MUX2X1 U3565 ( .B(n2823), .A(n2820), .S(n3081), .Y(n2827) );
  MUX2X1 U3566 ( .B(n2826), .A(n2811), .S(N181), .Y(n2829) );
  MUX2X1 U3567 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n3096), .Y(n2833) );
  MUX2X1 U3568 ( .B(\mem<60><4> ), .A(\mem<61><4> ), .S(n3096), .Y(n2832) );
  MUX2X1 U3569 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n3098), .Y(n2836) );
  MUX2X1 U3570 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n3096), .Y(n2835) );
  MUX2X1 U3571 ( .B(n2834), .A(n2831), .S(n3081), .Y(n2845) );
  MUX2X1 U3572 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n3098), .Y(n2839) );
  MUX2X1 U3573 ( .B(\mem<52><4> ), .A(\mem<53><4> ), .S(n3096), .Y(n2838) );
  MUX2X1 U3574 ( .B(\mem<50><4> ), .A(\mem<51><4> ), .S(n3098), .Y(n2842) );
  MUX2X1 U3575 ( .B(\mem<48><4> ), .A(\mem<49><4> ), .S(n3098), .Y(n2841) );
  MUX2X1 U3576 ( .B(n2840), .A(n2837), .S(n3082), .Y(n2844) );
  MUX2X1 U3577 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n3103), .Y(n2848) );
  MUX2X1 U3578 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n3103), .Y(n2847) );
  MUX2X1 U3579 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n3103), .Y(n2851) );
  MUX2X1 U3580 ( .B(\mem<40><4> ), .A(\mem<41><4> ), .S(n3103), .Y(n2850) );
  MUX2X1 U3581 ( .B(n2849), .A(n2846), .S(n3081), .Y(n2860) );
  MUX2X1 U3582 ( .B(\mem<38><4> ), .A(\mem<39><4> ), .S(n3103), .Y(n2854) );
  MUX2X1 U3583 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n3103), .Y(n2853) );
  MUX2X1 U3584 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n3103), .Y(n2857) );
  MUX2X1 U3585 ( .B(\mem<32><4> ), .A(\mem<33><4> ), .S(n3103), .Y(n2856) );
  MUX2X1 U3586 ( .B(n2855), .A(n2852), .S(n3082), .Y(n2859) );
  MUX2X1 U3587 ( .B(n2858), .A(n2843), .S(N181), .Y(n2892) );
  MUX2X1 U3588 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n3103), .Y(n2863) );
  MUX2X1 U3589 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n3103), .Y(n2862) );
  MUX2X1 U3590 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n3103), .Y(n2866) );
  MUX2X1 U3591 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n3103), .Y(n2865) );
  MUX2X1 U3592 ( .B(n2864), .A(n2861), .S(n3080), .Y(n2875) );
  MUX2X1 U3593 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n3104), .Y(n2869) );
  MUX2X1 U3594 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n3104), .Y(n2868) );
  MUX2X1 U3595 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n3104), .Y(n2872) );
  MUX2X1 U3596 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n3104), .Y(n2871) );
  MUX2X1 U3597 ( .B(n2870), .A(n2867), .S(n3080), .Y(n2874) );
  MUX2X1 U3598 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n3104), .Y(n2878) );
  MUX2X1 U3599 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n3104), .Y(n2877) );
  MUX2X1 U3600 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n3104), .Y(n2881) );
  MUX2X1 U3601 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n3104), .Y(n2880) );
  MUX2X1 U3602 ( .B(n2879), .A(n2876), .S(n3080), .Y(n2890) );
  MUX2X1 U3603 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n3104), .Y(n2884) );
  MUX2X1 U3604 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n3104), .Y(n2883) );
  MUX2X1 U3605 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n3104), .Y(n2887) );
  MUX2X1 U3606 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n3104), .Y(n2886) );
  MUX2X1 U3607 ( .B(n2885), .A(n2882), .S(n3080), .Y(n2889) );
  MUX2X1 U3608 ( .B(n2888), .A(n2873), .S(N181), .Y(n2891) );
  MUX2X1 U3609 ( .B(\mem<62><5> ), .A(\mem<63><5> ), .S(n3105), .Y(n2895) );
  MUX2X1 U3610 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n3105), .Y(n2894) );
  MUX2X1 U3611 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n3105), .Y(n2898) );
  MUX2X1 U3612 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n3105), .Y(n2897) );
  MUX2X1 U3613 ( .B(n2896), .A(n2893), .S(n3080), .Y(n2907) );
  MUX2X1 U3614 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n3105), .Y(n2901) );
  MUX2X1 U3615 ( .B(\mem<52><5> ), .A(\mem<53><5> ), .S(n3105), .Y(n2900) );
  MUX2X1 U3616 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n3105), .Y(n2904) );
  MUX2X1 U3617 ( .B(\mem<48><5> ), .A(\mem<49><5> ), .S(n3105), .Y(n2903) );
  MUX2X1 U3618 ( .B(n2902), .A(n2899), .S(n3080), .Y(n2906) );
  MUX2X1 U3619 ( .B(\mem<46><5> ), .A(\mem<47><5> ), .S(n3105), .Y(n2910) );
  MUX2X1 U3620 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n3105), .Y(n2909) );
  MUX2X1 U3621 ( .B(\mem<42><5> ), .A(\mem<43><5> ), .S(n3105), .Y(n2913) );
  MUX2X1 U3622 ( .B(\mem<40><5> ), .A(\mem<41><5> ), .S(n3105), .Y(n2912) );
  MUX2X1 U3623 ( .B(n2911), .A(n2908), .S(n3080), .Y(n2922) );
  MUX2X1 U3624 ( .B(\mem<38><5> ), .A(\mem<39><5> ), .S(n3106), .Y(n2916) );
  MUX2X1 U3625 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n3106), .Y(n2915) );
  MUX2X1 U3626 ( .B(\mem<34><5> ), .A(\mem<35><5> ), .S(n3106), .Y(n2919) );
  MUX2X1 U3627 ( .B(\mem<32><5> ), .A(\mem<33><5> ), .S(n3106), .Y(n2918) );
  MUX2X1 U3628 ( .B(n2917), .A(n2914), .S(n3080), .Y(n2921) );
  MUX2X1 U3629 ( .B(n2920), .A(n2905), .S(N181), .Y(n2954) );
  MUX2X1 U3630 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n3106), .Y(n2925) );
  MUX2X1 U3631 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n3106), .Y(n2924) );
  MUX2X1 U3632 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n3106), .Y(n2928) );
  MUX2X1 U3633 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n3106), .Y(n2927) );
  MUX2X1 U3634 ( .B(n2926), .A(n2923), .S(n3080), .Y(n2937) );
  MUX2X1 U3635 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n3106), .Y(n2931) );
  MUX2X1 U3636 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n3106), .Y(n2930) );
  MUX2X1 U3637 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n3106), .Y(n2934) );
  MUX2X1 U3638 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n3106), .Y(n2933) );
  MUX2X1 U3639 ( .B(n2932), .A(n2929), .S(n3080), .Y(n2936) );
  MUX2X1 U3640 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n3107), .Y(n2940) );
  MUX2X1 U3641 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n3107), .Y(n2939) );
  MUX2X1 U3642 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n3107), .Y(n2943) );
  MUX2X1 U3643 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n3107), .Y(n2942) );
  MUX2X1 U3644 ( .B(n2941), .A(n2938), .S(n3080), .Y(n2952) );
  MUX2X1 U3645 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n3107), .Y(n2946) );
  MUX2X1 U3646 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n3107), .Y(n2945) );
  MUX2X1 U3647 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n3107), .Y(n2949) );
  MUX2X1 U3648 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n3107), .Y(n2948) );
  MUX2X1 U3649 ( .B(n2947), .A(n2944), .S(n3080), .Y(n2951) );
  MUX2X1 U3650 ( .B(n2950), .A(n2935), .S(N181), .Y(n2953) );
  MUX2X1 U3651 ( .B(\mem<62><6> ), .A(\mem<63><6> ), .S(n3107), .Y(n2957) );
  MUX2X1 U3652 ( .B(\mem<60><6> ), .A(\mem<61><6> ), .S(n3107), .Y(n2956) );
  MUX2X1 U3653 ( .B(\mem<58><6> ), .A(\mem<59><6> ), .S(n3107), .Y(n2960) );
  MUX2X1 U3654 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n3107), .Y(n2959) );
  MUX2X1 U3655 ( .B(n2958), .A(n2955), .S(n3079), .Y(n2969) );
  MUX2X1 U3656 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n3108), .Y(n2963) );
  MUX2X1 U3657 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n3108), .Y(n2962) );
  MUX2X1 U3658 ( .B(\mem<50><6> ), .A(\mem<51><6> ), .S(n3108), .Y(n2966) );
  MUX2X1 U3659 ( .B(\mem<48><6> ), .A(\mem<49><6> ), .S(n3108), .Y(n2965) );
  MUX2X1 U3660 ( .B(n2964), .A(n2961), .S(n3079), .Y(n2968) );
  MUX2X1 U3661 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n3108), .Y(n2972) );
  MUX2X1 U3662 ( .B(\mem<44><6> ), .A(\mem<45><6> ), .S(n3108), .Y(n2971) );
  MUX2X1 U3663 ( .B(\mem<42><6> ), .A(\mem<43><6> ), .S(n3108), .Y(n2975) );
  MUX2X1 U3664 ( .B(\mem<40><6> ), .A(\mem<41><6> ), .S(n3108), .Y(n2974) );
  MUX2X1 U3665 ( .B(n2973), .A(n2970), .S(n3079), .Y(n2984) );
  MUX2X1 U3666 ( .B(\mem<38><6> ), .A(\mem<39><6> ), .S(n3108), .Y(n2978) );
  MUX2X1 U3667 ( .B(\mem<36><6> ), .A(\mem<37><6> ), .S(n3108), .Y(n2977) );
  MUX2X1 U3668 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n3108), .Y(n2981) );
  MUX2X1 U3669 ( .B(\mem<32><6> ), .A(\mem<33><6> ), .S(n3108), .Y(n2980) );
  MUX2X1 U3670 ( .B(n2979), .A(n2976), .S(n3079), .Y(n2983) );
  MUX2X1 U3671 ( .B(n2982), .A(n2967), .S(N181), .Y(n3016) );
  MUX2X1 U3672 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n3109), .Y(n2987) );
  MUX2X1 U3673 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n3109), .Y(n2986) );
  MUX2X1 U3674 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n3109), .Y(n2990) );
  MUX2X1 U3675 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n3109), .Y(n2989) );
  MUX2X1 U3676 ( .B(n2988), .A(n2985), .S(n3079), .Y(n2999) );
  MUX2X1 U3677 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n3109), .Y(n2993) );
  MUX2X1 U3678 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n3109), .Y(n2992) );
  MUX2X1 U3679 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n3109), .Y(n2996) );
  MUX2X1 U3680 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n3109), .Y(n2995) );
  MUX2X1 U3681 ( .B(n2994), .A(n2991), .S(n3079), .Y(n2998) );
  MUX2X1 U3682 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n3109), .Y(n3002) );
  MUX2X1 U3683 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n3109), .Y(n3001) );
  MUX2X1 U3684 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n3109), .Y(n3005) );
  MUX2X1 U3685 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n3109), .Y(n3004) );
  MUX2X1 U3686 ( .B(n3003), .A(n3000), .S(n3079), .Y(n3014) );
  MUX2X1 U3687 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n3110), .Y(n3008) );
  MUX2X1 U3688 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n3110), .Y(n3007) );
  MUX2X1 U3689 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n3110), .Y(n3011) );
  MUX2X1 U3690 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n3110), .Y(n3010) );
  MUX2X1 U3691 ( .B(n3009), .A(n3006), .S(n3079), .Y(n3013) );
  MUX2X1 U3692 ( .B(n3012), .A(n2997), .S(N181), .Y(n3015) );
  MUX2X1 U3693 ( .B(\mem<62><7> ), .A(\mem<63><7> ), .S(n3110), .Y(n3019) );
  MUX2X1 U3694 ( .B(\mem<60><7> ), .A(\mem<61><7> ), .S(n3110), .Y(n3018) );
  MUX2X1 U3695 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n3110), .Y(n3022) );
  MUX2X1 U3696 ( .B(\mem<56><7> ), .A(\mem<57><7> ), .S(n3110), .Y(n3021) );
  MUX2X1 U3697 ( .B(n3020), .A(n3017), .S(n3079), .Y(n3031) );
  MUX2X1 U3698 ( .B(\mem<54><7> ), .A(\mem<55><7> ), .S(n3110), .Y(n3025) );
  MUX2X1 U3699 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n3110), .Y(n3024) );
  MUX2X1 U3700 ( .B(\mem<50><7> ), .A(\mem<51><7> ), .S(n3110), .Y(n3028) );
  MUX2X1 U3701 ( .B(\mem<48><7> ), .A(\mem<49><7> ), .S(n3110), .Y(n3027) );
  MUX2X1 U3702 ( .B(n3026), .A(n3023), .S(n3079), .Y(n3030) );
  MUX2X1 U3703 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n3111), .Y(n3034) );
  MUX2X1 U3704 ( .B(\mem<44><7> ), .A(\mem<45><7> ), .S(n3111), .Y(n3033) );
  MUX2X1 U3705 ( .B(\mem<42><7> ), .A(\mem<43><7> ), .S(n3111), .Y(n3037) );
  MUX2X1 U3706 ( .B(\mem<40><7> ), .A(\mem<41><7> ), .S(n3111), .Y(n3036) );
  MUX2X1 U3707 ( .B(n3035), .A(n3032), .S(n3079), .Y(n3046) );
  MUX2X1 U3708 ( .B(\mem<38><7> ), .A(\mem<39><7> ), .S(n3111), .Y(n3040) );
  MUX2X1 U3709 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n3111), .Y(n3039) );
  MUX2X1 U3710 ( .B(\mem<34><7> ), .A(\mem<35><7> ), .S(n3111), .Y(n3043) );
  MUX2X1 U3711 ( .B(\mem<32><7> ), .A(\mem<33><7> ), .S(n3111), .Y(n3042) );
  MUX2X1 U3712 ( .B(n3041), .A(n3038), .S(n3079), .Y(n3045) );
  MUX2X1 U3713 ( .B(n3044), .A(n3029), .S(N181), .Y(n3078) );
  MUX2X1 U3714 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n3111), .Y(n3049) );
  MUX2X1 U3715 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n3111), .Y(n3048) );
  MUX2X1 U3716 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n3111), .Y(n3052) );
  MUX2X1 U3717 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n3111), .Y(n3051) );
  MUX2X1 U3718 ( .B(n3050), .A(n3047), .S(n3080), .Y(n3061) );
  MUX2X1 U3719 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n3095), .Y(n3055) );
  MUX2X1 U3720 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n3094), .Y(n3054) );
  MUX2X1 U3721 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n3094), .Y(n3058) );
  MUX2X1 U3722 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n3094), .Y(n3057) );
  MUX2X1 U3723 ( .B(n3056), .A(n3053), .S(n3079), .Y(n3060) );
  MUX2X1 U3724 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n3095), .Y(n3064) );
  MUX2X1 U3725 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n3095), .Y(n3063) );
  MUX2X1 U3726 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n3094), .Y(n3067) );
  MUX2X1 U3727 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n3095), .Y(n3066) );
  MUX2X1 U3728 ( .B(n3065), .A(n3062), .S(n3080), .Y(n3076) );
  MUX2X1 U3729 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n3094), .Y(n3070) );
  MUX2X1 U3730 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n3095), .Y(n3069) );
  MUX2X1 U3731 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n3095), .Y(n3073) );
  MUX2X1 U3732 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n3095), .Y(n3072) );
  MUX2X1 U3733 ( .B(n3071), .A(n3068), .S(n3079), .Y(n3075) );
  MUX2X1 U3734 ( .B(n3074), .A(n3059), .S(N181), .Y(n3077) );
endmodule


module cla16_2 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n5,
         n6, n7, n8, n1, n2, n4, n9, n10;

  AOI21X1 U5 ( .A(\P<3> ), .B(n4), .C(\G<3> ), .Y(n5) );
  AOI21X1 U6 ( .A(\P<2> ), .B(n9), .C(\G<2> ), .Y(n6) );
  AOI21X1 U7 ( .A(\P<1> ), .B(n10), .C(\G<1> ), .Y(n7) );
  AOI21X1 U8 ( .A(\P<0> ), .B(Cin), .C(\G<0> ), .Y(n8) );
  cla4_11 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_10 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n10), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_9 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n9), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_8 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n4), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  BUFX2 U1 ( .A(n7), .Y(n1) );
  INVX1 U2 ( .A(n6), .Y(n4) );
  INVX1 U3 ( .A(n8), .Y(n10) );
  BUFX2 U4 ( .A(n5), .Y(n2) );
  INVX1 U9 ( .A(n2), .Y(Cout) );
  INVX2 U10 ( .A(n1), .Y(n9) );
endmodule


module dff_355 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_356 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_357 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_358 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_359 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_360 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_361 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_362 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_363 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_364 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_365 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_366 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_367 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_368 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_369 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_370 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_339 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_340 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_341 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_342 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_343 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_344 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_345 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_346 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_347 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_348 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_349 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_350 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_351 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_352 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_353 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_354 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_371 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module rf_bypass ( .read1data({\read1data<15> , \read1data<14> , 
        \read1data<13> , \read1data<12> , \read1data<11> , \read1data<10> , 
        \read1data<9> , \read1data<8> , \read1data<7> , \read1data<6> , 
        \read1data<5> , \read1data<4> , \read1data<3> , \read1data<2> , 
        \read1data<1> , \read1data<0> }), .read2data({\read2data<15> , 
        \read2data<14> , \read2data<13> , \read2data<12> , \read2data<11> , 
        \read2data<10> , \read2data<9> , \read2data<8> , \read2data<7> , 
        \read2data<6> , \read2data<5> , \read2data<4> , \read2data<3> , 
        \read2data<2> , \read2data<1> , \read2data<0> }), err, clk, rst, 
    .read1regsel({\read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), 
    .read2regsel({\read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), 
    .writeregsel({\writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), 
    .writedata({\writedata<15> , \writedata<14> , \writedata<13> , 
        \writedata<12> , \writedata<11> , \writedata<10> , \writedata<9> , 
        \writedata<8> , \writedata<7> , \writedata<6> , \writedata<5> , 
        \writedata<4> , \writedata<3> , \writedata<2> , \writedata<1> , 
        \writedata<0> }), write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   \rf_r1_out<15> , \rf_r1_out<14> , \rf_r1_out<13> , \rf_r1_out<12> ,
         \rf_r1_out<11> , \rf_r1_out<10> , \rf_r1_out<9> , \rf_r1_out<8> ,
         \rf_r1_out<7> , \rf_r1_out<6> , \rf_r1_out<5> , \rf_r1_out<4> ,
         \rf_r1_out<3> , \rf_r1_out<2> , \rf_r1_out<1> , \rf_r1_out<0> ,
         \rf_r2_out<15> , \rf_r2_out<14> , \rf_r2_out<13> , \rf_r2_out<12> ,
         \rf_r2_out<11> , \rf_r2_out<10> , \rf_r2_out<9> , \rf_r2_out<8> ,
         \rf_r2_out<7> , \rf_r2_out<6> , \rf_r2_out<5> , \rf_r2_out<4> ,
         \rf_r2_out<3> , \rf_r2_out<2> , \rf_r2_out<1> , \rf_r2_out<0> , n19,
         n36, n37, n38, n39, n40, n57, n58, n59, n60, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;
  assign err = 1'b0;

  OAI21X1 U18 ( .A(n76), .B(n91), .C(n74), .Y(\read2data<9> ) );
  OAI21X1 U20 ( .A(n76), .B(n90), .C(n72), .Y(\read2data<8> ) );
  OAI21X1 U22 ( .A(n76), .B(n89), .C(n70), .Y(\read2data<7> ) );
  OAI21X1 U24 ( .A(n76), .B(n88), .C(n68), .Y(\read2data<6> ) );
  OAI21X1 U26 ( .A(n76), .B(n87), .C(n66), .Y(\read2data<5> ) );
  OAI21X1 U28 ( .A(n76), .B(n86), .C(n64), .Y(\read2data<4> ) );
  OAI21X1 U30 ( .A(n76), .B(n85), .C(n62), .Y(\read2data<3> ) );
  OAI21X1 U32 ( .A(n76), .B(n84), .C(n56), .Y(\read2data<2> ) );
  OAI21X1 U34 ( .A(n76), .B(n83), .C(n54), .Y(\read2data<1> ) );
  OAI21X1 U36 ( .A(n76), .B(n97), .C(n52), .Y(\read2data<15> ) );
  OAI21X1 U38 ( .A(n76), .B(n96), .C(n50), .Y(\read2data<14> ) );
  OAI21X1 U40 ( .A(n76), .B(n95), .C(n48), .Y(\read2data<13> ) );
  OAI21X1 U42 ( .A(n76), .B(n94), .C(n46), .Y(\read2data<12> ) );
  OAI21X1 U44 ( .A(n76), .B(n93), .C(n44), .Y(\read2data<11> ) );
  OAI21X1 U46 ( .A(n76), .B(n92), .C(n42), .Y(\read2data<10> ) );
  OAI21X1 U48 ( .A(n76), .B(n82), .C(n35), .Y(\read2data<0> ) );
  NAND3X1 U50 ( .A(n36), .B(n37), .C(n38), .Y(n19) );
  NOR2X1 U51 ( .A(n81), .B(n39), .Y(n38) );
  XOR2X1 U52 ( .A(n79), .B(\read2regsel<2> ), .Y(n39) );
  XNOR2X1 U53 ( .A(n77), .B(\read2regsel<1> ), .Y(n37) );
  XNOR2X1 U54 ( .A(\writeregsel<0> ), .B(\read2regsel<0> ), .Y(n36) );
  OAI21X1 U55 ( .A(n91), .B(n75), .C(n33), .Y(\read1data<9> ) );
  OAI21X1 U57 ( .A(n90), .B(n75), .C(n31), .Y(\read1data<8> ) );
  OAI21X1 U59 ( .A(n89), .B(n75), .C(n29), .Y(\read1data<7> ) );
  OAI21X1 U61 ( .A(n88), .B(n75), .C(n27), .Y(\read1data<6> ) );
  OAI21X1 U63 ( .A(n87), .B(n75), .C(n25), .Y(\read1data<5> ) );
  OAI21X1 U65 ( .A(n86), .B(n75), .C(n23), .Y(\read1data<4> ) );
  OAI21X1 U67 ( .A(n85), .B(n75), .C(n21), .Y(\read1data<3> ) );
  OAI21X1 U69 ( .A(n84), .B(n75), .C(n18), .Y(\read1data<2> ) );
  OAI21X1 U71 ( .A(n83), .B(n75), .C(n16), .Y(\read1data<1> ) );
  OAI21X1 U73 ( .A(n97), .B(n75), .C(n14), .Y(\read1data<15> ) );
  OAI21X1 U75 ( .A(n96), .B(n75), .C(n12), .Y(\read1data<14> ) );
  OAI21X1 U77 ( .A(n95), .B(n75), .C(n10), .Y(\read1data<13> ) );
  OAI21X1 U79 ( .A(n94), .B(n75), .C(n8), .Y(\read1data<12> ) );
  OAI21X1 U81 ( .A(n93), .B(n75), .C(n6), .Y(\read1data<11> ) );
  OAI21X1 U83 ( .A(n92), .B(n75), .C(n4), .Y(\read1data<10> ) );
  OAI21X1 U85 ( .A(n82), .B(n75), .C(n2), .Y(\read1data<0> ) );
  NAND3X1 U87 ( .A(n57), .B(n58), .C(n59), .Y(n40) );
  NOR2X1 U88 ( .A(n81), .B(n60), .Y(n59) );
  XOR2X1 U89 ( .A(n79), .B(\read1regsel<2> ), .Y(n60) );
  XNOR2X1 U90 ( .A(n77), .B(\read1regsel<1> ), .Y(n58) );
  XNOR2X1 U91 ( .A(\writeregsel<0> ), .B(\read1regsel<0> ), .Y(n57) );
  rf regfile ( .read1data({\rf_r1_out<15> , \rf_r1_out<14> , \rf_r1_out<13> , 
        \rf_r1_out<12> , \rf_r1_out<11> , \rf_r1_out<10> , \rf_r1_out<9> , 
        \rf_r1_out<8> , \rf_r1_out<7> , \rf_r1_out<6> , \rf_r1_out<5> , 
        \rf_r1_out<4> , \rf_r1_out<3> , \rf_r1_out<2> , \rf_r1_out<1> , 
        \rf_r1_out<0> }), .read2data({\rf_r2_out<15> , \rf_r2_out<14> , 
        \rf_r2_out<13> , \rf_r2_out<12> , \rf_r2_out<11> , \rf_r2_out<10> , 
        \rf_r2_out<9> , \rf_r2_out<8> , \rf_r2_out<7> , \rf_r2_out<6> , 
        \rf_r2_out<5> , \rf_r2_out<4> , \rf_r2_out<3> , \rf_r2_out<2> , 
        \rf_r2_out<1> , \rf_r2_out<0> }), .err(), .clk(clk), .rst(rst), 
        .read1regsel({\read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), 
        .read2regsel({\read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), 
        .writeregsel({n79, n77, \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        .write(write) );
  INVX1 U1 ( .A(\writedata<2> ), .Y(n84) );
  INVX1 U2 ( .A(\writedata<10> ), .Y(n92) );
  INVX1 U3 ( .A(write), .Y(n81) );
  INVX1 U4 ( .A(n80), .Y(n79) );
  INVX1 U5 ( .A(\writeregsel<2> ), .Y(n80) );
  INVX1 U6 ( .A(n78), .Y(n77) );
  INVX1 U7 ( .A(\writeregsel<1> ), .Y(n78) );
  INVX1 U8 ( .A(\writedata<0> ), .Y(n82) );
  INVX1 U9 ( .A(\writedata<1> ), .Y(n83) );
  INVX1 U10 ( .A(\writedata<3> ), .Y(n85) );
  INVX1 U11 ( .A(\writedata<4> ), .Y(n86) );
  INVX1 U12 ( .A(\writedata<5> ), .Y(n87) );
  INVX1 U13 ( .A(\writedata<6> ), .Y(n88) );
  INVX1 U14 ( .A(\writedata<7> ), .Y(n89) );
  INVX1 U15 ( .A(\writedata<8> ), .Y(n90) );
  INVX1 U16 ( .A(\writedata<9> ), .Y(n91) );
  INVX1 U17 ( .A(\writedata<11> ), .Y(n93) );
  INVX1 U19 ( .A(\writedata<12> ), .Y(n94) );
  INVX1 U21 ( .A(\writedata<13> ), .Y(n95) );
  INVX1 U23 ( .A(\writedata<14> ), .Y(n96) );
  INVX1 U25 ( .A(\writedata<15> ), .Y(n97) );
  AND2X1 U27 ( .A(\rf_r1_out<0> ), .B(n75), .Y(n1) );
  INVX1 U29 ( .A(n1), .Y(n2) );
  AND2X1 U31 ( .A(\rf_r1_out<10> ), .B(n75), .Y(n3) );
  INVX1 U33 ( .A(n3), .Y(n4) );
  AND2X1 U35 ( .A(\rf_r1_out<11> ), .B(n75), .Y(n5) );
  INVX1 U37 ( .A(n5), .Y(n6) );
  AND2X1 U39 ( .A(\rf_r1_out<12> ), .B(n75), .Y(n7) );
  INVX1 U41 ( .A(n7), .Y(n8) );
  AND2X1 U43 ( .A(\rf_r1_out<13> ), .B(n75), .Y(n9) );
  INVX1 U45 ( .A(n9), .Y(n10) );
  AND2X1 U47 ( .A(\rf_r1_out<14> ), .B(n75), .Y(n11) );
  INVX1 U49 ( .A(n11), .Y(n12) );
  AND2X1 U56 ( .A(\rf_r1_out<15> ), .B(n75), .Y(n13) );
  INVX1 U58 ( .A(n13), .Y(n14) );
  AND2X1 U60 ( .A(\rf_r1_out<1> ), .B(n75), .Y(n15) );
  INVX1 U62 ( .A(n15), .Y(n16) );
  AND2X1 U64 ( .A(\rf_r1_out<2> ), .B(n75), .Y(n17) );
  INVX1 U66 ( .A(n17), .Y(n18) );
  AND2X1 U68 ( .A(\rf_r1_out<3> ), .B(n75), .Y(n20) );
  INVX1 U70 ( .A(n20), .Y(n21) );
  AND2X1 U72 ( .A(\rf_r1_out<4> ), .B(n75), .Y(n22) );
  INVX1 U74 ( .A(n22), .Y(n23) );
  AND2X1 U76 ( .A(\rf_r1_out<5> ), .B(n75), .Y(n24) );
  INVX1 U78 ( .A(n24), .Y(n25) );
  AND2X1 U80 ( .A(\rf_r1_out<6> ), .B(n75), .Y(n26) );
  INVX1 U82 ( .A(n26), .Y(n27) );
  AND2X1 U84 ( .A(\rf_r1_out<7> ), .B(n75), .Y(n28) );
  INVX1 U86 ( .A(n28), .Y(n29) );
  AND2X1 U92 ( .A(\rf_r1_out<8> ), .B(n75), .Y(n30) );
  INVX1 U93 ( .A(n30), .Y(n31) );
  AND2X1 U94 ( .A(\rf_r1_out<9> ), .B(n75), .Y(n32) );
  INVX1 U95 ( .A(n32), .Y(n33) );
  AND2X1 U96 ( .A(\rf_r2_out<0> ), .B(n76), .Y(n34) );
  INVX1 U97 ( .A(n34), .Y(n35) );
  AND2X1 U98 ( .A(\rf_r2_out<10> ), .B(n76), .Y(n41) );
  INVX1 U99 ( .A(n41), .Y(n42) );
  AND2X1 U100 ( .A(\rf_r2_out<11> ), .B(n76), .Y(n43) );
  INVX1 U101 ( .A(n43), .Y(n44) );
  AND2X1 U102 ( .A(\rf_r2_out<12> ), .B(n76), .Y(n45) );
  INVX1 U103 ( .A(n45), .Y(n46) );
  AND2X1 U104 ( .A(\rf_r2_out<13> ), .B(n76), .Y(n47) );
  INVX1 U105 ( .A(n47), .Y(n48) );
  AND2X1 U106 ( .A(\rf_r2_out<14> ), .B(n76), .Y(n49) );
  INVX1 U107 ( .A(n49), .Y(n50) );
  AND2X1 U108 ( .A(\rf_r2_out<15> ), .B(n76), .Y(n51) );
  INVX1 U109 ( .A(n51), .Y(n52) );
  AND2X1 U110 ( .A(\rf_r2_out<1> ), .B(n76), .Y(n53) );
  INVX1 U111 ( .A(n53), .Y(n54) );
  AND2X1 U112 ( .A(\rf_r2_out<2> ), .B(n76), .Y(n55) );
  INVX1 U113 ( .A(n55), .Y(n56) );
  AND2X1 U114 ( .A(\rf_r2_out<3> ), .B(n76), .Y(n61) );
  INVX1 U115 ( .A(n61), .Y(n62) );
  AND2X1 U116 ( .A(\rf_r2_out<4> ), .B(n76), .Y(n63) );
  INVX1 U117 ( .A(n63), .Y(n64) );
  AND2X1 U118 ( .A(\rf_r2_out<5> ), .B(n76), .Y(n65) );
  INVX1 U119 ( .A(n65), .Y(n66) );
  AND2X1 U120 ( .A(\rf_r2_out<6> ), .B(n76), .Y(n67) );
  INVX1 U121 ( .A(n67), .Y(n68) );
  AND2X1 U122 ( .A(\rf_r2_out<7> ), .B(n76), .Y(n69) );
  INVX1 U123 ( .A(n69), .Y(n70) );
  AND2X1 U124 ( .A(\rf_r2_out<8> ), .B(n76), .Y(n71) );
  INVX1 U125 ( .A(n71), .Y(n72) );
  AND2X1 U126 ( .A(\rf_r2_out<9> ), .B(n76), .Y(n73) );
  INVX1 U127 ( .A(n73), .Y(n74) );
  BUFX2 U128 ( .A(n40), .Y(n75) );
  BUFX2 U129 ( .A(n19), .Y(n76) );
endmodule


module control_unit ( .opcode({\opcode<4> , \opcode<3> , \opcode<2> , 
        \opcode<1> , \opcode<0> }), .func({\func<1> , \func<0> }), .aluop({
        \aluop<2> , \aluop<1> , \aluop<0> }), alusrc, branch, jump, i1, i2, r, 
        jumpreg, set, btr, regwrite, memwrite, memread, memtoreg, invA, invB, 
        cin, excp, zeroext, halt, slbi, link, lbi, stu, rti );
  input \opcode<4> , \opcode<3> , \opcode<2> , \opcode<1> , \opcode<0> ,
         \func<1> , \func<0> ;
  output \aluop<2> , \aluop<1> , \aluop<0> , alusrc, branch, jump, i1, i2, r,
         jumpreg, set, btr, regwrite, memwrite, memread, memtoreg, invA, invB,
         cin, excp, zeroext, halt, slbi, link, lbi, stu, rti;
  wire   n81, N34, N55, n22, n23, n24, n25, n28, n29, n32, n33, n35, n36, n38,
         n41, n43, n44, n46, n47, n48, n49, n50, n51, n54, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20, n21,
         n30, n34, n39, n40, n42, n45, n53, n57, n58, n59, n61, n62, n63, n64,
         n66, n67, n68, n70, n71, n73, n74, n75, n76, n77, n78, n79, n80;

  AND2X2 U1 ( .A(n70), .B(n24), .Y(halt) );
  AND2X2 U2 ( .A(\opcode<1> ), .B(jump), .Y(link) );
  AND2X2 U3 ( .A(\opcode<0> ), .B(jump), .Y(jumpreg) );
  AND2X2 U4 ( .A(\opcode<2> ), .B(n24), .Y(jump) );
  AND2X2 U5 ( .A(n38), .B(n24), .Y(excp) );
  AND2X2 U6 ( .A(n47), .B(n48), .Y(n46) );
  OAI21X1 U26 ( .A(\opcode<4> ), .B(n15), .C(n64), .Y(zeroext) );
  NOR3X1 U27 ( .A(n71), .B(n75), .C(n22), .Y(stu) );
  NOR3X1 U28 ( .A(n23), .B(\opcode<2> ), .C(n75), .Y(rti) );
  NAND2X1 U29 ( .A(n24), .B(\opcode<0> ), .Y(n23) );
  NAND3X1 U32 ( .A(\opcode<1> ), .B(n78), .C(\opcode<2> ), .Y(n25) );
  OAI21X1 U36 ( .A(n73), .B(n17), .C(n35), .Y(invB) );
  NAND3X1 U37 ( .A(n62), .B(n36), .C(n64), .Y(i2) );
  AOI21X1 U38 ( .A(n7), .B(\opcode<0> ), .C(branch), .Y(n36) );
  OAI21X1 U40 ( .A(n38), .B(n13), .C(n4), .Y(i1) );
  NOR2X1 U42 ( .A(\opcode<3> ), .B(\opcode<4> ), .Y(n24) );
  OAI21X1 U43 ( .A(n73), .B(n17), .C(n67), .Y(cin) );
  OAI21X1 U44 ( .A(n41), .B(n6), .C(n43), .Y(invA) );
  NAND3X1 U45 ( .A(n1), .B(n80), .C(n74), .Y(n43) );
  NAND3X1 U47 ( .A(n14), .B(n68), .C(\opcode<4> ), .Y(n41) );
  NOR3X1 U48 ( .A(n33), .B(n2), .C(n80), .Y(btr) );
  NOR2X1 U49 ( .A(n8), .B(n78), .Y(branch) );
  OAI21X1 U52 ( .A(n70), .B(n80), .C(\opcode<3> ), .Y(n44) );
  NAND3X1 U53 ( .A(n75), .B(n76), .C(n71), .Y(n28) );
  NAND3X1 U54 ( .A(n35), .B(n64), .C(n46), .Y(N55) );
  NAND3X1 U55 ( .A(\opcode<0> ), .B(n77), .C(\opcode<2> ), .Y(n48) );
  NAND3X1 U56 ( .A(n38), .B(\opcode<4> ), .C(\func<0> ), .Y(n47) );
  NOR3X1 U58 ( .A(\opcode<0> ), .B(\opcode<2> ), .C(n75), .Y(n38) );
  NAND3X1 U59 ( .A(n14), .B(n49), .C(\opcode<0> ), .Y(n35) );
  OAI21X1 U60 ( .A(n66), .B(n68), .C(\opcode<4> ), .Y(n49) );
  NAND3X1 U61 ( .A(n50), .B(n51), .C(n58), .Y(N34) );
  NOR2X1 U65 ( .A(\opcode<1> ), .B(\opcode<0> ), .Y(n29) );
  NAND3X1 U66 ( .A(n77), .B(\opcode<1> ), .C(\opcode<2> ), .Y(n51) );
  OAI21X1 U67 ( .A(\func<1> ), .B(n80), .C(n14), .Y(n50) );
  NAND3X1 U72 ( .A(n32), .B(n76), .C(\opcode<4> ), .Y(n54) );
  OAI21X1 U73 ( .A(\opcode<0> ), .B(n75), .C(n33), .Y(n32) );
  NAND2X1 U74 ( .A(\opcode<0> ), .B(n75), .Y(n33) );
  NAND2X1 U75 ( .A(n77), .B(n76), .Y(n22) );
  INVX1 U7 ( .A(\func<1> ), .Y(n68) );
  INVX1 U8 ( .A(invA), .Y(n67) );
  INVX1 U9 ( .A(n62), .Y(lbi) );
  INVX1 U10 ( .A(n64), .Y(slbi) );
  INVX1 U11 ( .A(\func<0> ), .Y(n66) );
  INVX1 U12 ( .A(n32), .Y(n73) );
  AND2X2 U13 ( .A(\opcode<3> ), .B(n76), .Y(n1) );
  INVX1 U14 ( .A(n1), .Y(n2) );
  INVX2 U15 ( .A(\opcode<2> ), .Y(n76) );
  AND2X2 U16 ( .A(n1), .B(n80), .Y(n3) );
  INVX1 U17 ( .A(n3), .Y(n4) );
  AND2X2 U18 ( .A(\func<0> ), .B(\opcode<0> ), .Y(n5) );
  INVX1 U19 ( .A(n5), .Y(n6) );
  AND2X2 U20 ( .A(\opcode<2> ), .B(n80), .Y(n7) );
  INVX1 U21 ( .A(n7), .Y(n8) );
  AND2X2 U22 ( .A(\opcode<4> ), .B(\opcode<3> ), .Y(n9) );
  INVX1 U23 ( .A(n9), .Y(n10) );
  INVX1 U24 ( .A(n9), .Y(n11) );
  AND2X2 U25 ( .A(\opcode<4> ), .B(n78), .Y(n12) );
  INVX1 U30 ( .A(n12), .Y(n13) );
  AND2X2 U31 ( .A(\opcode<1> ), .B(n1), .Y(n14) );
  INVX1 U33 ( .A(n14), .Y(n15) );
  AND2X2 U34 ( .A(\opcode<2> ), .B(n79), .Y(set) );
  INVX1 U35 ( .A(set), .Y(n17) );
  AND2X2 U39 ( .A(\opcode<3> ), .B(n54), .Y(n18) );
  AND2X2 U41 ( .A(\opcode<2> ), .B(n78), .Y(n19) );
  AND2X2 U46 ( .A(\opcode<4> ), .B(n28), .Y(n20) );
  INVX1 U50 ( .A(n28), .Y(n70) );
  INVX1 U51 ( .A(\opcode<4> ), .Y(n80) );
  INVX1 U57 ( .A(\opcode<3> ), .Y(n78) );
  INVX1 U62 ( .A(n81), .Y(n21) );
  INVX2 U63 ( .A(n21), .Y(r) );
  OR2X1 U64 ( .A(n40), .B(n30), .Y(alusrc) );
  OR2X1 U68 ( .A(n19), .B(n77), .Y(n30) );
  OR2X1 U69 ( .A(n42), .B(n34), .Y(regwrite) );
  OR2X1 U70 ( .A(n20), .B(n1), .Y(n34) );
  OR2X1 U71 ( .A(n7), .B(n39), .Y(\aluop<2> ) );
  OR2X1 U76 ( .A(n18), .B(n53), .Y(n39) );
  INVX1 U77 ( .A(n44), .Y(n40) );
  INVX1 U78 ( .A(n25), .Y(n42) );
  OR2X2 U79 ( .A(n32), .B(n22), .Y(n45) );
  INVX1 U80 ( .A(n45), .Y(memwrite) );
  INVX1 U81 ( .A(n33), .Y(n74) );
  INVX1 U82 ( .A(n22), .Y(n53) );
  BUFX2 U83 ( .A(N34), .Y(\aluop<1> ) );
  BUFX2 U84 ( .A(N55), .Y(\aluop<0> ) );
  AND2X2 U85 ( .A(n29), .B(set), .Y(n57) );
  INVX1 U86 ( .A(n57), .Y(n58) );
  OR2X2 U87 ( .A(n33), .B(n22), .Y(n59) );
  INVX1 U88 ( .A(n59), .Y(memtoreg) );
  AND2X1 U89 ( .A(n70), .B(n79), .Y(n61) );
  INVX1 U90 ( .A(n61), .Y(n62) );
  INVX1 U91 ( .A(n11), .Y(n79) );
  AND2X1 U92 ( .A(n77), .B(n38), .Y(n63) );
  INVX1 U93 ( .A(n63), .Y(n64) );
  INVX1 U94 ( .A(n13), .Y(n77) );
  AOI21X1 U95 ( .A(n76), .B(n29), .C(n10), .Y(n81) );
  BUFX2 U96 ( .A(memtoreg), .Y(memread) );
  INVX2 U97 ( .A(\opcode<0> ), .Y(n71) );
  INVX2 U98 ( .A(\opcode<1> ), .Y(n75) );
endmodule


module dff_338 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_304 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_305 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_306 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_307 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_308 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_309 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_310 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_311 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_312 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_313 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_314 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_315 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_316 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_317 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_318 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_319 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_337 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_336 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_335 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_301 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_302 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_303 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_285 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_286 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_287 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_288 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_289 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_290 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_291 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_292 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_293 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_294 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_295 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_296 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_297 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_298 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_299 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_300 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_334 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_282 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_283 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_284 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_279 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_280 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_281 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_276 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_277 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_278 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_264 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_265 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_266 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_267 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_268 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_269 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_270 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_271 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_272 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_273 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_274 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_275 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_333 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_332 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_331 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_330 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_329 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_328 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_327 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_326 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_325 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_324 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_323 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_322 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_321 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_320 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module alu ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , 
        \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> 
        }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , 
        \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> 
        }), Cin, .Op({\Op<2> , \Op<1> , \Op<0> }), invA, invB, sign, .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }), Ofl, Z, Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<2> , \Op<1> , \Op<0> , invA, invB, sign;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Ofl, Z, Cout;
  wire   \A_real<15> , \A_real<14> , \A_real<13> , \A_real<12> , \A_real<11> ,
         \A_real<10> , \A_real<9> , \A_real<8> , \A_real<7> , \A_real<6> ,
         \A_real<5> , \A_real<4> , \A_real<3> , \A_real<2> , \A_real<1> ,
         \A_real<0> , \B_real<15> , \B_real<14> , \B_real<13> , \B_real<12> ,
         \B_real<11> , \B_real<10> , \B_real<9> , \B_real<8> , \B_real<7> ,
         \B_real<6> , \B_real<5> , \B_real<4> , \B_real<3> , \B_real<2> ,
         \B_real<1> , \B_real<0> , \op0_out<15> , \op0_out<14> , \op0_out<13> ,
         \op0_out<12> , \op0_out<11> , \op0_out<10> , \op0_out<9> ,
         \op0_out<8> , \op0_out<7> , \op0_out<6> , \op0_out<5> , \op0_out<4> ,
         \op0_out<3> , \op0_out<2> , \op0_out<1> , \op0_out<0> , \op1_out<15> ,
         \op1_out<14> , \op1_out<13> , \op1_out<12> , \op1_out<11> ,
         \op1_out<10> , \op1_out<9> , \op1_out<8> , \op1_out<7> , \op1_out<6> ,
         \op1_out<5> , \op1_out<4> , \op1_out<3> , \op1_out<2> , \op1_out<1> ,
         \op1_out<0> , \op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> ,
         \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> ,
         \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> ,
         \op0_A<1> , \op0_A<0> , \op0_B<15> , \op0_B<14> , \op0_B<13> ,
         \op0_B<12> , \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> ,
         \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> ,
         \op0_B<2> , \op0_B<1> , \op0_B<0> , \op1_A<3> , \op1_A<2> ,
         \op1_A<1> , \op1_A<0> , \op1_B<15> , \op1_B<14> , \op1_B<13> ,
         \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> ,
         \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> ,
         \op1_B<2> , \op1_B<1> , \op1_B<0> , n59, n60, n62, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n61, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n116;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  OR2X2 U4 ( .A(n71), .B(n72), .Y(n62) );
  OAI21X1 U74 ( .A(n81), .B(n116), .C(n44), .Y(\Out<0> ) );
  NAND3X1 U76 ( .A(Cout), .B(n81), .C(n68), .Y(n59) );
  demux1to2_16_1 demux0 ( .In({\A_real<15> , \A_real<14> , \A_real<13> , 
        \A_real<12> , \A_real<11> , \A_real<10> , \A_real<9> , \A_real<8> , 
        \A_real<7> , \A_real<6> , \A_real<5> , \A_real<4> , \A_real<3> , 
        \A_real<2> , \A_real<1> , \A_real<0> }), .S(n81), .Out0({\op0_A<15> , 
        \op0_A<14> , \op0_A<13> , \op0_A<12> , \op0_A<11> , \op0_A<10> , 
        \op0_A<9> , \op0_A<8> , \op0_A<7> , \op0_A<6> , \op0_A<5> , \op0_A<4> , 
        \op0_A<3> , \op0_A<2> , \op0_A<1> , \op0_A<0> }), .Out1({\op0_B<15> , 
        \op0_B<14> , \op0_B<13> , \op0_B<12> , \op0_B<11> , \op0_B<10> , 
        \op0_B<9> , \op0_B<8> , \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , 
        \op0_B<3> , \op0_B<2> , \op0_B<1> , \op0_B<0> }) );
  demux1to2_16_0 demux1 ( .In({\B_real<15> , \B_real<14> , \B_real<13> , 
        \B_real<12> , \B_real<11> , \B_real<10> , \B_real<9> , \B_real<8> , 
        \B_real<7> , \B_real<6> , \B_real<5> , \B_real<4> , \B_real<3> , 
        \B_real<2> , \B_real<1> , \B_real<0> }), .S(n81), .Out0({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, \op1_A<3> , 
        \op1_A<2> , \op1_A<1> , \op1_A<0> }), .Out1({\op1_B<15> , \op1_B<14> , 
        \op1_B<13> , \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , 
        \op1_B<8> , \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , 
        \op1_B<2> , \op1_B<1> , \op1_B<0> }) );
  cla_or_xor_and coxa0 ( .A({\op0_B<15> , \op0_B<14> , \op0_B<13> , 
        \op0_B<12> , \op0_B<11> , \op0_B<10> , \op0_B<9> , \op0_B<8> , 
        \op0_B<7> , \op0_B<6> , \op0_B<5> , \op0_B<4> , \op0_B<3> , \op0_B<2> , 
        \op0_B<1> , \op0_B<0> }), .B({\op1_B<15> , \op1_B<14> , \op1_B<13> , 
        \op1_B<12> , \op1_B<11> , \op1_B<10> , \op1_B<9> , \op1_B<8> , 
        \op1_B<7> , \op1_B<6> , \op1_B<5> , \op1_B<4> , \op1_B<3> , \op1_B<2> , 
        \op1_B<1> , \op1_B<0> }), .Cin(Cin), .Op({\Op<1> , \Op<0> }), .Out({
        \op0_out<15> , \op0_out<14> , \op0_out<13> , \op0_out<12> , 
        \op0_out<11> , \op0_out<10> , \op0_out<9> , \op0_out<8> , \op0_out<7> , 
        \op0_out<6> , \op0_out<5> , \op0_out<4> , \op0_out<3> , \op0_out<2> , 
        \op0_out<1> , \op0_out<0> }), .Cout(Cout) );
  shifter shift ( .In({\op0_A<15> , \op0_A<14> , \op0_A<13> , \op0_A<12> , 
        \op0_A<11> , \op0_A<10> , \op0_A<9> , \op0_A<8> , \op0_A<7> , 
        \op0_A<6> , \op0_A<5> , \op0_A<4> , \op0_A<3> , \op0_A<2> , \op0_A<1> , 
        \op0_A<0> }), .Cnt({\op1_A<3> , \op1_A<2> , \op1_A<1> , \op1_A<0> }), 
        .Op({n71, n72}), .Out({\op1_out<15> , \op1_out<14> , \op1_out<13> , 
        \op1_out<12> , \op1_out<11> , \op1_out<10> , \op1_out<9> , 
        \op1_out<8> , \op1_out<7> , \op1_out<6> , \op1_out<5> , \op1_out<4> , 
        \op1_out<3> , \op1_out<2> , \op1_out<1> , \op1_out<0> }) );
  BUFX2 U1 ( .A(n74), .Y(n1) );
  BUFX2 U2 ( .A(\op0_out<5> ), .Y(n2) );
  AND2X2 U3 ( .A(n10), .B(n88), .Y(n3) );
  OR2X2 U5 ( .A(n81), .B(\op1_out<0> ), .Y(n4) );
  AND2X2 U6 ( .A(n22), .B(n64), .Y(n55) );
  AND2X1 U7 ( .A(n26), .B(n34), .Y(n65) );
  INVX1 U8 ( .A(n111), .Y(\A_real<15> ) );
  OR2X1 U9 ( .A(\op1_out<12> ), .B(\op1_out<13> ), .Y(n27) );
  OR2X1 U10 ( .A(\op1_out<8> ), .B(\op1_out<9> ), .Y(n29) );
  INVX1 U11 ( .A(n76), .Y(n9) );
  AND2X1 U12 ( .A(n50), .B(n46), .Y(n39) );
  INVX1 U13 ( .A(n80), .Y(n73) );
  INVX1 U14 ( .A(\op1_out<7> ), .Y(n96) );
  INVX1 U15 ( .A(\op0_out<3> ), .Y(n88) );
  INVX1 U16 ( .A(\op1_out<4> ), .Y(n91) );
  INVX1 U17 ( .A(\op1_out<6> ), .Y(n95) );
  INVX1 U18 ( .A(\op0_out<6> ), .Y(n94) );
  INVX1 U19 ( .A(\op1_out<8> ), .Y(n98) );
  INVX1 U20 ( .A(\op1_out<9> ), .Y(n100) );
  INVX1 U21 ( .A(\op1_out<10> ), .Y(n102) );
  INVX1 U22 ( .A(\op1_out<11> ), .Y(n104) );
  INVX1 U23 ( .A(\op1_out<12> ), .Y(n106) );
  INVX1 U24 ( .A(\op1_out<13> ), .Y(n108) );
  INVX1 U25 ( .A(\op1_out<14> ), .Y(n110) );
  INVX1 U26 ( .A(\op1_out<0> ), .Y(n116) );
  INVX1 U27 ( .A(\op0_out<7> ), .Y(n5) );
  MUX2X1 U28 ( .B(n107), .A(n108), .S(n82), .Y(\Out<13> ) );
  BUFX2 U29 ( .A(\op0_out<4> ), .Y(n6) );
  XNOR2X1 U30 ( .A(\A<9> ), .B(n78), .Y(\A_real<9> ) );
  XOR2X1 U31 ( .A(\B<1> ), .B(n76), .Y(\B_real<1> ) );
  INVX1 U32 ( .A(n77), .Y(n8) );
  XOR2X1 U33 ( .A(n7), .B(n8), .Y(\B_real<7> ) );
  INVX1 U34 ( .A(\B<7> ), .Y(n7) );
  INVX4 U35 ( .A(n75), .Y(n77) );
  MUX2X1 U36 ( .B(n105), .A(n106), .S(n82), .Y(\Out<12> ) );
  INVX1 U37 ( .A(\op0_out<13> ), .Y(n107) );
  MUX2X1 U38 ( .B(n5), .A(n96), .S(n82), .Y(\Out<7> ) );
  XNOR2X1 U39 ( .A(\B<2> ), .B(n9), .Y(\B_real<2> ) );
  INVX1 U40 ( .A(\op1_out<3> ), .Y(n89) );
  XOR2X1 U41 ( .A(\B<3> ), .B(n77), .Y(\B_real<3> ) );
  OR2X2 U42 ( .A(\op1_out<3> ), .B(\op1_out<2> ), .Y(n19) );
  AND2X2 U43 ( .A(n55), .B(n97), .Y(n10) );
  INVX1 U44 ( .A(\op0_out<2> ), .Y(n86) );
  INVX1 U45 ( .A(n2), .Y(n92) );
  XOR2X1 U46 ( .A(\B<0> ), .B(n76), .Y(\B_real<0> ) );
  INVX1 U47 ( .A(n6), .Y(n90) );
  OR2X2 U48 ( .A(\op0_out<1> ), .B(\op0_out<0> ), .Y(n11) );
  OR2X2 U49 ( .A(n67), .B(n13), .Y(n12) );
  OR2X2 U50 ( .A(n19), .B(n4), .Y(n13) );
  OR2X2 U51 ( .A(n20), .B(n16), .Y(n14) );
  OR2X2 U52 ( .A(\op0_out<9> ), .B(\op0_out<6> ), .Y(n15) );
  OR2X2 U53 ( .A(n61), .B(n15), .Y(n16) );
  AND2X2 U54 ( .A(n84), .B(n83), .Y(n17) );
  INVX1 U55 ( .A(n17), .Y(n18) );
  OR2X2 U56 ( .A(n74), .B(n63), .Y(n20) );
  OR2X2 U57 ( .A(\op0_out<4> ), .B(\op0_out<2> ), .Y(n21) );
  INVX1 U58 ( .A(n21), .Y(n22) );
  AND2X2 U59 ( .A(n52), .B(n48), .Y(n23) );
  INVX1 U60 ( .A(n23), .Y(\Out<1> ) );
  OR2X1 U61 ( .A(\op1_out<4> ), .B(\op1_out<5> ), .Y(n25) );
  INVX1 U62 ( .A(n25), .Y(n26) );
  INVX1 U63 ( .A(n27), .Y(n28) );
  INVX1 U64 ( .A(n29), .Y(n30) );
  OR2X2 U65 ( .A(\op0_out<5> ), .B(\op0_out<12> ), .Y(n31) );
  INVX1 U66 ( .A(n31), .Y(n32) );
  OR2X1 U67 ( .A(\op1_out<6> ), .B(\op1_out<7> ), .Y(n33) );
  INVX1 U68 ( .A(n33), .Y(n34) );
  OR2X2 U69 ( .A(\op1_out<14> ), .B(\op1_out<15> ), .Y(n35) );
  INVX1 U70 ( .A(n35), .Y(n36) );
  OR2X2 U71 ( .A(\op1_out<10> ), .B(\op1_out<11> ), .Y(n37) );
  INVX1 U72 ( .A(n37), .Y(n38) );
  INVX1 U73 ( .A(n39), .Y(n40) );
  AND2X2 U75 ( .A(\op1_out<15> ), .B(n82), .Y(n41) );
  INVX1 U77 ( .A(n41), .Y(n42) );
  AND2X2 U78 ( .A(\op0_out<0> ), .B(n81), .Y(n43) );
  INVX1 U79 ( .A(n43), .Y(n44) );
  OR2X2 U80 ( .A(n54), .B(n57), .Y(n45) );
  INVX1 U81 ( .A(n45), .Y(n46) );
  AND2X2 U82 ( .A(\op1_out<1> ), .B(n82), .Y(n47) );
  INVX1 U83 ( .A(n47), .Y(n48) );
  OR2X2 U84 ( .A(n66), .B(n12), .Y(n49) );
  INVX1 U85 ( .A(n49), .Y(n50) );
  AND2X2 U86 ( .A(\op0_out<1> ), .B(n81), .Y(n51) );
  INVX1 U87 ( .A(n51), .Y(n52) );
  AND2X2 U88 ( .A(n28), .B(n36), .Y(n53) );
  INVX1 U89 ( .A(n53), .Y(n54) );
  AND2X2 U90 ( .A(n30), .B(n38), .Y(n56) );
  INVX1 U91 ( .A(n56), .Y(n57) );
  AND2X2 U92 ( .A(n32), .B(n3), .Y(n58) );
  INVX1 U93 ( .A(n58), .Y(n61) );
  BUFX2 U94 ( .A(\op0_out<15> ), .Y(n63) );
  INVX1 U95 ( .A(n11), .Y(n64) );
  INVX1 U96 ( .A(n65), .Y(n66) );
  INVX1 U97 ( .A(n85), .Y(n67) );
  INVX1 U98 ( .A(\op1_out<1> ), .Y(n85) );
  INVX1 U99 ( .A(n59), .Y(Ofl) );
  BUFX2 U100 ( .A(n60), .Y(n68) );
  INVX1 U101 ( .A(\op0_out<11> ), .Y(n103) );
  OAI21X1 U102 ( .A(n69), .B(n82), .C(n42), .Y(\Out<15> ) );
  INVX1 U103 ( .A(n63), .Y(n69) );
  OAI21X1 U104 ( .A(n14), .B(n18), .C(n40), .Y(Z) );
  INVX1 U105 ( .A(\op1_out<5> ), .Y(n93) );
  XNOR2X1 U106 ( .A(\A<1> ), .B(n78), .Y(\A_real<1> ) );
  INVX2 U107 ( .A(n78), .Y(n80) );
  INVX1 U108 ( .A(\op1_out<2> ), .Y(n87) );
  XNOR2X1 U109 ( .A(\A<4> ), .B(n70), .Y(\A_real<4> ) );
  INVX8 U110 ( .A(n79), .Y(n70) );
  XOR2X1 U111 ( .A(\A<5> ), .B(n80), .Y(\A_real<5> ) );
  XOR2X1 U112 ( .A(\B<11> ), .B(invB), .Y(\B_real<11> ) );
  BUFX2 U113 ( .A(\Op<1> ), .Y(n71) );
  BUFX2 U114 ( .A(\Op<0> ), .Y(n72) );
  XNOR2X1 U115 ( .A(\A<7> ), .B(n78), .Y(\A_real<7> ) );
  XNOR2X1 U116 ( .A(\A<10> ), .B(n78), .Y(\A_real<10> ) );
  XNOR2X1 U117 ( .A(\A<0> ), .B(n70), .Y(\A_real<0> ) );
  XNOR2X1 U118 ( .A(\A<11> ), .B(n73), .Y(\A_real<11> ) );
  INVX1 U119 ( .A(\op0_out<9> ), .Y(n99) );
  XNOR2X1 U120 ( .A(\A<3> ), .B(n78), .Y(\A_real<3> ) );
  XNOR2X1 U121 ( .A(\A<2> ), .B(n70), .Y(\A_real<2> ) );
  INVX1 U122 ( .A(\op0_out<10> ), .Y(n101) );
  XNOR2X1 U123 ( .A(\A<8> ), .B(n70), .Y(\A_real<8> ) );
  BUFX2 U124 ( .A(\op0_out<14> ), .Y(n74) );
  INVX1 U125 ( .A(\op0_out<12> ), .Y(n105) );
  INVX1 U126 ( .A(n1), .Y(n109) );
  INVX1 U127 ( .A(\op0_out<8> ), .Y(n97) );
  INVX8 U128 ( .A(invB), .Y(n75) );
  INVX8 U129 ( .A(n75), .Y(n76) );
  INVX8 U130 ( .A(invA), .Y(n78) );
  INVX8 U131 ( .A(n78), .Y(n79) );
  INVX8 U132 ( .A(n82), .Y(n81) );
  INVX8 U133 ( .A(\Op<2> ), .Y(n82) );
  XNOR2X1 U134 ( .A(\B<15> ), .B(n77), .Y(n112) );
  INVX2 U135 ( .A(n112), .Y(\B_real<15> ) );
  XOR2X1 U136 ( .A(\B<14> ), .B(n76), .Y(\B_real<14> ) );
  XOR2X1 U137 ( .A(\B<13> ), .B(n77), .Y(\B_real<13> ) );
  XOR2X1 U138 ( .A(\B<12> ), .B(n76), .Y(\B_real<12> ) );
  XOR2X1 U139 ( .A(\B<10> ), .B(n76), .Y(\B_real<10> ) );
  XOR2X1 U140 ( .A(\B<9> ), .B(n77), .Y(\B_real<9> ) );
  XOR2X1 U141 ( .A(\B<8> ), .B(n76), .Y(\B_real<8> ) );
  XOR2X1 U142 ( .A(\B<6> ), .B(n76), .Y(\B_real<6> ) );
  XOR2X1 U143 ( .A(\B<5> ), .B(n77), .Y(\B_real<5> ) );
  XOR2X1 U144 ( .A(\B<4> ), .B(n76), .Y(\B_real<4> ) );
  XNOR2X1 U145 ( .A(\A<15> ), .B(n80), .Y(n111) );
  XOR2X1 U146 ( .A(\A<14> ), .B(n79), .Y(\A_real<14> ) );
  XOR2X1 U147 ( .A(\A<13> ), .B(n80), .Y(\A_real<13> ) );
  XOR2X1 U148 ( .A(\A<12> ), .B(n79), .Y(\A_real<12> ) );
  XOR2X1 U149 ( .A(\A<6> ), .B(n79), .Y(\A_real<6> ) );
  NOR2X1 U150 ( .A(\op0_out<11> ), .B(n82), .Y(n84) );
  NOR3X1 U151 ( .A(\op0_out<13> ), .B(\op0_out<10> ), .C(\op0_out<7> ), .Y(n83) );
  MUX2X1 U152 ( .B(n87), .A(n86), .S(n81), .Y(\Out<2> ) );
  MUX2X1 U153 ( .B(n89), .A(n88), .S(n81), .Y(\Out<3> ) );
  MUX2X1 U154 ( .B(n91), .A(n90), .S(n81), .Y(\Out<4> ) );
  MUX2X1 U155 ( .B(n93), .A(n92), .S(n81), .Y(\Out<5> ) );
  MUX2X1 U156 ( .B(n95), .A(n94), .S(n81), .Y(\Out<6> ) );
  MUX2X1 U157 ( .B(n98), .A(n97), .S(n81), .Y(\Out<8> ) );
  MUX2X1 U158 ( .B(n100), .A(n99), .S(n81), .Y(\Out<9> ) );
  MUX2X1 U159 ( .B(n102), .A(n101), .S(n81), .Y(\Out<10> ) );
  MUX2X1 U160 ( .B(n104), .A(n103), .S(n81), .Y(\Out<11> ) );
  MUX2X1 U161 ( .B(n110), .A(n109), .S(n81), .Y(\Out<14> ) );
  XNOR2X1 U162 ( .A(n112), .B(n111), .Y(n113) );
  AOI21X1 U163 ( .A(sign), .B(n113), .C(n62), .Y(n60) );
endmodule


module mux4to1_16_5 ( .InA({\InA<15> , \InA<14> , \InA<13> , \InA<12> , 
        \InA<11> , \InA<10> , \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , 
        \InA<4> , \InA<3> , \InA<2> , \InA<1> , \InA<0> }), .InB({\InB<15> , 
        \InB<14> , \InB<13> , \InB<12> , \InB<11> , \InB<10> , \InB<9> , 
        \InB<8> , \InB<7> , \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , 
        \InB<1> , \InB<0> }), .InC({\InC<15> , \InC<14> , \InC<13> , \InC<12> , 
        \InC<11> , \InC<10> , \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , 
        \InC<4> , \InC<3> , \InC<2> , \InC<1> , \InC<0> }), .InD({\InD<15> , 
        \InD<14> , \InD<13> , \InD<12> , \InD<11> , \InD<10> , \InD<9> , 
        \InD<8> , \InD<7> , \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , 
        \InD<1> , \InD<0> }), .S({\S<1> , \S<0> }), .Out({\Out<15> , \Out<14> , 
        \Out<13> , \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , 
        \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , 
        \Out<0> }) );
  input \InA<15> , \InA<14> , \InA<13> , \InA<12> , \InA<11> , \InA<10> ,
         \InA<9> , \InA<8> , \InA<7> , \InA<6> , \InA<5> , \InA<4> , \InA<3> ,
         \InA<2> , \InA<1> , \InA<0> , \InB<15> , \InB<14> , \InB<13> ,
         \InB<12> , \InB<11> , \InB<10> , \InB<9> , \InB<8> , \InB<7> ,
         \InB<6> , \InB<5> , \InB<4> , \InB<3> , \InB<2> , \InB<1> , \InB<0> ,
         \InC<15> , \InC<14> , \InC<13> , \InC<12> , \InC<11> , \InC<10> ,
         \InC<9> , \InC<8> , \InC<7> , \InC<6> , \InC<5> , \InC<4> , \InC<3> ,
         \InC<2> , \InC<1> , \InC<0> , \InD<15> , \InD<14> , \InD<13> ,
         \InD<12> , \InD<11> , \InD<10> , \InD<9> , \InD<8> , \InD<7> ,
         \InD<6> , \InD<5> , \InD<4> , \InD<3> , \InD<2> , \InD<1> , \InD<0> ,
         \S<1> , \S<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n3, n4, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n1, n2, n5, n6, n7, n8, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71, n73,
         n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, n100,
         n101, n102, n103, n104;

  AOI22X1 U5 ( .A(\InA<9> ), .B(n104), .C(\InB<9> ), .D(n5), .Y(n4) );
  AOI22X1 U6 ( .A(\InC<9> ), .B(n7), .C(\InD<9> ), .D(n6), .Y(n3) );
  AOI22X1 U8 ( .A(\InA<8> ), .B(n104), .C(\InB<8> ), .D(n5), .Y(n10) );
  AOI22X1 U9 ( .A(\InC<8> ), .B(n7), .C(\InD<8> ), .D(n6), .Y(n9) );
  AOI22X1 U11 ( .A(\InA<7> ), .B(n104), .C(\InB<7> ), .D(n5), .Y(n12) );
  AOI22X1 U12 ( .A(\InC<7> ), .B(n7), .C(\InD<7> ), .D(n6), .Y(n11) );
  AOI22X1 U14 ( .A(\InA<6> ), .B(n104), .C(\InB<6> ), .D(n5), .Y(n14) );
  AOI22X1 U15 ( .A(\InC<6> ), .B(n7), .C(\InD<6> ), .D(n6), .Y(n13) );
  AOI22X1 U17 ( .A(\InA<5> ), .B(n104), .C(\InB<5> ), .D(n5), .Y(n16) );
  AOI22X1 U18 ( .A(\InC<5> ), .B(n7), .C(\InD<5> ), .D(n6), .Y(n15) );
  AOI22X1 U20 ( .A(\InA<4> ), .B(n104), .C(\InB<4> ), .D(n5), .Y(n18) );
  AOI22X1 U21 ( .A(\InC<4> ), .B(n7), .C(\InD<4> ), .D(n6), .Y(n17) );
  AOI22X1 U23 ( .A(\InA<3> ), .B(n104), .C(\InB<3> ), .D(n5), .Y(n20) );
  AOI22X1 U24 ( .A(\InC<3> ), .B(n7), .C(\InD<3> ), .D(n6), .Y(n19) );
  AOI22X1 U26 ( .A(\InA<2> ), .B(n104), .C(\InB<2> ), .D(n5), .Y(n22) );
  AOI22X1 U27 ( .A(\InC<2> ), .B(n7), .C(\InD<2> ), .D(n6), .Y(n21) );
  AOI22X1 U29 ( .A(\InA<1> ), .B(n104), .C(\InB<1> ), .D(n5), .Y(n24) );
  AOI22X1 U30 ( .A(\InC<1> ), .B(n7), .C(\InD<1> ), .D(n6), .Y(n23) );
  AOI22X1 U32 ( .A(\InA<15> ), .B(n104), .C(\InB<15> ), .D(n5), .Y(n26) );
  AOI22X1 U33 ( .A(\InC<15> ), .B(n7), .C(\InD<15> ), .D(n6), .Y(n25) );
  AOI22X1 U35 ( .A(\InA<14> ), .B(n104), .C(\InB<14> ), .D(n5), .Y(n28) );
  AOI22X1 U36 ( .A(\InC<14> ), .B(n7), .C(\InD<14> ), .D(n6), .Y(n27) );
  AOI22X1 U38 ( .A(\InA<13> ), .B(n104), .C(\InB<13> ), .D(n5), .Y(n30) );
  AOI22X1 U39 ( .A(\InC<13> ), .B(n7), .C(\InD<13> ), .D(n6), .Y(n29) );
  AOI22X1 U41 ( .A(\InA<12> ), .B(n104), .C(\InB<12> ), .D(n5), .Y(n32) );
  AOI22X1 U42 ( .A(\InC<12> ), .B(n7), .C(\InD<12> ), .D(n6), .Y(n31) );
  AOI22X1 U44 ( .A(\InA<11> ), .B(n104), .C(\InB<11> ), .D(n5), .Y(n34) );
  AOI22X1 U45 ( .A(\InC<11> ), .B(n7), .C(\InD<11> ), .D(n6), .Y(n33) );
  AOI22X1 U47 ( .A(\InA<10> ), .B(n104), .C(\InB<10> ), .D(n5), .Y(n36) );
  AOI22X1 U48 ( .A(\InC<10> ), .B(n7), .C(\InD<10> ), .D(n6), .Y(n35) );
  INVX1 U1 ( .A(\S<0> ), .Y(n101) );
  OR2X1 U2 ( .A(\S<1> ), .B(\S<0> ), .Y(n100) );
  INVX1 U3 ( .A(\S<1> ), .Y(n99) );
  AND2X1 U4 ( .A(n43), .B(n58), .Y(n69) );
  AND2X1 U7 ( .A(n44), .B(n59), .Y(n83) );
  AND2X1 U10 ( .A(n45), .B(n60), .Y(n85) );
  AND2X1 U13 ( .A(n46), .B(n61), .Y(n87) );
  AND2X1 U16 ( .A(n47), .B(n62), .Y(n89) );
  AND2X1 U19 ( .A(n48), .B(n63), .Y(n91) );
  AND2X1 U22 ( .A(n49), .B(n64), .Y(n93) );
  AND2X1 U25 ( .A(n50), .B(n65), .Y(n95) );
  AND2X1 U28 ( .A(n51), .B(n66), .Y(n97) );
  AND2X1 U31 ( .A(n37), .B(n52), .Y(n71) );
  AND2X1 U34 ( .A(n38), .B(n53), .Y(n73) );
  AND2X1 U37 ( .A(n39), .B(n54), .Y(n75) );
  AND2X1 U40 ( .A(n40), .B(n55), .Y(n77) );
  AND2X1 U43 ( .A(n41), .B(n56), .Y(n79) );
  AND2X1 U46 ( .A(n42), .B(n57), .Y(n81) );
  BUFX2 U49 ( .A(n102), .Y(n1) );
  BUFX2 U50 ( .A(n103), .Y(n2) );
  AND2X1 U51 ( .A(\S<0> ), .B(n99), .Y(n5) );
  AND2X1 U52 ( .A(\S<0> ), .B(\S<1> ), .Y(n6) );
  AND2X1 U53 ( .A(n101), .B(\S<1> ), .Y(n7) );
  AND2X1 U54 ( .A(\InD<0> ), .B(n6), .Y(n8) );
  BUFX2 U55 ( .A(n35), .Y(n37) );
  BUFX2 U56 ( .A(n33), .Y(n38) );
  BUFX2 U57 ( .A(n31), .Y(n39) );
  BUFX2 U58 ( .A(n29), .Y(n40) );
  BUFX2 U59 ( .A(n27), .Y(n41) );
  BUFX2 U60 ( .A(n25), .Y(n42) );
  BUFX2 U61 ( .A(n23), .Y(n43) );
  BUFX2 U62 ( .A(n21), .Y(n44) );
  BUFX2 U63 ( .A(n19), .Y(n45) );
  BUFX2 U64 ( .A(n17), .Y(n46) );
  BUFX2 U65 ( .A(n15), .Y(n47) );
  BUFX2 U66 ( .A(n13), .Y(n48) );
  BUFX2 U67 ( .A(n11), .Y(n49) );
  BUFX2 U68 ( .A(n9), .Y(n50) );
  BUFX2 U69 ( .A(n3), .Y(n51) );
  BUFX2 U70 ( .A(n36), .Y(n52) );
  BUFX2 U71 ( .A(n34), .Y(n53) );
  BUFX2 U72 ( .A(n32), .Y(n54) );
  BUFX2 U73 ( .A(n30), .Y(n55) );
  BUFX2 U74 ( .A(n28), .Y(n56) );
  BUFX2 U75 ( .A(n26), .Y(n57) );
  BUFX2 U76 ( .A(n24), .Y(n58) );
  BUFX2 U77 ( .A(n22), .Y(n59) );
  BUFX2 U78 ( .A(n20), .Y(n60) );
  BUFX2 U79 ( .A(n18), .Y(n61) );
  BUFX2 U80 ( .A(n16), .Y(n62) );
  BUFX2 U81 ( .A(n14), .Y(n63) );
  BUFX2 U82 ( .A(n12), .Y(n64) );
  BUFX2 U83 ( .A(n10), .Y(n65) );
  BUFX2 U84 ( .A(n4), .Y(n66) );
  OR2X1 U85 ( .A(n5), .B(n8), .Y(n67) );
  INVX1 U86 ( .A(n67), .Y(n68) );
  INVX1 U87 ( .A(n69), .Y(\Out<1> ) );
  INVX1 U88 ( .A(n71), .Y(\Out<10> ) );
  INVX1 U89 ( .A(n73), .Y(\Out<11> ) );
  INVX1 U90 ( .A(n75), .Y(\Out<12> ) );
  INVX1 U91 ( .A(n77), .Y(\Out<13> ) );
  INVX1 U92 ( .A(n79), .Y(\Out<14> ) );
  INVX1 U93 ( .A(n81), .Y(\Out<15> ) );
  INVX1 U94 ( .A(n83), .Y(\Out<2> ) );
  INVX1 U95 ( .A(n85), .Y(\Out<3> ) );
  INVX1 U96 ( .A(n87), .Y(\Out<4> ) );
  INVX1 U97 ( .A(n89), .Y(\Out<5> ) );
  INVX1 U98 ( .A(n91), .Y(\Out<6> ) );
  INVX1 U99 ( .A(n93), .Y(\Out<7> ) );
  INVX1 U100 ( .A(n95), .Y(\Out<8> ) );
  INVX1 U101 ( .A(n97), .Y(\Out<9> ) );
  AOI21X1 U102 ( .A(n6), .B(\InD<0> ), .C(\InB<0> ), .Y(n103) );
  AOI22X1 U103 ( .A(n104), .B(\InA<0> ), .C(n7), .D(\InC<0> ), .Y(n102) );
  INVX1 U104 ( .A(n100), .Y(n104) );
  OAI21X1 U105 ( .A(n68), .B(n2), .C(n1), .Y(\Out<0> ) );
endmodule


module cla16_1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), Cout );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   \G<3> , \G<2> , \G<1> , \G<0> , \P<3> , \P<2> , \P<1> , \P<0> , n1,
         n2, n3, n9, n10, n11, n12, n13, n14, n15;

  AOI21X1 U5 ( .A(\P<3> ), .B(n9), .C(\G<3> ), .Y(n15) );
  AOI21X1 U6 ( .A(\P<2> ), .B(n10), .C(\G<2> ), .Y(n14) );
  AOI21X1 U7 ( .A(\P<1> ), .B(n11), .C(\G<1> ), .Y(n13) );
  AOI21X1 U8 ( .A(\P<0> ), .B(Cin), .C(\G<0> ), .Y(n12) );
  cla4_7 ca0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        .Cout(), .PG(\P<0> ), .GG(\G<0> ) );
  cla4_6 ca1 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(n2), .S({\S<7> , \S<6> , \S<5> , \S<4> }), 
        .Cout(), .PG(\P<1> ), .GG(\G<1> ) );
  cla4_5 ca2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(n10), .S({\S<11> , \S<10> , \S<9> , \S<8> }), 
        .Cout(), .PG(\P<2> ), .GG(\G<2> ) );
  cla4_4 ca3 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> }), .Cin(n9), .S({\S<15> , \S<14> , \S<13> , \S<12> }), 
        .Cout(), .PG(\P<3> ), .GG(\G<3> ) );
  BUFX2 U1 ( .A(n14), .Y(n1) );
  BUFX2 U2 ( .A(n11), .Y(n2) );
  INVX1 U3 ( .A(n12), .Y(n11) );
  INVX1 U4 ( .A(n13), .Y(n10) );
  BUFX2 U9 ( .A(n15), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(Cout) );
  INVX2 U11 ( .A(n1), .Y(n9) );
endmodule


module mux4to1 ( InA, InB, InC, InD, .S({\S<1> , \S<0> }), Out );
  input InA, InB, InC, InD, \S<1> , \S<0> ;
  output Out;
  wire   n4, n5, n6, n1, n2;

  OAI21X1 U3 ( .A(\S<1> ), .B(n4), .C(n5), .Y(Out) );
  NAND2X1 U4 ( .A(n1), .B(\S<1> ), .Y(n5) );
  AOI22X1 U5 ( .A(InC), .B(n2), .C(InD), .D(\S<0> ), .Y(n6) );
  AOI22X1 U6 ( .A(InA), .B(n2), .C(\S<0> ), .D(InB), .Y(n4) );
  INVX1 U1 ( .A(\S<0> ), .Y(n2) );
  INVX1 U2 ( .A(n6), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memory2c_0 ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, \mem<0><7> , \mem<0><6> , \mem<0><5> ,
         \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> ,
         \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> ,
         \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> ,
         \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> ,
         \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> ,
         \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> ,
         \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> ,
         \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> ,
         \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> ,
         \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> ,
         \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> ,
         \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> ,
         \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> ,
         \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> ,
         \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> ,
         \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> ,
         \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> ,
         \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> ,
         \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> ,
         \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> ,
         \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> ,
         \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> ,
         \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> ,
         \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> ,
         \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> ,
         \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> ,
         \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> ,
         \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> ,
         \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> ,
         \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> ,
         \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> ,
         \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> ,
         \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> ,
         \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> ,
         \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> ,
         \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> ,
         \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> ,
         \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> ,
         \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> , \mem<33><4> ,
         \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> , \mem<34><7> ,
         \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> , \mem<34><2> ,
         \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> , \mem<35><5> ,
         \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> , \mem<35><0> ,
         \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> , \mem<36><3> ,
         \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> , \mem<37><6> ,
         \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> , \mem<37><1> ,
         \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> , \mem<38><4> ,
         \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> , \mem<39><7> ,
         \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> , \mem<39><2> ,
         \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> , \mem<40><5> ,
         \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> , \mem<40><0> ,
         \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> , \mem<41><3> ,
         \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> , \mem<42><6> ,
         \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> , \mem<42><1> ,
         \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> , \mem<43><4> ,
         \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> , \mem<44><7> ,
         \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> , \mem<44><2> ,
         \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> , \mem<45><5> ,
         \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> , \mem<45><0> ,
         \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> , \mem<46><3> ,
         \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> , \mem<47><6> ,
         \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> , \mem<47><1> ,
         \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> , \mem<48><4> ,
         \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> , \mem<49><7> ,
         \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> , \mem<49><2> ,
         \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> , \mem<50><5> ,
         \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> , \mem<50><0> ,
         \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> , \mem<51><3> ,
         \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> , \mem<52><6> ,
         \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> , \mem<52><1> ,
         \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> , \mem<53><4> ,
         \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> , \mem<54><7> ,
         \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> , \mem<54><2> ,
         \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> , \mem<55><5> ,
         \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> , \mem<55><0> ,
         \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> , \mem<56><3> ,
         \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> , \mem<57><6> ,
         \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> , \mem<57><1> ,
         \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> , \mem<58><4> ,
         \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> , \mem<59><7> ,
         \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> , \mem<59><2> ,
         \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> , \mem<60><5> ,
         \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> , \mem<60><0> ,
         \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> , \mem<61><3> ,
         \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> , \mem<62><6> ,
         \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> , \mem<62><1> ,
         \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> , \mem<63><4> ,
         \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> , N185, N186,
         N187, N188, N189, N190, N191, N192, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n609, n611, n624, n637, n649, n661, n673, n685, n697, n709, n721,
         n733, n745, n757, n769, n781, n793, n805, n817, n829, n841, n853,
         n865, n877, n889, n901, n913, n925, n937, n949, n961, n973, n985,
         n997, n1009, n1021, n1033, n1045, n1057, n1069, n1081, n1093, n1105,
         n1117, n1129, n1141, n1153, n1165, n1177, n1189, n1201, n1213, n1225,
         n1237, n1249, n1261, n1273, n1285, n1297, n1309, n1321, n1333, n1345,
         n1357, n1358, n1371, n1372, n1383, n1384, n1396, n1397, n1409, n1410,
         n1424, n1425, n1436, n1437, n1449, n1450, n1461, n1462, n1476, n1477,
         n1488, n1489, n1501, n1502, n1513, n1514, n1528, n1529, n1540, n1541,
         n1553, n1554, n1565, n1566, n1580, n1581, n1592, n1593, n1605, n1606,
         n1617, n1618, n1632, n1633, n1644, n1645, n1657, n1658, n1669, n1670,
         n1684, n1685, n1696, n1697, n1709, n1710, n1721, n1722, n1736, n1737,
         n1758, n1759, n1771, n1773, n1775, n1776, n1783, n1793, n1795, n1796,
         n1802, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n3206), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n3207), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n3208), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n3209), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n3210), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n3211), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n3212), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n3213), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n3214), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n3215), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n3216), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n3217), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n3218), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n3219), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n3220), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n3221), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n3222), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n3223), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n3224), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n3225), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n3226), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n3227), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n3228), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n3229), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n3230), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n3231), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n3232), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n3233), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n3234), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n3235), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n3236), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n3237), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n3238), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n3239), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n3240), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n3241), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n3242), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n3243), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n3244), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n3245), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n3246), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n3247), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n3248), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n3249), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n3250), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n3251), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n3252), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n3253), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n3254), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n3255), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n3256), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n3257), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n3258), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n3259), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n3260), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n3261), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n3262), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n3263), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n3264), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n3265), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n3266), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n3267), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n3268), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n3269), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n3270), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n3271), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n3272), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n3273), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n3274), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n3275), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n3276), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n3277), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n3278), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n3279), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n3280), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n3281), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n3282), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n3283), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n3284), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n3285), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n3286), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n3287), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n3288), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n3289), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n3290), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n3291), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n3292), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n3293), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n3294), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n3295), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n3296), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n3297), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n3298), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n3299), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n3300), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n3301), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n3302), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n3303), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n3304), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n3305), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n3306), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n3307), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n3308), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n3309), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n3310), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n3311), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n3312), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n3313), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n3314), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n3315), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n3316), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n3317), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n3318), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n3319), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n3320), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n3321), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n3322), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n3323), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n3324), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n3325), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n3326), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n3327), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n3328), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n3329), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n3330), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n3331), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n3332), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n3333), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n3334), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n3335), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n3336), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n3337), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n3338), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n3339), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n3340), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n3341), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n3342), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n3343), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n3344), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n3345), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n3346), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n3347), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n3348), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n3349), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n3350), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n3351), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n3352), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n3353), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n3354), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n3355), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n3356), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n3357), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n3358), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n3359), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n3360), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n3361), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n3362), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n3363), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n3364), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n3365), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n3366), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n3367), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n3368), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n3369), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n3370), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n3371), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n3372), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n3373), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n3374), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n3375), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n3376), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n3377), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n3378), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n3379), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n3380), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n3381), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n3382), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n3383), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n3384), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n3385), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n3386), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n3387), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n3388), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n3389), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n3390), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n3391), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n3392), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n3393), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n3394), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n3395), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n3396), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n3397), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n3398), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n3399), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n3400), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n3401), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n3402), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n3403), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n3404), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n3405), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n3406), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n3407), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n3408), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n3409), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n3410), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n3411), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n3412), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n3413), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n3414), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n3415), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n3416), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n3417), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n3418), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n3419), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n3420), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n3421), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n3422), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n3423), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n3424), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n3425), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n3426), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n3427), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n3428), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n3429), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n3430), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n3431), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n3432), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n3433), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n3434), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n3435), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n3436), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n3437), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n3438), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n3439), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n3440), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n3441), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n3442), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n3443), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n3444), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n3445), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n3446), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n3447), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n3448), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n3449), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n3450), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n3451), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n3452), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n3453), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n3454), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n3455), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n3456), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n3457), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n3458), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n3459), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n3460), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n3461), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n3462), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n3463), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n3464), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n3465), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n3466), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n3467), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n3468), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n3469), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n3470), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n3471), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n3472), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n3473), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n3474), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n3475), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n3476), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n3477), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n3478), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n3479), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n3480), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n3481), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n3482), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n3483), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n3484), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n3485), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n3486), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n3487), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n3488), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n3489), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n3490), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n3491), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n3492), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n3493), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n3494), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n3495), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n3496), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n3497), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n3498), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n3499), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n3500), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n3501), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n3502), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n3503), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n3504), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n3505), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n3506), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n3507), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n3508), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n3509), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n3510), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n3511), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n3512), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n3513), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n3514), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n3515), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n3516), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n3517), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n3518), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n3519), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n3520), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n3521), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n3522), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n3523), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n3524), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n3525), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n3526), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n3527), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n3528), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n3529), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n3530), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n3531), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n3532), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n3533), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n3534), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n3535), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n3536), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n3537), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n3538), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n3539), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n3540), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n3541), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n3542), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n3543), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n3544), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n3545), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n3546), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n3547), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n3548), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n3549), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n3550), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n3551), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n3552), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n3553), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n3554), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n3555), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n3556), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n3557), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n3558), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n3559), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n3560), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n3561), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n3562), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n3563), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n3564), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n3565), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n3566), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n3567), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n3568), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n3569), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n3570), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n3571), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n3572), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n3573), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n3574), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n3575), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n3576), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n3577), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n3578), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n3579), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n3580), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n3581), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n3582), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n3583), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n3584), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n3585), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n3586), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n3587), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n3588), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n3589), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n3590), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n3591), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n3592), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n3593), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n3594), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n3595), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n3596), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n3597), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n3598), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n3599), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n3600), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n3601), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n3602), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n3603), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n3604), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n3605), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n3606), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n3607), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n3608), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n3609), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n3610), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n3611), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n3612), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n3613), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n3614), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n3615), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n3616), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n3617), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n3618), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n3619), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n3620), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n3621), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n3622), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n3623), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n3624), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n3625), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n3626), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n3627), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n3628), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n3629), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n3630), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n3631), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n3632), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n3633), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n3634), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n3635), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n3636), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n3637), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n3638), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n3639), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n3640), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n3641), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n3642), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n3643), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n3644), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n3645), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n3646), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n3647), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n3648), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n3649), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n3650), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n3651), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n3652), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n3653), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n3654), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n3655), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n3656), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n3657), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n3658), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n3659), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n3660), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n3661), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n3662), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n3663), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n3664), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n3665), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n3666), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n3667), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n3668), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n3669), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n3670), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n3671), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n3672), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n3673), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n3674), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n3675), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n3676), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n3677), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n3678), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n3679), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n3680), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n3681), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n3682), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n3683), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n3684), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n3685), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n3686), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n3687), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n3688), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n3689), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n3690), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n3691), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n3692), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n3693), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n3694), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n3695), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n3696), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n3697), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n3698), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n3699), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n3700), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n3701), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n3702), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n3703), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n3704), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n3705), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n3706), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n3707), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n3708), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n3709), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n3710), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n3711), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n3712), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n3713), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n3714), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n3715), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n3716), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n3717), .CLK(clk), .Q(\mem<63><0> ) );
  AND2X2 U132 ( .A(n4090), .B(n4089), .Y(n4091) );
  AND2X2 U133 ( .A(n4085), .B(n4084), .Y(n4086) );
  AND2X2 U135 ( .A(n4080), .B(n4079), .Y(n4081) );
  AND2X2 U136 ( .A(n4075), .B(n4074), .Y(n4076) );
  AND2X2 U137 ( .A(n4069), .B(n4068), .Y(n4070) );
  AND2X2 U138 ( .A(n4063), .B(n4062), .Y(n4064) );
  AND2X2 U140 ( .A(n4058), .B(n4057), .Y(n4059) );
  AND2X2 U141 ( .A(n4053), .B(n4052), .Y(n4054) );
  AND2X2 U142 ( .A(n4045), .B(n4044), .Y(n4046) );
  AND2X2 U143 ( .A(n4040), .B(n4039), .Y(n4041) );
  AND2X2 U145 ( .A(n4035), .B(n4034), .Y(n4036) );
  AND2X2 U146 ( .A(n4030), .B(n4029), .Y(n4031) );
  AND2X2 U147 ( .A(n4024), .B(n4023), .Y(n4025) );
  AND2X2 U148 ( .A(n4019), .B(n4018), .Y(n4020) );
  AND2X2 U150 ( .A(n4014), .B(n4013), .Y(n4015) );
  AND2X2 U151 ( .A(n4009), .B(n4008), .Y(n4010) );
  AND2X2 U152 ( .A(n4001), .B(n4000), .Y(n4002) );
  AND2X2 U153 ( .A(n3996), .B(n3995), .Y(n3997) );
  AND2X2 U155 ( .A(n3991), .B(n3990), .Y(n3992) );
  AND2X2 U156 ( .A(n3986), .B(n3985), .Y(n3987) );
  AND2X2 U157 ( .A(n3980), .B(n3979), .Y(n3981) );
  AND2X2 U158 ( .A(n3975), .B(n3974), .Y(n3976) );
  AND2X2 U160 ( .A(n3970), .B(n3969), .Y(n3971) );
  AND2X2 U161 ( .A(n3965), .B(n3964), .Y(n3966) );
  AND2X2 U162 ( .A(n3957), .B(n3956), .Y(n3958) );
  AND2X2 U163 ( .A(n3952), .B(n3951), .Y(n3953) );
  AND2X2 U165 ( .A(n3947), .B(n3946), .Y(n3948) );
  AND2X2 U166 ( .A(n3942), .B(n3941), .Y(n3943) );
  AND2X2 U167 ( .A(n3936), .B(n3935), .Y(n3937) );
  AND2X2 U168 ( .A(n3931), .B(n3930), .Y(n3932) );
  AND2X2 U170 ( .A(n3926), .B(n3925), .Y(n3927) );
  AND2X2 U171 ( .A(n3921), .B(n3920), .Y(n3922) );
  AND2X2 U172 ( .A(n3913), .B(n3912), .Y(n3914) );
  AND2X2 U173 ( .A(n3908), .B(n3907), .Y(n3909) );
  AND2X2 U175 ( .A(n3903), .B(n3902), .Y(n3904) );
  AND2X2 U176 ( .A(n3898), .B(n3897), .Y(n3899) );
  AND2X2 U177 ( .A(n3892), .B(n3891), .Y(n3893) );
  AND2X2 U178 ( .A(n3887), .B(n3886), .Y(n3888) );
  AND2X2 U180 ( .A(n3882), .B(n3881), .Y(n3883) );
  AND2X2 U181 ( .A(n3877), .B(n3876), .Y(n3878) );
  AND2X2 U182 ( .A(n3869), .B(n3868), .Y(n3870) );
  AND2X2 U183 ( .A(n3864), .B(n3863), .Y(n3865) );
  AND2X2 U185 ( .A(n3859), .B(n3858), .Y(n3860) );
  AND2X2 U186 ( .A(n3854), .B(n3853), .Y(n3855) );
  AND2X2 U187 ( .A(n3848), .B(n3847), .Y(n3849) );
  AND2X2 U188 ( .A(n3843), .B(n3842), .Y(n3844) );
  AND2X2 U190 ( .A(n3838), .B(n3837), .Y(n3839) );
  AND2X2 U191 ( .A(n3833), .B(n3832), .Y(n3834) );
  AND2X2 U192 ( .A(n3825), .B(n3824), .Y(n3826) );
  AND2X2 U193 ( .A(n3820), .B(n3819), .Y(n3821) );
  AND2X2 U195 ( .A(n3815), .B(n3814), .Y(n3816) );
  AND2X2 U196 ( .A(n3810), .B(n3809), .Y(n3811) );
  AND2X2 U197 ( .A(n3804), .B(n3803), .Y(n3805) );
  AND2X2 U198 ( .A(n3799), .B(n3798), .Y(n3800) );
  AND2X2 U200 ( .A(n3794), .B(n3793), .Y(n3795) );
  AND2X2 U201 ( .A(n3789), .B(n3788), .Y(n3790) );
  AND2X2 U208 ( .A(n3781), .B(n3780), .Y(n3782) );
  AND2X2 U209 ( .A(n3769), .B(n3768), .Y(n3770) );
  AND2X2 U212 ( .A(n3761), .B(n3760), .Y(n3762) );
  AND2X2 U213 ( .A(n3756), .B(n3755), .Y(n3757) );
  AND2X2 U214 ( .A(n3748), .B(n3747), .Y(n3749) );
  OR2X2 U215 ( .A(n3744), .B(n3743), .Y(n3745) );
  AND2X2 U216 ( .A(n3738), .B(n3737), .Y(n3739) );
  AND2X2 U218 ( .A(n3732), .B(n3731), .Y(n3733) );
  AND2X2 U219 ( .A(n3727), .B(n3726), .Y(n3728) );
  OAI21X1 U817 ( .A(n4801), .B(n3191), .C(n4800), .Y(n3717) );
  AOI22X1 U818 ( .A(\data_in<8> ), .B(n4799), .C(\data_in<0> ), .D(n4798), .Y(
        n4800) );
  OAI21X1 U819 ( .A(n4801), .B(n3190), .C(n4797), .Y(n3716) );
  AOI22X1 U820 ( .A(\data_in<9> ), .B(n4799), .C(\data_in<1> ), .D(n4798), .Y(
        n4797) );
  OAI21X1 U821 ( .A(n4801), .B(n3189), .C(n4796), .Y(n3715) );
  AOI22X1 U822 ( .A(\data_in<10> ), .B(n4799), .C(\data_in<2> ), .D(n4798), 
        .Y(n4796) );
  OAI21X1 U823 ( .A(n4801), .B(n3188), .C(n4795), .Y(n3714) );
  AOI22X1 U824 ( .A(\data_in<11> ), .B(n4799), .C(\data_in<3> ), .D(n4798), 
        .Y(n4795) );
  OAI21X1 U825 ( .A(n4801), .B(n3187), .C(n4794), .Y(n3713) );
  AOI22X1 U826 ( .A(\data_in<12> ), .B(n4799), .C(\data_in<4> ), .D(n4798), 
        .Y(n4794) );
  OAI21X1 U827 ( .A(n4801), .B(n3186), .C(n4793), .Y(n3712) );
  AOI22X1 U828 ( .A(\data_in<13> ), .B(n4799), .C(\data_in<5> ), .D(n4798), 
        .Y(n4793) );
  OAI21X1 U829 ( .A(n4801), .B(n3185), .C(n4792), .Y(n3711) );
  AOI22X1 U830 ( .A(\data_in<14> ), .B(n4799), .C(\data_in<6> ), .D(n4798), 
        .Y(n4792) );
  OAI21X1 U831 ( .A(n4801), .B(n3184), .C(n4791), .Y(n3710) );
  AOI22X1 U832 ( .A(\data_in<15> ), .B(n4799), .C(\data_in<7> ), .D(n4798), 
        .Y(n4791) );
  OAI21X1 U833 ( .A(n350), .B(n4789), .C(n355), .Y(n4790) );
  OAI21X1 U834 ( .A(n2671), .B(n3183), .C(n4787), .Y(n3709) );
  AOI22X1 U835 ( .A(n4786), .B(\data_in<8> ), .C(n4785), .D(\data_in<0> ), .Y(
        n4787) );
  OAI21X1 U836 ( .A(n2671), .B(n3182), .C(n4784), .Y(n3708) );
  AOI22X1 U837 ( .A(n4786), .B(\data_in<9> ), .C(n4785), .D(\data_in<1> ), .Y(
        n4784) );
  OAI21X1 U838 ( .A(n2671), .B(n3181), .C(n4783), .Y(n3707) );
  AOI22X1 U839 ( .A(n4786), .B(\data_in<10> ), .C(n4785), .D(\data_in<2> ), 
        .Y(n4783) );
  OAI21X1 U840 ( .A(n2671), .B(n3180), .C(n4782), .Y(n3706) );
  AOI22X1 U841 ( .A(n4786), .B(\data_in<11> ), .C(n4785), .D(\data_in<3> ), 
        .Y(n4782) );
  OAI21X1 U842 ( .A(n2671), .B(n3179), .C(n4781), .Y(n3705) );
  AOI22X1 U843 ( .A(n4786), .B(\data_in<12> ), .C(n4785), .D(\data_in<4> ), 
        .Y(n4781) );
  OAI21X1 U844 ( .A(n2671), .B(n3178), .C(n4780), .Y(n3704) );
  AOI22X1 U845 ( .A(n4786), .B(\data_in<13> ), .C(n4785), .D(\data_in<5> ), 
        .Y(n4780) );
  OAI21X1 U846 ( .A(n2671), .B(n3177), .C(n4779), .Y(n3703) );
  AOI22X1 U847 ( .A(n4786), .B(\data_in<14> ), .C(n4785), .D(\data_in<6> ), 
        .Y(n4779) );
  OAI21X1 U848 ( .A(n2671), .B(n3176), .C(n4778), .Y(n3702) );
  AOI22X1 U849 ( .A(n4786), .B(\data_in<15> ), .C(n4785), .D(\data_in<7> ), 
        .Y(n4778) );
  AOI21X1 U850 ( .A(n355), .B(n460), .C(n2673), .Y(n4788) );
  OAI21X1 U851 ( .A(n2670), .B(n3175), .C(n4775), .Y(n3701) );
  AOI22X1 U852 ( .A(n4774), .B(\data_in<8> ), .C(n4773), .D(\data_in<0> ), .Y(
        n4775) );
  OAI21X1 U853 ( .A(n2670), .B(n3174), .C(n4772), .Y(n3700) );
  AOI22X1 U854 ( .A(n4774), .B(\data_in<9> ), .C(n4773), .D(\data_in<1> ), .Y(
        n4772) );
  OAI21X1 U855 ( .A(n2670), .B(n3173), .C(n4771), .Y(n3699) );
  AOI22X1 U856 ( .A(n4774), .B(\data_in<10> ), .C(n4773), .D(\data_in<2> ), 
        .Y(n4771) );
  OAI21X1 U857 ( .A(n2670), .B(n3172), .C(n4770), .Y(n3698) );
  AOI22X1 U858 ( .A(n4774), .B(\data_in<11> ), .C(n4773), .D(\data_in<3> ), 
        .Y(n4770) );
  OAI21X1 U859 ( .A(n2670), .B(n3171), .C(n4769), .Y(n3697) );
  AOI22X1 U860 ( .A(n4774), .B(\data_in<12> ), .C(n4773), .D(\data_in<4> ), 
        .Y(n4769) );
  OAI21X1 U861 ( .A(n2670), .B(n3170), .C(n4768), .Y(n3696) );
  AOI22X1 U862 ( .A(n4774), .B(\data_in<13> ), .C(n4773), .D(\data_in<5> ), 
        .Y(n4768) );
  OAI21X1 U863 ( .A(n2670), .B(n3169), .C(n4767), .Y(n3695) );
  AOI22X1 U864 ( .A(n4774), .B(\data_in<14> ), .C(n4773), .D(\data_in<6> ), 
        .Y(n4767) );
  OAI21X1 U865 ( .A(n2670), .B(n3168), .C(n4766), .Y(n3694) );
  AOI22X1 U866 ( .A(n4774), .B(\data_in<15> ), .C(n4773), .D(\data_in<7> ), 
        .Y(n4766) );
  AOI21X1 U867 ( .A(n460), .B(n455), .C(n2673), .Y(n4776) );
  OAI21X1 U868 ( .A(n2669), .B(n3167), .C(n4764), .Y(n3693) );
  AOI22X1 U869 ( .A(n4763), .B(\data_in<8> ), .C(n4762), .D(\data_in<0> ), .Y(
        n4764) );
  OAI21X1 U870 ( .A(n2669), .B(n3166), .C(n4761), .Y(n3692) );
  AOI22X1 U871 ( .A(n4763), .B(\data_in<9> ), .C(n4762), .D(\data_in<1> ), .Y(
        n4761) );
  OAI21X1 U872 ( .A(n2669), .B(n3165), .C(n4760), .Y(n3691) );
  AOI22X1 U873 ( .A(n4763), .B(\data_in<10> ), .C(n4762), .D(\data_in<2> ), 
        .Y(n4760) );
  OAI21X1 U874 ( .A(n2669), .B(n3164), .C(n4759), .Y(n3690) );
  AOI22X1 U875 ( .A(n4763), .B(\data_in<11> ), .C(n4762), .D(\data_in<3> ), 
        .Y(n4759) );
  OAI21X1 U876 ( .A(n2669), .B(n3163), .C(n4758), .Y(n3689) );
  AOI22X1 U877 ( .A(n4763), .B(\data_in<12> ), .C(n4762), .D(\data_in<4> ), 
        .Y(n4758) );
  OAI21X1 U878 ( .A(n2669), .B(n3162), .C(n4757), .Y(n3688) );
  AOI22X1 U879 ( .A(n4763), .B(\data_in<13> ), .C(n4762), .D(\data_in<5> ), 
        .Y(n4757) );
  OAI21X1 U880 ( .A(n2669), .B(n3161), .C(n4756), .Y(n3687) );
  AOI22X1 U881 ( .A(n4763), .B(\data_in<14> ), .C(n4762), .D(\data_in<6> ), 
        .Y(n4756) );
  OAI21X1 U882 ( .A(n2669), .B(n3160), .C(n4755), .Y(n3686) );
  AOI22X1 U883 ( .A(n4763), .B(\data_in<15> ), .C(n4762), .D(\data_in<7> ), 
        .Y(n4755) );
  AOI21X1 U884 ( .A(n455), .B(n458), .C(n2673), .Y(n4765) );
  OAI21X1 U885 ( .A(n2668), .B(n3159), .C(n4753), .Y(n3685) );
  AOI22X1 U886 ( .A(n4752), .B(\data_in<8> ), .C(n4751), .D(\data_in<0> ), .Y(
        n4753) );
  OAI21X1 U887 ( .A(n2668), .B(n3158), .C(n4750), .Y(n3684) );
  AOI22X1 U888 ( .A(n4752), .B(\data_in<9> ), .C(n4751), .D(\data_in<1> ), .Y(
        n4750) );
  OAI21X1 U889 ( .A(n2668), .B(n3157), .C(n4749), .Y(n3683) );
  AOI22X1 U890 ( .A(n4752), .B(\data_in<10> ), .C(n4751), .D(\data_in<2> ), 
        .Y(n4749) );
  OAI21X1 U891 ( .A(n2668), .B(n3156), .C(n4748), .Y(n3682) );
  AOI22X1 U892 ( .A(n4752), .B(\data_in<11> ), .C(n4751), .D(\data_in<3> ), 
        .Y(n4748) );
  OAI21X1 U893 ( .A(n2668), .B(n3155), .C(n4747), .Y(n3681) );
  AOI22X1 U894 ( .A(n4752), .B(\data_in<12> ), .C(n4751), .D(\data_in<4> ), 
        .Y(n4747) );
  OAI21X1 U895 ( .A(n2668), .B(n3154), .C(n4746), .Y(n3680) );
  AOI22X1 U896 ( .A(n4752), .B(\data_in<13> ), .C(n4751), .D(\data_in<5> ), 
        .Y(n4746) );
  OAI21X1 U897 ( .A(n2668), .B(n3153), .C(n4745), .Y(n3679) );
  AOI22X1 U898 ( .A(n4752), .B(\data_in<14> ), .C(n4751), .D(\data_in<6> ), 
        .Y(n4745) );
  OAI21X1 U899 ( .A(n2668), .B(n3152), .C(n4744), .Y(n3678) );
  AOI22X1 U900 ( .A(n4752), .B(\data_in<15> ), .C(n4751), .D(\data_in<7> ), 
        .Y(n4744) );
  AOI21X1 U901 ( .A(n458), .B(n451), .C(n2673), .Y(n4754) );
  OAI21X1 U902 ( .A(n2667), .B(n3151), .C(n4742), .Y(n3677) );
  AOI22X1 U903 ( .A(n4741), .B(\data_in<8> ), .C(n4740), .D(\data_in<0> ), .Y(
        n4742) );
  OAI21X1 U904 ( .A(n2667), .B(n3150), .C(n4739), .Y(n3676) );
  AOI22X1 U905 ( .A(n4741), .B(\data_in<9> ), .C(n4740), .D(\data_in<1> ), .Y(
        n4739) );
  OAI21X1 U906 ( .A(n2667), .B(n3149), .C(n4738), .Y(n3675) );
  AOI22X1 U907 ( .A(n4741), .B(\data_in<10> ), .C(n4740), .D(\data_in<2> ), 
        .Y(n4738) );
  OAI21X1 U908 ( .A(n2667), .B(n3148), .C(n4737), .Y(n3674) );
  AOI22X1 U909 ( .A(n4741), .B(\data_in<11> ), .C(n4740), .D(\data_in<3> ), 
        .Y(n4737) );
  OAI21X1 U910 ( .A(n2667), .B(n3147), .C(n4736), .Y(n3673) );
  AOI22X1 U911 ( .A(n4741), .B(\data_in<12> ), .C(n4740), .D(\data_in<4> ), 
        .Y(n4736) );
  OAI21X1 U912 ( .A(n2667), .B(n3146), .C(n4735), .Y(n3672) );
  AOI22X1 U913 ( .A(n4741), .B(\data_in<13> ), .C(n4740), .D(\data_in<5> ), 
        .Y(n4735) );
  OAI21X1 U914 ( .A(n2667), .B(n3145), .C(n4734), .Y(n3671) );
  AOI22X1 U915 ( .A(n4741), .B(\data_in<14> ), .C(n4740), .D(\data_in<6> ), 
        .Y(n4734) );
  OAI21X1 U916 ( .A(n2667), .B(n3144), .C(n4733), .Y(n3670) );
  AOI22X1 U917 ( .A(n4741), .B(\data_in<15> ), .C(n4740), .D(\data_in<7> ), 
        .Y(n4733) );
  AOI21X1 U918 ( .A(n451), .B(n454), .C(n2672), .Y(n4743) );
  OAI21X1 U919 ( .A(n2666), .B(n3143), .C(n4731), .Y(n3669) );
  AOI22X1 U920 ( .A(n4730), .B(\data_in<8> ), .C(n4729), .D(\data_in<0> ), .Y(
        n4731) );
  OAI21X1 U921 ( .A(n2666), .B(n3142), .C(n4728), .Y(n3668) );
  AOI22X1 U922 ( .A(n4730), .B(\data_in<9> ), .C(n4729), .D(\data_in<1> ), .Y(
        n4728) );
  OAI21X1 U923 ( .A(n2666), .B(n3141), .C(n4727), .Y(n3667) );
  AOI22X1 U924 ( .A(n4730), .B(\data_in<10> ), .C(n4729), .D(\data_in<2> ), 
        .Y(n4727) );
  OAI21X1 U925 ( .A(n2666), .B(n3140), .C(n4726), .Y(n3666) );
  AOI22X1 U926 ( .A(n4730), .B(\data_in<11> ), .C(n4729), .D(\data_in<3> ), 
        .Y(n4726) );
  OAI21X1 U927 ( .A(n2666), .B(n3139), .C(n4725), .Y(n3665) );
  AOI22X1 U928 ( .A(n4730), .B(\data_in<12> ), .C(n4729), .D(\data_in<4> ), 
        .Y(n4725) );
  OAI21X1 U929 ( .A(n2666), .B(n3138), .C(n4724), .Y(n3664) );
  AOI22X1 U930 ( .A(n4730), .B(\data_in<13> ), .C(n4729), .D(\data_in<5> ), 
        .Y(n4724) );
  OAI21X1 U931 ( .A(n2666), .B(n3137), .C(n4723), .Y(n3663) );
  AOI22X1 U932 ( .A(n4730), .B(\data_in<14> ), .C(n4729), .D(\data_in<6> ), 
        .Y(n4723) );
  OAI21X1 U933 ( .A(n2666), .B(n3136), .C(n4722), .Y(n3662) );
  AOI22X1 U934 ( .A(n4730), .B(\data_in<15> ), .C(n4729), .D(\data_in<7> ), 
        .Y(n4722) );
  AOI21X1 U935 ( .A(n454), .B(n447), .C(n2672), .Y(n4732) );
  OAI21X1 U936 ( .A(n2665), .B(n3135), .C(n4720), .Y(n3661) );
  AOI22X1 U937 ( .A(n4719), .B(\data_in<8> ), .C(n4718), .D(\data_in<0> ), .Y(
        n4720) );
  OAI21X1 U938 ( .A(n2665), .B(n3134), .C(n4717), .Y(n3660) );
  AOI22X1 U939 ( .A(n4719), .B(\data_in<9> ), .C(n4718), .D(\data_in<1> ), .Y(
        n4717) );
  OAI21X1 U940 ( .A(n2665), .B(n3133), .C(n4716), .Y(n3659) );
  AOI22X1 U941 ( .A(n4719), .B(\data_in<10> ), .C(n4718), .D(\data_in<2> ), 
        .Y(n4716) );
  OAI21X1 U942 ( .A(n2665), .B(n3132), .C(n4715), .Y(n3658) );
  AOI22X1 U943 ( .A(n4719), .B(\data_in<11> ), .C(n4718), .D(\data_in<3> ), 
        .Y(n4715) );
  OAI21X1 U944 ( .A(n2665), .B(n3131), .C(n4714), .Y(n3657) );
  AOI22X1 U945 ( .A(n4719), .B(\data_in<12> ), .C(n4718), .D(\data_in<4> ), 
        .Y(n4714) );
  OAI21X1 U946 ( .A(n2665), .B(n3130), .C(n4713), .Y(n3656) );
  AOI22X1 U947 ( .A(n4719), .B(\data_in<13> ), .C(n4718), .D(\data_in<5> ), 
        .Y(n4713) );
  OAI21X1 U948 ( .A(n2665), .B(n3129), .C(n4712), .Y(n3655) );
  AOI22X1 U949 ( .A(n4719), .B(\data_in<14> ), .C(n4718), .D(\data_in<6> ), 
        .Y(n4712) );
  OAI21X1 U950 ( .A(n2665), .B(n3128), .C(n4711), .Y(n3654) );
  AOI22X1 U951 ( .A(n4719), .B(\data_in<15> ), .C(n4718), .D(\data_in<7> ), 
        .Y(n4711) );
  AOI21X1 U952 ( .A(n447), .B(n450), .C(n2672), .Y(n4721) );
  OAI21X1 U953 ( .A(n2664), .B(n3127), .C(n4709), .Y(n3653) );
  AOI22X1 U954 ( .A(n4708), .B(\data_in<8> ), .C(n4707), .D(\data_in<0> ), .Y(
        n4709) );
  OAI21X1 U955 ( .A(n2664), .B(n3126), .C(n4706), .Y(n3652) );
  AOI22X1 U956 ( .A(n4708), .B(\data_in<9> ), .C(n4707), .D(\data_in<1> ), .Y(
        n4706) );
  OAI21X1 U957 ( .A(n2664), .B(n3125), .C(n4705), .Y(n3651) );
  AOI22X1 U958 ( .A(n4708), .B(\data_in<10> ), .C(n4707), .D(\data_in<2> ), 
        .Y(n4705) );
  OAI21X1 U959 ( .A(n2664), .B(n3124), .C(n4704), .Y(n3650) );
  AOI22X1 U960 ( .A(n4708), .B(\data_in<11> ), .C(n4707), .D(\data_in<3> ), 
        .Y(n4704) );
  OAI21X1 U961 ( .A(n2664), .B(n3123), .C(n4703), .Y(n3649) );
  AOI22X1 U962 ( .A(n4708), .B(\data_in<12> ), .C(n4707), .D(\data_in<4> ), 
        .Y(n4703) );
  OAI21X1 U963 ( .A(n2664), .B(n3122), .C(n4702), .Y(n3648) );
  AOI22X1 U964 ( .A(n4708), .B(\data_in<13> ), .C(n4707), .D(\data_in<5> ), 
        .Y(n4702) );
  OAI21X1 U965 ( .A(n2664), .B(n3121), .C(n4701), .Y(n3647) );
  AOI22X1 U966 ( .A(n4708), .B(\data_in<14> ), .C(n4707), .D(\data_in<6> ), 
        .Y(n4701) );
  OAI21X1 U967 ( .A(n2664), .B(n3120), .C(n4700), .Y(n3646) );
  AOI22X1 U968 ( .A(n4708), .B(\data_in<15> ), .C(n4707), .D(\data_in<7> ), 
        .Y(n4700) );
  AOI21X1 U969 ( .A(n450), .B(n474), .C(n2672), .Y(n4710) );
  OAI21X1 U970 ( .A(n2663), .B(n3119), .C(n4698), .Y(n3645) );
  AOI22X1 U971 ( .A(n4697), .B(\data_in<8> ), .C(n4696), .D(\data_in<0> ), .Y(
        n4698) );
  OAI21X1 U972 ( .A(n2663), .B(n3118), .C(n4695), .Y(n3644) );
  AOI22X1 U973 ( .A(n4697), .B(\data_in<9> ), .C(n4696), .D(\data_in<1> ), .Y(
        n4695) );
  OAI21X1 U974 ( .A(n2663), .B(n3117), .C(n4694), .Y(n3643) );
  AOI22X1 U975 ( .A(n4697), .B(\data_in<10> ), .C(n4696), .D(\data_in<2> ), 
        .Y(n4694) );
  OAI21X1 U976 ( .A(n2663), .B(n3116), .C(n4693), .Y(n3642) );
  AOI22X1 U977 ( .A(n4697), .B(\data_in<11> ), .C(n4696), .D(\data_in<3> ), 
        .Y(n4693) );
  OAI21X1 U978 ( .A(n2663), .B(n3115), .C(n4692), .Y(n3641) );
  AOI22X1 U979 ( .A(n4697), .B(\data_in<12> ), .C(n4696), .D(\data_in<4> ), 
        .Y(n4692) );
  OAI21X1 U980 ( .A(n2663), .B(n3114), .C(n4691), .Y(n3640) );
  AOI22X1 U981 ( .A(n4697), .B(\data_in<13> ), .C(n4696), .D(\data_in<5> ), 
        .Y(n4691) );
  OAI21X1 U982 ( .A(n2663), .B(n3113), .C(n4690), .Y(n3639) );
  AOI22X1 U983 ( .A(n4697), .B(\data_in<14> ), .C(n4696), .D(\data_in<6> ), 
        .Y(n4690) );
  OAI21X1 U984 ( .A(n2663), .B(n3112), .C(n4689), .Y(n3638) );
  AOI22X1 U985 ( .A(n4697), .B(\data_in<15> ), .C(n4696), .D(\data_in<7> ), 
        .Y(n4689) );
  AOI21X1 U986 ( .A(n474), .B(n476), .C(n2672), .Y(n4699) );
  OAI21X1 U987 ( .A(n2662), .B(n3111), .C(n4687), .Y(n3637) );
  AOI22X1 U988 ( .A(n4686), .B(\data_in<8> ), .C(n4685), .D(\data_in<0> ), .Y(
        n4687) );
  OAI21X1 U989 ( .A(n2662), .B(n3110), .C(n4684), .Y(n3636) );
  AOI22X1 U990 ( .A(n4686), .B(\data_in<9> ), .C(n4685), .D(\data_in<1> ), .Y(
        n4684) );
  OAI21X1 U991 ( .A(n2662), .B(n3109), .C(n4683), .Y(n3635) );
  AOI22X1 U992 ( .A(n4686), .B(\data_in<10> ), .C(n4685), .D(\data_in<2> ), 
        .Y(n4683) );
  OAI21X1 U993 ( .A(n2662), .B(n3108), .C(n4682), .Y(n3634) );
  AOI22X1 U994 ( .A(n4686), .B(\data_in<11> ), .C(n4685), .D(\data_in<3> ), 
        .Y(n4682) );
  OAI21X1 U995 ( .A(n2662), .B(n3107), .C(n4681), .Y(n3633) );
  AOI22X1 U996 ( .A(n4686), .B(\data_in<12> ), .C(n4685), .D(\data_in<4> ), 
        .Y(n4681) );
  OAI21X1 U997 ( .A(n2662), .B(n3106), .C(n4680), .Y(n3632) );
  AOI22X1 U998 ( .A(n4686), .B(\data_in<13> ), .C(n4685), .D(\data_in<5> ), 
        .Y(n4680) );
  OAI21X1 U999 ( .A(n2662), .B(n3105), .C(n4679), .Y(n3631) );
  AOI22X1 U1000 ( .A(n4686), .B(\data_in<14> ), .C(n4685), .D(\data_in<6> ), 
        .Y(n4679) );
  OAI21X1 U1001 ( .A(n2662), .B(n3104), .C(n4678), .Y(n3630) );
  AOI22X1 U1002 ( .A(n4686), .B(\data_in<15> ), .C(n4685), .D(\data_in<7> ), 
        .Y(n4678) );
  AOI21X1 U1003 ( .A(n476), .B(n470), .C(n2672), .Y(n4688) );
  OAI21X1 U1004 ( .A(n2661), .B(n3103), .C(n4676), .Y(n3629) );
  AOI22X1 U1005 ( .A(n4675), .B(\data_in<8> ), .C(n4674), .D(\data_in<0> ), 
        .Y(n4676) );
  OAI21X1 U1006 ( .A(n2661), .B(n3102), .C(n4673), .Y(n3628) );
  AOI22X1 U1007 ( .A(n4675), .B(\data_in<9> ), .C(n4674), .D(\data_in<1> ), 
        .Y(n4673) );
  OAI21X1 U1008 ( .A(n2661), .B(n3101), .C(n4672), .Y(n3627) );
  AOI22X1 U1009 ( .A(n4675), .B(\data_in<10> ), .C(n4674), .D(\data_in<2> ), 
        .Y(n4672) );
  OAI21X1 U1010 ( .A(n2661), .B(n3100), .C(n4671), .Y(n3626) );
  AOI22X1 U1011 ( .A(n4675), .B(\data_in<11> ), .C(n4674), .D(\data_in<3> ), 
        .Y(n4671) );
  OAI21X1 U1012 ( .A(n2661), .B(n3099), .C(n4670), .Y(n3625) );
  AOI22X1 U1013 ( .A(n4675), .B(\data_in<12> ), .C(n4674), .D(\data_in<4> ), 
        .Y(n4670) );
  OAI21X1 U1014 ( .A(n2661), .B(n3098), .C(n4669), .Y(n3624) );
  AOI22X1 U1015 ( .A(n4675), .B(\data_in<13> ), .C(n4674), .D(\data_in<5> ), 
        .Y(n4669) );
  OAI21X1 U1016 ( .A(n2661), .B(n3097), .C(n4668), .Y(n3623) );
  AOI22X1 U1017 ( .A(n4675), .B(\data_in<14> ), .C(n4674), .D(\data_in<6> ), 
        .Y(n4668) );
  OAI21X1 U1018 ( .A(n2661), .B(n3096), .C(n4667), .Y(n3622) );
  AOI22X1 U1019 ( .A(n4675), .B(\data_in<15> ), .C(n4674), .D(\data_in<7> ), 
        .Y(n4667) );
  AOI21X1 U1020 ( .A(n470), .B(n472), .C(n2672), .Y(n4677) );
  OAI21X1 U1021 ( .A(n2660), .B(n3095), .C(n4665), .Y(n3621) );
  AOI22X1 U1022 ( .A(n4664), .B(\data_in<8> ), .C(n4663), .D(\data_in<0> ), 
        .Y(n4665) );
  OAI21X1 U1023 ( .A(n2660), .B(n3094), .C(n4662), .Y(n3620) );
  AOI22X1 U1024 ( .A(n4664), .B(\data_in<9> ), .C(n4663), .D(\data_in<1> ), 
        .Y(n4662) );
  OAI21X1 U1025 ( .A(n2660), .B(n3093), .C(n4661), .Y(n3619) );
  AOI22X1 U1026 ( .A(n4664), .B(\data_in<10> ), .C(n4663), .D(\data_in<2> ), 
        .Y(n4661) );
  OAI21X1 U1027 ( .A(n2660), .B(n3092), .C(n4660), .Y(n3618) );
  AOI22X1 U1028 ( .A(n4664), .B(\data_in<11> ), .C(n4663), .D(\data_in<3> ), 
        .Y(n4660) );
  OAI21X1 U1029 ( .A(n2660), .B(n3091), .C(n4659), .Y(n3617) );
  AOI22X1 U1030 ( .A(n4664), .B(\data_in<12> ), .C(n4663), .D(\data_in<4> ), 
        .Y(n4659) );
  OAI21X1 U1031 ( .A(n2660), .B(n3090), .C(n4658), .Y(n3616) );
  AOI22X1 U1032 ( .A(n4664), .B(\data_in<13> ), .C(n4663), .D(\data_in<5> ), 
        .Y(n4658) );
  OAI21X1 U1033 ( .A(n2660), .B(n3089), .C(n4657), .Y(n3615) );
  AOI22X1 U1034 ( .A(n4664), .B(\data_in<14> ), .C(n4663), .D(\data_in<6> ), 
        .Y(n4657) );
  OAI21X1 U1035 ( .A(n2660), .B(n3088), .C(n4656), .Y(n3614) );
  AOI22X1 U1036 ( .A(n4664), .B(\data_in<15> ), .C(n4663), .D(\data_in<7> ), 
        .Y(n4656) );
  AOI21X1 U1037 ( .A(n472), .B(n466), .C(n2672), .Y(n4666) );
  OAI21X1 U1038 ( .A(n2659), .B(n3087), .C(n4654), .Y(n3613) );
  AOI22X1 U1039 ( .A(n4653), .B(\data_in<8> ), .C(n4652), .D(\data_in<0> ), 
        .Y(n4654) );
  OAI21X1 U1040 ( .A(n2659), .B(n3086), .C(n4651), .Y(n3612) );
  AOI22X1 U1041 ( .A(n4653), .B(\data_in<9> ), .C(n4652), .D(\data_in<1> ), 
        .Y(n4651) );
  OAI21X1 U1042 ( .A(n2659), .B(n3085), .C(n4650), .Y(n3611) );
  AOI22X1 U1043 ( .A(n4653), .B(\data_in<10> ), .C(n4652), .D(\data_in<2> ), 
        .Y(n4650) );
  OAI21X1 U1044 ( .A(n2659), .B(n3084), .C(n4649), .Y(n3610) );
  AOI22X1 U1045 ( .A(n4653), .B(\data_in<11> ), .C(n4652), .D(\data_in<3> ), 
        .Y(n4649) );
  OAI21X1 U1046 ( .A(n2659), .B(n3083), .C(n4648), .Y(n3609) );
  AOI22X1 U1047 ( .A(n4653), .B(\data_in<12> ), .C(n4652), .D(\data_in<4> ), 
        .Y(n4648) );
  OAI21X1 U1048 ( .A(n2659), .B(n3082), .C(n4647), .Y(n3608) );
  AOI22X1 U1049 ( .A(n4653), .B(\data_in<13> ), .C(n4652), .D(\data_in<5> ), 
        .Y(n4647) );
  OAI21X1 U1050 ( .A(n2659), .B(n3081), .C(n4646), .Y(n3607) );
  AOI22X1 U1051 ( .A(n4653), .B(\data_in<14> ), .C(n4652), .D(\data_in<6> ), 
        .Y(n4646) );
  OAI21X1 U1052 ( .A(n2659), .B(n3080), .C(n4645), .Y(n3606) );
  AOI22X1 U1053 ( .A(n4653), .B(\data_in<15> ), .C(n4652), .D(\data_in<7> ), 
        .Y(n4645) );
  AOI21X1 U1054 ( .A(n466), .B(n468), .C(n2672), .Y(n4655) );
  OAI21X1 U1055 ( .A(n2658), .B(n3079), .C(n4643), .Y(n3605) );
  AOI22X1 U1056 ( .A(n4642), .B(\data_in<8> ), .C(n4641), .D(\data_in<0> ), 
        .Y(n4643) );
  OAI21X1 U1057 ( .A(n2658), .B(n3078), .C(n4640), .Y(n3604) );
  AOI22X1 U1058 ( .A(n4642), .B(\data_in<9> ), .C(n4641), .D(\data_in<1> ), 
        .Y(n4640) );
  OAI21X1 U1059 ( .A(n2658), .B(n3077), .C(n4639), .Y(n3603) );
  AOI22X1 U1060 ( .A(n4642), .B(\data_in<10> ), .C(n4641), .D(\data_in<2> ), 
        .Y(n4639) );
  OAI21X1 U1061 ( .A(n2658), .B(n3076), .C(n4638), .Y(n3602) );
  AOI22X1 U1062 ( .A(n4642), .B(\data_in<11> ), .C(n4641), .D(\data_in<3> ), 
        .Y(n4638) );
  OAI21X1 U1063 ( .A(n2658), .B(n3075), .C(n4637), .Y(n3601) );
  AOI22X1 U1064 ( .A(n4642), .B(\data_in<12> ), .C(n4641), .D(\data_in<4> ), 
        .Y(n4637) );
  OAI21X1 U1065 ( .A(n2658), .B(n3074), .C(n4636), .Y(n3600) );
  AOI22X1 U1066 ( .A(n4642), .B(\data_in<13> ), .C(n4641), .D(\data_in<5> ), 
        .Y(n4636) );
  OAI21X1 U1067 ( .A(n2658), .B(n3073), .C(n4635), .Y(n3599) );
  AOI22X1 U1068 ( .A(n4642), .B(\data_in<14> ), .C(n4641), .D(\data_in<6> ), 
        .Y(n4635) );
  OAI21X1 U1069 ( .A(n2658), .B(n3072), .C(n4634), .Y(n3598) );
  AOI22X1 U1070 ( .A(n4642), .B(\data_in<15> ), .C(n4641), .D(\data_in<7> ), 
        .Y(n4634) );
  AOI21X1 U1071 ( .A(n468), .B(n462), .C(n2672), .Y(n4644) );
  OAI21X1 U1072 ( .A(n2657), .B(n3071), .C(n4632), .Y(n3597) );
  AOI22X1 U1073 ( .A(n4631), .B(\data_in<8> ), .C(n4630), .D(\data_in<0> ), 
        .Y(n4632) );
  OAI21X1 U1074 ( .A(n2657), .B(n3070), .C(n4629), .Y(n3596) );
  AOI22X1 U1075 ( .A(n4631), .B(\data_in<9> ), .C(n4630), .D(\data_in<1> ), 
        .Y(n4629) );
  OAI21X1 U1076 ( .A(n2657), .B(n3069), .C(n4628), .Y(n3595) );
  AOI22X1 U1077 ( .A(n4631), .B(\data_in<10> ), .C(n4630), .D(\data_in<2> ), 
        .Y(n4628) );
  OAI21X1 U1078 ( .A(n2657), .B(n3068), .C(n4627), .Y(n3594) );
  AOI22X1 U1079 ( .A(n4631), .B(\data_in<11> ), .C(n4630), .D(\data_in<3> ), 
        .Y(n4627) );
  OAI21X1 U1080 ( .A(n2657), .B(n3067), .C(n4626), .Y(n3593) );
  AOI22X1 U1081 ( .A(n4631), .B(\data_in<12> ), .C(n4630), .D(\data_in<4> ), 
        .Y(n4626) );
  OAI21X1 U1082 ( .A(n2657), .B(n3066), .C(n4625), .Y(n3592) );
  AOI22X1 U1083 ( .A(n4631), .B(\data_in<13> ), .C(n4630), .D(\data_in<5> ), 
        .Y(n4625) );
  OAI21X1 U1084 ( .A(n2657), .B(n3065), .C(n4624), .Y(n3591) );
  AOI22X1 U1085 ( .A(n4631), .B(\data_in<14> ), .C(n4630), .D(\data_in<6> ), 
        .Y(n4624) );
  OAI21X1 U1086 ( .A(n2657), .B(n3064), .C(n4623), .Y(n3590) );
  AOI22X1 U1087 ( .A(n4631), .B(\data_in<15> ), .C(n4630), .D(\data_in<7> ), 
        .Y(n4623) );
  AOI21X1 U1088 ( .A(n462), .B(n464), .C(n2672), .Y(n4633) );
  OAI21X1 U1089 ( .A(n2656), .B(n3063), .C(n4621), .Y(n3589) );
  AOI22X1 U1090 ( .A(n4620), .B(\data_in<8> ), .C(n4619), .D(\data_in<0> ), 
        .Y(n4621) );
  OAI21X1 U1091 ( .A(n2656), .B(n3062), .C(n4618), .Y(n3588) );
  AOI22X1 U1092 ( .A(n4620), .B(\data_in<9> ), .C(n4619), .D(\data_in<1> ), 
        .Y(n4618) );
  OAI21X1 U1093 ( .A(n2656), .B(n3061), .C(n4617), .Y(n3587) );
  AOI22X1 U1094 ( .A(n4620), .B(\data_in<10> ), .C(n4619), .D(\data_in<2> ), 
        .Y(n4617) );
  OAI21X1 U1095 ( .A(n2656), .B(n3060), .C(n4616), .Y(n3586) );
  AOI22X1 U1096 ( .A(n4620), .B(\data_in<11> ), .C(n4619), .D(\data_in<3> ), 
        .Y(n4616) );
  OAI21X1 U1097 ( .A(n2656), .B(n3059), .C(n4615), .Y(n3585) );
  AOI22X1 U1098 ( .A(n4620), .B(\data_in<12> ), .C(n4619), .D(\data_in<4> ), 
        .Y(n4615) );
  OAI21X1 U1099 ( .A(n2656), .B(n3058), .C(n4614), .Y(n3584) );
  AOI22X1 U1100 ( .A(n4620), .B(\data_in<13> ), .C(n4619), .D(\data_in<5> ), 
        .Y(n4614) );
  OAI21X1 U1101 ( .A(n2656), .B(n3057), .C(n4613), .Y(n3583) );
  AOI22X1 U1102 ( .A(n4620), .B(\data_in<14> ), .C(n4619), .D(\data_in<6> ), 
        .Y(n4613) );
  OAI21X1 U1103 ( .A(n2656), .B(n3056), .C(n4612), .Y(n3582) );
  AOI22X1 U1104 ( .A(n4620), .B(\data_in<15> ), .C(n4619), .D(\data_in<7> ), 
        .Y(n4612) );
  AOI21X1 U1105 ( .A(n464), .B(n428), .C(n2672), .Y(n4622) );
  OAI21X1 U1106 ( .A(n2655), .B(n3055), .C(n4610), .Y(n3581) );
  AOI22X1 U1107 ( .A(n4609), .B(\data_in<8> ), .C(n4608), .D(\data_in<0> ), 
        .Y(n4610) );
  OAI21X1 U1108 ( .A(n2655), .B(n3054), .C(n4607), .Y(n3580) );
  AOI22X1 U1109 ( .A(n4609), .B(\data_in<9> ), .C(n4608), .D(\data_in<1> ), 
        .Y(n4607) );
  OAI21X1 U1110 ( .A(n2655), .B(n3053), .C(n4606), .Y(n3579) );
  AOI22X1 U1111 ( .A(n4609), .B(\data_in<10> ), .C(n4608), .D(\data_in<2> ), 
        .Y(n4606) );
  OAI21X1 U1112 ( .A(n2655), .B(n3052), .C(n4605), .Y(n3578) );
  AOI22X1 U1113 ( .A(n4609), .B(\data_in<11> ), .C(n4608), .D(\data_in<3> ), 
        .Y(n4605) );
  OAI21X1 U1114 ( .A(n2655), .B(n3051), .C(n4604), .Y(n3577) );
  AOI22X1 U1115 ( .A(n4609), .B(\data_in<12> ), .C(n4608), .D(\data_in<4> ), 
        .Y(n4604) );
  OAI21X1 U1116 ( .A(n2655), .B(n3050), .C(n4603), .Y(n3576) );
  AOI22X1 U1117 ( .A(n4609), .B(\data_in<13> ), .C(n4608), .D(\data_in<5> ), 
        .Y(n4603) );
  OAI21X1 U1118 ( .A(n2655), .B(n3049), .C(n4602), .Y(n3575) );
  AOI22X1 U1119 ( .A(n4609), .B(\data_in<14> ), .C(n4608), .D(\data_in<6> ), 
        .Y(n4602) );
  OAI21X1 U1120 ( .A(n2655), .B(n3048), .C(n4601), .Y(n3574) );
  AOI22X1 U1121 ( .A(n4609), .B(\data_in<15> ), .C(n4608), .D(\data_in<7> ), 
        .Y(n4601) );
  AOI21X1 U1122 ( .A(n428), .B(n430), .C(n2672), .Y(n4611) );
  OAI21X1 U1123 ( .A(n2654), .B(n3047), .C(n4599), .Y(n3573) );
  AOI22X1 U1124 ( .A(n4598), .B(\data_in<8> ), .C(n4597), .D(\data_in<0> ), 
        .Y(n4599) );
  OAI21X1 U1125 ( .A(n2654), .B(n3046), .C(n4596), .Y(n3572) );
  AOI22X1 U1126 ( .A(n4598), .B(\data_in<9> ), .C(n4597), .D(\data_in<1> ), 
        .Y(n4596) );
  OAI21X1 U1127 ( .A(n2654), .B(n3045), .C(n4595), .Y(n3571) );
  AOI22X1 U1128 ( .A(n4598), .B(\data_in<10> ), .C(n4597), .D(\data_in<2> ), 
        .Y(n4595) );
  OAI21X1 U1129 ( .A(n2654), .B(n3044), .C(n4594), .Y(n3570) );
  AOI22X1 U1130 ( .A(n4598), .B(\data_in<11> ), .C(n4597), .D(\data_in<3> ), 
        .Y(n4594) );
  OAI21X1 U1131 ( .A(n2654), .B(n3043), .C(n4593), .Y(n3569) );
  AOI22X1 U1132 ( .A(n4598), .B(\data_in<12> ), .C(n4597), .D(\data_in<4> ), 
        .Y(n4593) );
  OAI21X1 U1133 ( .A(n2654), .B(n3042), .C(n4592), .Y(n3568) );
  AOI22X1 U1134 ( .A(n4598), .B(\data_in<13> ), .C(n4597), .D(\data_in<5> ), 
        .Y(n4592) );
  OAI21X1 U1135 ( .A(n2654), .B(n3041), .C(n4591), .Y(n3567) );
  AOI22X1 U1136 ( .A(n4598), .B(\data_in<14> ), .C(n4597), .D(\data_in<6> ), 
        .Y(n4591) );
  OAI21X1 U1137 ( .A(n2654), .B(n3040), .C(n4590), .Y(n3566) );
  AOI22X1 U1138 ( .A(n4598), .B(\data_in<15> ), .C(n4597), .D(\data_in<7> ), 
        .Y(n4590) );
  AOI21X1 U1139 ( .A(n430), .B(n424), .C(n2672), .Y(n4600) );
  OAI21X1 U1140 ( .A(n2653), .B(n3039), .C(n4588), .Y(n3565) );
  AOI22X1 U1141 ( .A(n4587), .B(\data_in<8> ), .C(n4586), .D(\data_in<0> ), 
        .Y(n4588) );
  OAI21X1 U1142 ( .A(n2653), .B(n3038), .C(n4585), .Y(n3564) );
  AOI22X1 U1143 ( .A(n4587), .B(\data_in<9> ), .C(n4586), .D(\data_in<1> ), 
        .Y(n4585) );
  OAI21X1 U1144 ( .A(n2653), .B(n3037), .C(n4584), .Y(n3563) );
  AOI22X1 U1145 ( .A(n4587), .B(\data_in<10> ), .C(n4586), .D(\data_in<2> ), 
        .Y(n4584) );
  OAI21X1 U1146 ( .A(n2653), .B(n3036), .C(n4583), .Y(n3562) );
  AOI22X1 U1147 ( .A(n4587), .B(\data_in<11> ), .C(n4586), .D(\data_in<3> ), 
        .Y(n4583) );
  OAI21X1 U1148 ( .A(n2653), .B(n3035), .C(n4582), .Y(n3561) );
  AOI22X1 U1149 ( .A(n4587), .B(\data_in<12> ), .C(n4586), .D(\data_in<4> ), 
        .Y(n4582) );
  OAI21X1 U1150 ( .A(n2653), .B(n3034), .C(n4581), .Y(n3560) );
  AOI22X1 U1151 ( .A(n4587), .B(\data_in<13> ), .C(n4586), .D(\data_in<5> ), 
        .Y(n4581) );
  OAI21X1 U1152 ( .A(n2653), .B(n3033), .C(n4580), .Y(n3559) );
  AOI22X1 U1153 ( .A(n4587), .B(\data_in<14> ), .C(n4586), .D(\data_in<6> ), 
        .Y(n4580) );
  OAI21X1 U1154 ( .A(n2653), .B(n3032), .C(n4579), .Y(n3558) );
  AOI22X1 U1155 ( .A(n4587), .B(\data_in<15> ), .C(n4586), .D(\data_in<7> ), 
        .Y(n4579) );
  AOI21X1 U1156 ( .A(n424), .B(n426), .C(n2672), .Y(n4589) );
  OAI21X1 U1157 ( .A(n2652), .B(n3031), .C(n4577), .Y(n3557) );
  AOI22X1 U1158 ( .A(n4576), .B(\data_in<8> ), .C(n4575), .D(\data_in<0> ), 
        .Y(n4577) );
  OAI21X1 U1159 ( .A(n2652), .B(n3030), .C(n4574), .Y(n3556) );
  AOI22X1 U1160 ( .A(n4576), .B(\data_in<9> ), .C(n4575), .D(\data_in<1> ), 
        .Y(n4574) );
  OAI21X1 U1161 ( .A(n2652), .B(n3029), .C(n4573), .Y(n3555) );
  AOI22X1 U1162 ( .A(n4576), .B(\data_in<10> ), .C(n4575), .D(\data_in<2> ), 
        .Y(n4573) );
  OAI21X1 U1163 ( .A(n2652), .B(n3028), .C(n4572), .Y(n3554) );
  AOI22X1 U1164 ( .A(n4576), .B(\data_in<11> ), .C(n4575), .D(\data_in<3> ), 
        .Y(n4572) );
  OAI21X1 U1165 ( .A(n2652), .B(n3027), .C(n4571), .Y(n3553) );
  AOI22X1 U1166 ( .A(n4576), .B(\data_in<12> ), .C(n4575), .D(\data_in<4> ), 
        .Y(n4571) );
  OAI21X1 U1167 ( .A(n2652), .B(n3026), .C(n4570), .Y(n3552) );
  AOI22X1 U1168 ( .A(n4576), .B(\data_in<13> ), .C(n4575), .D(\data_in<5> ), 
        .Y(n4570) );
  OAI21X1 U1169 ( .A(n2652), .B(n3025), .C(n4569), .Y(n3551) );
  AOI22X1 U1170 ( .A(n4576), .B(\data_in<14> ), .C(n4575), .D(\data_in<6> ), 
        .Y(n4569) );
  OAI21X1 U1171 ( .A(n2652), .B(n3024), .C(n4568), .Y(n3550) );
  AOI22X1 U1172 ( .A(n4576), .B(\data_in<15> ), .C(n4575), .D(\data_in<7> ), 
        .Y(n4568) );
  AOI21X1 U1173 ( .A(n426), .B(n420), .C(n2672), .Y(n4578) );
  OAI21X1 U1174 ( .A(n2651), .B(n3023), .C(n4566), .Y(n3549) );
  AOI22X1 U1175 ( .A(n4565), .B(\data_in<8> ), .C(n4564), .D(\data_in<0> ), 
        .Y(n4566) );
  OAI21X1 U1176 ( .A(n2651), .B(n3022), .C(n4563), .Y(n3548) );
  AOI22X1 U1177 ( .A(n4565), .B(\data_in<9> ), .C(n4564), .D(\data_in<1> ), 
        .Y(n4563) );
  OAI21X1 U1178 ( .A(n2651), .B(n3021), .C(n4562), .Y(n3547) );
  AOI22X1 U1179 ( .A(n4565), .B(\data_in<10> ), .C(n4564), .D(\data_in<2> ), 
        .Y(n4562) );
  OAI21X1 U1180 ( .A(n2651), .B(n3020), .C(n4561), .Y(n3546) );
  AOI22X1 U1181 ( .A(n4565), .B(\data_in<11> ), .C(n4564), .D(\data_in<3> ), 
        .Y(n4561) );
  OAI21X1 U1182 ( .A(n2651), .B(n3019), .C(n4560), .Y(n3545) );
  AOI22X1 U1183 ( .A(n4565), .B(\data_in<12> ), .C(n4564), .D(\data_in<4> ), 
        .Y(n4560) );
  OAI21X1 U1184 ( .A(n2651), .B(n3018), .C(n4559), .Y(n3544) );
  AOI22X1 U1185 ( .A(n4565), .B(\data_in<13> ), .C(n4564), .D(\data_in<5> ), 
        .Y(n4559) );
  OAI21X1 U1186 ( .A(n2651), .B(n3017), .C(n4558), .Y(n3543) );
  AOI22X1 U1187 ( .A(n4565), .B(\data_in<14> ), .C(n4564), .D(\data_in<6> ), 
        .Y(n4558) );
  OAI21X1 U1188 ( .A(n2651), .B(n3016), .C(n4557), .Y(n3542) );
  AOI22X1 U1189 ( .A(n4565), .B(\data_in<15> ), .C(n4564), .D(\data_in<7> ), 
        .Y(n4557) );
  AOI21X1 U1190 ( .A(n420), .B(n422), .C(n2673), .Y(n4567) );
  OAI21X1 U1191 ( .A(n2650), .B(n3015), .C(n4555), .Y(n3541) );
  AOI22X1 U1192 ( .A(n4554), .B(\data_in<8> ), .C(n4553), .D(\data_in<0> ), 
        .Y(n4555) );
  OAI21X1 U1193 ( .A(n2650), .B(n3014), .C(n4552), .Y(n3540) );
  AOI22X1 U1194 ( .A(n4554), .B(\data_in<9> ), .C(n4553), .D(\data_in<1> ), 
        .Y(n4552) );
  OAI21X1 U1195 ( .A(n2650), .B(n3013), .C(n4551), .Y(n3539) );
  AOI22X1 U1196 ( .A(n4554), .B(\data_in<10> ), .C(n4553), .D(\data_in<2> ), 
        .Y(n4551) );
  OAI21X1 U1197 ( .A(n2650), .B(n3012), .C(n4550), .Y(n3538) );
  AOI22X1 U1198 ( .A(n4554), .B(\data_in<11> ), .C(n4553), .D(\data_in<3> ), 
        .Y(n4550) );
  OAI21X1 U1199 ( .A(n2650), .B(n3011), .C(n4549), .Y(n3537) );
  AOI22X1 U1200 ( .A(n4554), .B(\data_in<12> ), .C(n4553), .D(\data_in<4> ), 
        .Y(n4549) );
  OAI21X1 U1201 ( .A(n2650), .B(n3010), .C(n4548), .Y(n3536) );
  AOI22X1 U1202 ( .A(n4554), .B(\data_in<13> ), .C(n4553), .D(\data_in<5> ), 
        .Y(n4548) );
  OAI21X1 U1203 ( .A(n2650), .B(n3009), .C(n4547), .Y(n3535) );
  AOI22X1 U1204 ( .A(n4554), .B(\data_in<14> ), .C(n4553), .D(\data_in<6> ), 
        .Y(n4547) );
  OAI21X1 U1205 ( .A(n2650), .B(n3008), .C(n4546), .Y(n3534) );
  AOI22X1 U1206 ( .A(n4554), .B(\data_in<15> ), .C(n4553), .D(\data_in<7> ), 
        .Y(n4546) );
  AOI21X1 U1207 ( .A(n422), .B(n416), .C(n2673), .Y(n4556) );
  OAI21X1 U1208 ( .A(n2649), .B(n3007), .C(n4544), .Y(n3533) );
  AOI22X1 U1209 ( .A(n4543), .B(\data_in<8> ), .C(n4542), .D(\data_in<0> ), 
        .Y(n4544) );
  OAI21X1 U1210 ( .A(n2649), .B(n3006), .C(n4541), .Y(n3532) );
  AOI22X1 U1211 ( .A(n4543), .B(\data_in<9> ), .C(n4542), .D(\data_in<1> ), 
        .Y(n4541) );
  OAI21X1 U1212 ( .A(n2649), .B(n3005), .C(n4540), .Y(n3531) );
  AOI22X1 U1213 ( .A(n4543), .B(\data_in<10> ), .C(n4542), .D(\data_in<2> ), 
        .Y(n4540) );
  OAI21X1 U1214 ( .A(n2649), .B(n3004), .C(n4539), .Y(n3530) );
  AOI22X1 U1215 ( .A(n4543), .B(\data_in<11> ), .C(n4542), .D(\data_in<3> ), 
        .Y(n4539) );
  OAI21X1 U1216 ( .A(n2649), .B(n3003), .C(n4538), .Y(n3529) );
  AOI22X1 U1217 ( .A(n4543), .B(\data_in<12> ), .C(n4542), .D(\data_in<4> ), 
        .Y(n4538) );
  OAI21X1 U1218 ( .A(n2649), .B(n3002), .C(n4537), .Y(n3528) );
  AOI22X1 U1219 ( .A(n4543), .B(\data_in<13> ), .C(n4542), .D(\data_in<5> ), 
        .Y(n4537) );
  OAI21X1 U1220 ( .A(n2649), .B(n3001), .C(n4536), .Y(n3527) );
  AOI22X1 U1221 ( .A(n4543), .B(\data_in<14> ), .C(n4542), .D(\data_in<6> ), 
        .Y(n4536) );
  OAI21X1 U1222 ( .A(n2649), .B(n3000), .C(n4535), .Y(n3526) );
  AOI22X1 U1223 ( .A(n4543), .B(\data_in<15> ), .C(n4542), .D(\data_in<7> ), 
        .Y(n4535) );
  AOI21X1 U1224 ( .A(n416), .B(n418), .C(n2673), .Y(n4545) );
  OAI21X1 U1225 ( .A(n2648), .B(n2999), .C(n4533), .Y(n3525) );
  AOI22X1 U1226 ( .A(n4532), .B(\data_in<8> ), .C(n4531), .D(\data_in<0> ), 
        .Y(n4533) );
  OAI21X1 U1227 ( .A(n2648), .B(n2998), .C(n4530), .Y(n3524) );
  AOI22X1 U1228 ( .A(n4532), .B(\data_in<9> ), .C(n4531), .D(\data_in<1> ), 
        .Y(n4530) );
  OAI21X1 U1229 ( .A(n2648), .B(n2997), .C(n4529), .Y(n3523) );
  AOI22X1 U1230 ( .A(n4532), .B(\data_in<10> ), .C(n4531), .D(\data_in<2> ), 
        .Y(n4529) );
  OAI21X1 U1231 ( .A(n2648), .B(n2996), .C(n4528), .Y(n3522) );
  AOI22X1 U1232 ( .A(n4532), .B(\data_in<11> ), .C(n4531), .D(\data_in<3> ), 
        .Y(n4528) );
  OAI21X1 U1233 ( .A(n2648), .B(n2995), .C(n4527), .Y(n3521) );
  AOI22X1 U1234 ( .A(n4532), .B(\data_in<12> ), .C(n4531), .D(\data_in<4> ), 
        .Y(n4527) );
  OAI21X1 U1235 ( .A(n2648), .B(n2994), .C(n4526), .Y(n3520) );
  AOI22X1 U1236 ( .A(n4532), .B(\data_in<13> ), .C(n4531), .D(\data_in<5> ), 
        .Y(n4526) );
  OAI21X1 U1237 ( .A(n2648), .B(n2993), .C(n4525), .Y(n3519) );
  AOI22X1 U1238 ( .A(n4532), .B(\data_in<14> ), .C(n4531), .D(\data_in<6> ), 
        .Y(n4525) );
  OAI21X1 U1239 ( .A(n2648), .B(n2992), .C(n4524), .Y(n3518) );
  AOI22X1 U1240 ( .A(n4532), .B(\data_in<15> ), .C(n4531), .D(\data_in<7> ), 
        .Y(n4524) );
  AOI21X1 U1241 ( .A(n418), .B(n444), .C(n2673), .Y(n4534) );
  OAI21X1 U1242 ( .A(n2647), .B(n2991), .C(n4522), .Y(n3517) );
  AOI22X1 U1243 ( .A(n4521), .B(\data_in<8> ), .C(n4520), .D(\data_in<0> ), 
        .Y(n4522) );
  OAI21X1 U1244 ( .A(n2647), .B(n2990), .C(n4519), .Y(n3516) );
  AOI22X1 U1245 ( .A(n4521), .B(\data_in<9> ), .C(n4520), .D(\data_in<1> ), 
        .Y(n4519) );
  OAI21X1 U1246 ( .A(n2647), .B(n2989), .C(n4518), .Y(n3515) );
  AOI22X1 U1247 ( .A(n4521), .B(\data_in<10> ), .C(n4520), .D(\data_in<2> ), 
        .Y(n4518) );
  OAI21X1 U1248 ( .A(n2647), .B(n2988), .C(n4517), .Y(n3514) );
  AOI22X1 U1249 ( .A(n4521), .B(\data_in<11> ), .C(n4520), .D(\data_in<3> ), 
        .Y(n4517) );
  OAI21X1 U1250 ( .A(n2647), .B(n2987), .C(n4516), .Y(n3513) );
  AOI22X1 U1251 ( .A(n4521), .B(\data_in<12> ), .C(n4520), .D(\data_in<4> ), 
        .Y(n4516) );
  OAI21X1 U1252 ( .A(n2647), .B(n2986), .C(n4515), .Y(n3512) );
  AOI22X1 U1253 ( .A(n4521), .B(\data_in<13> ), .C(n4520), .D(\data_in<5> ), 
        .Y(n4515) );
  OAI21X1 U1254 ( .A(n2647), .B(n2985), .C(n4514), .Y(n3511) );
  AOI22X1 U1255 ( .A(n4521), .B(\data_in<14> ), .C(n4520), .D(\data_in<6> ), 
        .Y(n4514) );
  OAI21X1 U1256 ( .A(n2647), .B(n2984), .C(n4513), .Y(n3510) );
  AOI22X1 U1257 ( .A(n4521), .B(\data_in<15> ), .C(n4520), .D(\data_in<7> ), 
        .Y(n4513) );
  AOI21X1 U1258 ( .A(n444), .B(n445), .C(n2673), .Y(n4523) );
  OAI21X1 U1259 ( .A(n2646), .B(n2983), .C(n4511), .Y(n3509) );
  AOI22X1 U1260 ( .A(n4510), .B(\data_in<8> ), .C(n4509), .D(\data_in<0> ), 
        .Y(n4511) );
  OAI21X1 U1261 ( .A(n2646), .B(n2982), .C(n4508), .Y(n3508) );
  AOI22X1 U1262 ( .A(n4510), .B(\data_in<9> ), .C(n4509), .D(\data_in<1> ), 
        .Y(n4508) );
  OAI21X1 U1263 ( .A(n2646), .B(n2981), .C(n4507), .Y(n3507) );
  AOI22X1 U1264 ( .A(n4510), .B(\data_in<10> ), .C(n4509), .D(\data_in<2> ), 
        .Y(n4507) );
  OAI21X1 U1265 ( .A(n2646), .B(n2980), .C(n4506), .Y(n3506) );
  AOI22X1 U1266 ( .A(n4510), .B(\data_in<11> ), .C(n4509), .D(\data_in<3> ), 
        .Y(n4506) );
  OAI21X1 U1267 ( .A(n2646), .B(n2979), .C(n4505), .Y(n3505) );
  AOI22X1 U1268 ( .A(n4510), .B(\data_in<12> ), .C(n4509), .D(\data_in<4> ), 
        .Y(n4505) );
  OAI21X1 U1269 ( .A(n2646), .B(n2978), .C(n4504), .Y(n3504) );
  AOI22X1 U1270 ( .A(n4510), .B(\data_in<13> ), .C(n4509), .D(\data_in<5> ), 
        .Y(n4504) );
  OAI21X1 U1271 ( .A(n2646), .B(n2977), .C(n4503), .Y(n3503) );
  AOI22X1 U1272 ( .A(n4510), .B(\data_in<14> ), .C(n4509), .D(\data_in<6> ), 
        .Y(n4503) );
  OAI21X1 U1273 ( .A(n2646), .B(n2976), .C(n4502), .Y(n3502) );
  AOI22X1 U1274 ( .A(n4510), .B(\data_in<15> ), .C(n4509), .D(\data_in<7> ), 
        .Y(n4502) );
  AOI21X1 U1275 ( .A(n445), .B(n440), .C(n2673), .Y(n4512) );
  OAI21X1 U1276 ( .A(n2645), .B(n2975), .C(n4500), .Y(n3501) );
  AOI22X1 U1277 ( .A(n4499), .B(\data_in<8> ), .C(n4498), .D(\data_in<0> ), 
        .Y(n4500) );
  OAI21X1 U1278 ( .A(n2645), .B(n2974), .C(n4497), .Y(n3500) );
  AOI22X1 U1279 ( .A(n4499), .B(\data_in<9> ), .C(n4498), .D(\data_in<1> ), 
        .Y(n4497) );
  OAI21X1 U1280 ( .A(n2645), .B(n2973), .C(n4496), .Y(n3499) );
  AOI22X1 U1281 ( .A(n4499), .B(\data_in<10> ), .C(n4498), .D(\data_in<2> ), 
        .Y(n4496) );
  OAI21X1 U1282 ( .A(n2645), .B(n2972), .C(n4495), .Y(n3498) );
  AOI22X1 U1283 ( .A(n4499), .B(\data_in<11> ), .C(n4498), .D(\data_in<3> ), 
        .Y(n4495) );
  OAI21X1 U1284 ( .A(n2645), .B(n2971), .C(n4494), .Y(n3497) );
  AOI22X1 U1285 ( .A(n4499), .B(\data_in<12> ), .C(n4498), .D(\data_in<4> ), 
        .Y(n4494) );
  OAI21X1 U1286 ( .A(n2645), .B(n2970), .C(n4493), .Y(n3496) );
  AOI22X1 U1287 ( .A(n4499), .B(\data_in<13> ), .C(n4498), .D(\data_in<5> ), 
        .Y(n4493) );
  OAI21X1 U1288 ( .A(n2645), .B(n2969), .C(n4492), .Y(n3495) );
  AOI22X1 U1289 ( .A(n4499), .B(\data_in<14> ), .C(n4498), .D(\data_in<6> ), 
        .Y(n4492) );
  OAI21X1 U1290 ( .A(n2645), .B(n2968), .C(n4491), .Y(n3494) );
  AOI22X1 U1291 ( .A(n4499), .B(\data_in<15> ), .C(n4498), .D(\data_in<7> ), 
        .Y(n4491) );
  AOI21X1 U1292 ( .A(n440), .B(n441), .C(n2673), .Y(n4501) );
  OAI21X1 U1293 ( .A(n2644), .B(n2967), .C(n4489), .Y(n3493) );
  AOI22X1 U1294 ( .A(n4488), .B(\data_in<8> ), .C(n4487), .D(\data_in<0> ), 
        .Y(n4489) );
  OAI21X1 U1295 ( .A(n2644), .B(n2966), .C(n4486), .Y(n3492) );
  AOI22X1 U1296 ( .A(n4488), .B(\data_in<9> ), .C(n4487), .D(\data_in<1> ), 
        .Y(n4486) );
  OAI21X1 U1297 ( .A(n2644), .B(n2965), .C(n4485), .Y(n3491) );
  AOI22X1 U1298 ( .A(n4488), .B(\data_in<10> ), .C(n4487), .D(\data_in<2> ), 
        .Y(n4485) );
  OAI21X1 U1299 ( .A(n2644), .B(n2964), .C(n4484), .Y(n3490) );
  AOI22X1 U1300 ( .A(n4488), .B(\data_in<11> ), .C(n4487), .D(\data_in<3> ), 
        .Y(n4484) );
  OAI21X1 U1301 ( .A(n2644), .B(n2963), .C(n4483), .Y(n3489) );
  AOI22X1 U1302 ( .A(n4488), .B(\data_in<12> ), .C(n4487), .D(\data_in<4> ), 
        .Y(n4483) );
  OAI21X1 U1303 ( .A(n2644), .B(n2962), .C(n4482), .Y(n3488) );
  AOI22X1 U1304 ( .A(n4488), .B(\data_in<13> ), .C(n4487), .D(\data_in<5> ), 
        .Y(n4482) );
  OAI21X1 U1305 ( .A(n2644), .B(n2961), .C(n4481), .Y(n3487) );
  AOI22X1 U1306 ( .A(n4488), .B(\data_in<14> ), .C(n4487), .D(\data_in<6> ), 
        .Y(n4481) );
  OAI21X1 U1307 ( .A(n2644), .B(n2960), .C(n4480), .Y(n3486) );
  AOI22X1 U1308 ( .A(n4488), .B(\data_in<15> ), .C(n4487), .D(\data_in<7> ), 
        .Y(n4480) );
  AOI21X1 U1309 ( .A(n441), .B(n436), .C(n2673), .Y(n4490) );
  OAI21X1 U1310 ( .A(n2643), .B(n2959), .C(n4478), .Y(n3485) );
  AOI22X1 U1311 ( .A(n4477), .B(\data_in<8> ), .C(n4476), .D(\data_in<0> ), 
        .Y(n4478) );
  OAI21X1 U1312 ( .A(n2643), .B(n2958), .C(n4475), .Y(n3484) );
  AOI22X1 U1313 ( .A(n4477), .B(\data_in<9> ), .C(n4476), .D(\data_in<1> ), 
        .Y(n4475) );
  OAI21X1 U1314 ( .A(n2643), .B(n2957), .C(n4474), .Y(n3483) );
  AOI22X1 U1315 ( .A(n4477), .B(\data_in<10> ), .C(n4476), .D(\data_in<2> ), 
        .Y(n4474) );
  OAI21X1 U1316 ( .A(n2643), .B(n2956), .C(n4473), .Y(n3482) );
  AOI22X1 U1317 ( .A(n4477), .B(\data_in<11> ), .C(n4476), .D(\data_in<3> ), 
        .Y(n4473) );
  OAI21X1 U1318 ( .A(n2643), .B(n2955), .C(n4472), .Y(n3481) );
  AOI22X1 U1319 ( .A(n4477), .B(\data_in<12> ), .C(n4476), .D(\data_in<4> ), 
        .Y(n4472) );
  OAI21X1 U1320 ( .A(n2643), .B(n2954), .C(n4471), .Y(n3480) );
  AOI22X1 U1321 ( .A(n4477), .B(\data_in<13> ), .C(n4476), .D(\data_in<5> ), 
        .Y(n4471) );
  OAI21X1 U1322 ( .A(n2643), .B(n2953), .C(n4470), .Y(n3479) );
  AOI22X1 U1323 ( .A(n4477), .B(\data_in<14> ), .C(n4476), .D(\data_in<6> ), 
        .Y(n4470) );
  OAI21X1 U1324 ( .A(n2643), .B(n2952), .C(n4469), .Y(n3478) );
  AOI22X1 U1325 ( .A(n4477), .B(\data_in<15> ), .C(n4476), .D(\data_in<7> ), 
        .Y(n4469) );
  AOI21X1 U1326 ( .A(n436), .B(n438), .C(n2673), .Y(n4479) );
  OAI21X1 U1327 ( .A(n2642), .B(n2951), .C(n4467), .Y(n3477) );
  AOI22X1 U1328 ( .A(n4466), .B(\data_in<8> ), .C(n4465), .D(\data_in<0> ), 
        .Y(n4467) );
  OAI21X1 U1329 ( .A(n2642), .B(n2950), .C(n4464), .Y(n3476) );
  AOI22X1 U1330 ( .A(n4466), .B(\data_in<9> ), .C(n4465), .D(\data_in<1> ), 
        .Y(n4464) );
  OAI21X1 U1331 ( .A(n2642), .B(n2949), .C(n4463), .Y(n3475) );
  AOI22X1 U1332 ( .A(n4466), .B(\data_in<10> ), .C(n4465), .D(\data_in<2> ), 
        .Y(n4463) );
  OAI21X1 U1333 ( .A(n2642), .B(n2948), .C(n4462), .Y(n3474) );
  AOI22X1 U1334 ( .A(n4466), .B(\data_in<11> ), .C(n4465), .D(\data_in<3> ), 
        .Y(n4462) );
  OAI21X1 U1335 ( .A(n2642), .B(n2947), .C(n4461), .Y(n3473) );
  AOI22X1 U1336 ( .A(n4466), .B(\data_in<12> ), .C(n4465), .D(\data_in<4> ), 
        .Y(n4461) );
  OAI21X1 U1337 ( .A(n2642), .B(n2946), .C(n4460), .Y(n3472) );
  AOI22X1 U1338 ( .A(n4466), .B(\data_in<13> ), .C(n4465), .D(\data_in<5> ), 
        .Y(n4460) );
  OAI21X1 U1339 ( .A(n2642), .B(n2945), .C(n4459), .Y(n3471) );
  AOI22X1 U1340 ( .A(n4466), .B(\data_in<14> ), .C(n4465), .D(\data_in<6> ), 
        .Y(n4459) );
  OAI21X1 U1341 ( .A(n2642), .B(n2944), .C(n4458), .Y(n3470) );
  AOI22X1 U1342 ( .A(n4466), .B(\data_in<15> ), .C(n4465), .D(\data_in<7> ), 
        .Y(n4458) );
  AOI21X1 U1343 ( .A(n438), .B(n432), .C(n2673), .Y(n4468) );
  OAI21X1 U1344 ( .A(n2641), .B(n2943), .C(n4456), .Y(n3469) );
  AOI22X1 U1345 ( .A(n4455), .B(\data_in<8> ), .C(n4454), .D(\data_in<0> ), 
        .Y(n4456) );
  OAI21X1 U1346 ( .A(n2641), .B(n2942), .C(n4453), .Y(n3468) );
  AOI22X1 U1347 ( .A(n4455), .B(\data_in<9> ), .C(n4454), .D(\data_in<1> ), 
        .Y(n4453) );
  OAI21X1 U1348 ( .A(n2641), .B(n2941), .C(n4452), .Y(n3467) );
  AOI22X1 U1349 ( .A(n4455), .B(\data_in<10> ), .C(n4454), .D(\data_in<2> ), 
        .Y(n4452) );
  OAI21X1 U1350 ( .A(n2641), .B(n2940), .C(n4451), .Y(n3466) );
  AOI22X1 U1351 ( .A(n4455), .B(\data_in<11> ), .C(n4454), .D(\data_in<3> ), 
        .Y(n4451) );
  OAI21X1 U1352 ( .A(n2641), .B(n2939), .C(n4450), .Y(n3465) );
  AOI22X1 U1353 ( .A(n4455), .B(\data_in<12> ), .C(n4454), .D(\data_in<4> ), 
        .Y(n4450) );
  OAI21X1 U1354 ( .A(n2641), .B(n2938), .C(n4449), .Y(n3464) );
  AOI22X1 U1355 ( .A(n4455), .B(\data_in<13> ), .C(n4454), .D(\data_in<5> ), 
        .Y(n4449) );
  OAI21X1 U1356 ( .A(n2641), .B(n2937), .C(n4448), .Y(n3463) );
  AOI22X1 U1357 ( .A(n4455), .B(\data_in<14> ), .C(n4454), .D(\data_in<6> ), 
        .Y(n4448) );
  OAI21X1 U1358 ( .A(n2641), .B(n2936), .C(n4447), .Y(n3462) );
  AOI22X1 U1359 ( .A(n4455), .B(\data_in<15> ), .C(n4454), .D(\data_in<7> ), 
        .Y(n4447) );
  AOI21X1 U1360 ( .A(n432), .B(n434), .C(n2673), .Y(n4457) );
  OAI21X1 U1361 ( .A(n2640), .B(n2935), .C(n4445), .Y(n3461) );
  AOI22X1 U1362 ( .A(n4444), .B(\data_in<8> ), .C(n4443), .D(\data_in<0> ), 
        .Y(n4445) );
  OAI21X1 U1363 ( .A(n2640), .B(n2934), .C(n4442), .Y(n3460) );
  AOI22X1 U1364 ( .A(n4444), .B(\data_in<9> ), .C(n4443), .D(\data_in<1> ), 
        .Y(n4442) );
  OAI21X1 U1365 ( .A(n2640), .B(n2933), .C(n4441), .Y(n3459) );
  AOI22X1 U1366 ( .A(n4444), .B(\data_in<10> ), .C(n4443), .D(\data_in<2> ), 
        .Y(n4441) );
  OAI21X1 U1367 ( .A(n2640), .B(n2932), .C(n4440), .Y(n3458) );
  AOI22X1 U1368 ( .A(n4444), .B(\data_in<11> ), .C(n4443), .D(\data_in<3> ), 
        .Y(n4440) );
  OAI21X1 U1369 ( .A(n2640), .B(n2931), .C(n4439), .Y(n3457) );
  AOI22X1 U1370 ( .A(n4444), .B(\data_in<12> ), .C(n4443), .D(\data_in<4> ), 
        .Y(n4439) );
  OAI21X1 U1371 ( .A(n2640), .B(n2930), .C(n4438), .Y(n3456) );
  AOI22X1 U1372 ( .A(n4444), .B(\data_in<13> ), .C(n4443), .D(\data_in<5> ), 
        .Y(n4438) );
  OAI21X1 U1373 ( .A(n2640), .B(n2929), .C(n4437), .Y(n3455) );
  AOI22X1 U1374 ( .A(n4444), .B(\data_in<14> ), .C(n4443), .D(\data_in<6> ), 
        .Y(n4437) );
  OAI21X1 U1375 ( .A(n2640), .B(n2928), .C(n4436), .Y(n3454) );
  AOI22X1 U1376 ( .A(n4444), .B(\data_in<15> ), .C(n4443), .D(\data_in<7> ), 
        .Y(n4436) );
  AOI21X1 U1377 ( .A(n434), .B(n370), .C(n2673), .Y(n4446) );
  OAI21X1 U1378 ( .A(n2639), .B(n2927), .C(n4434), .Y(n3453) );
  AOI22X1 U1379 ( .A(n4433), .B(\data_in<8> ), .C(n4432), .D(\data_in<0> ), 
        .Y(n4434) );
  OAI21X1 U1380 ( .A(n2639), .B(n2926), .C(n4431), .Y(n3452) );
  AOI22X1 U1381 ( .A(n4433), .B(\data_in<9> ), .C(n4432), .D(\data_in<1> ), 
        .Y(n4431) );
  OAI21X1 U1382 ( .A(n2639), .B(n2925), .C(n4430), .Y(n3451) );
  AOI22X1 U1383 ( .A(n4433), .B(\data_in<10> ), .C(n4432), .D(\data_in<2> ), 
        .Y(n4430) );
  OAI21X1 U1384 ( .A(n2639), .B(n2924), .C(n4429), .Y(n3450) );
  AOI22X1 U1385 ( .A(n4433), .B(\data_in<11> ), .C(n4432), .D(\data_in<3> ), 
        .Y(n4429) );
  OAI21X1 U1386 ( .A(n2639), .B(n2923), .C(n4428), .Y(n3449) );
  AOI22X1 U1387 ( .A(n4433), .B(\data_in<12> ), .C(n4432), .D(\data_in<4> ), 
        .Y(n4428) );
  OAI21X1 U1388 ( .A(n2639), .B(n2922), .C(n4427), .Y(n3448) );
  AOI22X1 U1389 ( .A(n4433), .B(\data_in<13> ), .C(n4432), .D(\data_in<5> ), 
        .Y(n4427) );
  OAI21X1 U1390 ( .A(n2639), .B(n2921), .C(n4426), .Y(n3447) );
  AOI22X1 U1391 ( .A(n4433), .B(\data_in<14> ), .C(n4432), .D(\data_in<6> ), 
        .Y(n4426) );
  OAI21X1 U1392 ( .A(n2639), .B(n2920), .C(n4425), .Y(n3446) );
  AOI22X1 U1393 ( .A(n4433), .B(\data_in<15> ), .C(n4432), .D(\data_in<7> ), 
        .Y(n4425) );
  AOI21X1 U1394 ( .A(n370), .B(n372), .C(n2673), .Y(n4435) );
  OAI21X1 U1395 ( .A(n2638), .B(n2919), .C(n4423), .Y(n3445) );
  AOI22X1 U1396 ( .A(n4422), .B(\data_in<8> ), .C(n4421), .D(\data_in<0> ), 
        .Y(n4423) );
  OAI21X1 U1397 ( .A(n2638), .B(n2918), .C(n4420), .Y(n3444) );
  AOI22X1 U1398 ( .A(n4422), .B(\data_in<9> ), .C(n4421), .D(\data_in<1> ), 
        .Y(n4420) );
  OAI21X1 U1399 ( .A(n2638), .B(n2917), .C(n4419), .Y(n3443) );
  AOI22X1 U1400 ( .A(n4422), .B(\data_in<10> ), .C(n4421), .D(\data_in<2> ), 
        .Y(n4419) );
  OAI21X1 U1401 ( .A(n2638), .B(n2916), .C(n4418), .Y(n3442) );
  AOI22X1 U1402 ( .A(n4422), .B(\data_in<11> ), .C(n4421), .D(\data_in<3> ), 
        .Y(n4418) );
  OAI21X1 U1403 ( .A(n2638), .B(n2915), .C(n4417), .Y(n3441) );
  AOI22X1 U1404 ( .A(n4422), .B(\data_in<12> ), .C(n4421), .D(\data_in<4> ), 
        .Y(n4417) );
  OAI21X1 U1405 ( .A(n2638), .B(n2914), .C(n4416), .Y(n3440) );
  AOI22X1 U1406 ( .A(n4422), .B(\data_in<13> ), .C(n4421), .D(\data_in<5> ), 
        .Y(n4416) );
  OAI21X1 U1407 ( .A(n2638), .B(n2913), .C(n4415), .Y(n3439) );
  AOI22X1 U1408 ( .A(n4422), .B(\data_in<14> ), .C(n4421), .D(\data_in<6> ), 
        .Y(n4415) );
  OAI21X1 U1409 ( .A(n2638), .B(n2912), .C(n4414), .Y(n3438) );
  AOI22X1 U1410 ( .A(n4422), .B(\data_in<15> ), .C(n4421), .D(\data_in<7> ), 
        .Y(n4414) );
  AOI21X1 U1411 ( .A(n372), .B(n366), .C(n2672), .Y(n4424) );
  OAI21X1 U1412 ( .A(n2637), .B(n2911), .C(n4412), .Y(n3437) );
  AOI22X1 U1413 ( .A(n4411), .B(\data_in<8> ), .C(n4410), .D(\data_in<0> ), 
        .Y(n4412) );
  OAI21X1 U1414 ( .A(n2637), .B(n2910), .C(n4409), .Y(n3436) );
  AOI22X1 U1415 ( .A(n4411), .B(\data_in<9> ), .C(n4410), .D(\data_in<1> ), 
        .Y(n4409) );
  OAI21X1 U1416 ( .A(n2637), .B(n2909), .C(n4408), .Y(n3435) );
  AOI22X1 U1417 ( .A(n4411), .B(\data_in<10> ), .C(n4410), .D(\data_in<2> ), 
        .Y(n4408) );
  OAI21X1 U1418 ( .A(n2637), .B(n2908), .C(n4407), .Y(n3434) );
  AOI22X1 U1419 ( .A(n4411), .B(\data_in<11> ), .C(n4410), .D(\data_in<3> ), 
        .Y(n4407) );
  OAI21X1 U1420 ( .A(n2637), .B(n2907), .C(n4406), .Y(n3433) );
  AOI22X1 U1421 ( .A(n4411), .B(\data_in<12> ), .C(n4410), .D(\data_in<4> ), 
        .Y(n4406) );
  OAI21X1 U1422 ( .A(n2637), .B(n2906), .C(n4405), .Y(n3432) );
  AOI22X1 U1423 ( .A(n4411), .B(\data_in<13> ), .C(n4410), .D(\data_in<5> ), 
        .Y(n4405) );
  OAI21X1 U1424 ( .A(n2637), .B(n2905), .C(n4404), .Y(n3431) );
  AOI22X1 U1425 ( .A(n4411), .B(\data_in<14> ), .C(n4410), .D(\data_in<6> ), 
        .Y(n4404) );
  OAI21X1 U1426 ( .A(n2637), .B(n2904), .C(n4403), .Y(n3430) );
  AOI22X1 U1427 ( .A(n4411), .B(\data_in<15> ), .C(n4410), .D(\data_in<7> ), 
        .Y(n4403) );
  AOI21X1 U1428 ( .A(n366), .B(n368), .C(n2673), .Y(n4413) );
  OAI21X1 U1429 ( .A(n2636), .B(n2903), .C(n4401), .Y(n3429) );
  AOI22X1 U1430 ( .A(n4400), .B(\data_in<8> ), .C(n4399), .D(\data_in<0> ), 
        .Y(n4401) );
  OAI21X1 U1431 ( .A(n2636), .B(n2902), .C(n4398), .Y(n3428) );
  AOI22X1 U1432 ( .A(n4400), .B(\data_in<9> ), .C(n4399), .D(\data_in<1> ), 
        .Y(n4398) );
  OAI21X1 U1433 ( .A(n2636), .B(n2901), .C(n4397), .Y(n3427) );
  AOI22X1 U1434 ( .A(n4400), .B(\data_in<10> ), .C(n4399), .D(\data_in<2> ), 
        .Y(n4397) );
  OAI21X1 U1435 ( .A(n2636), .B(n2900), .C(n4396), .Y(n3426) );
  AOI22X1 U1436 ( .A(n4400), .B(\data_in<11> ), .C(n4399), .D(\data_in<3> ), 
        .Y(n4396) );
  OAI21X1 U1437 ( .A(n2636), .B(n2899), .C(n4395), .Y(n3425) );
  AOI22X1 U1438 ( .A(n4400), .B(\data_in<12> ), .C(n4399), .D(\data_in<4> ), 
        .Y(n4395) );
  OAI21X1 U1439 ( .A(n2636), .B(n2898), .C(n4394), .Y(n3424) );
  AOI22X1 U1440 ( .A(n4400), .B(\data_in<13> ), .C(n4399), .D(\data_in<5> ), 
        .Y(n4394) );
  OAI21X1 U1441 ( .A(n2636), .B(n2897), .C(n4393), .Y(n3423) );
  AOI22X1 U1442 ( .A(n4400), .B(\data_in<14> ), .C(n4399), .D(\data_in<6> ), 
        .Y(n4393) );
  OAI21X1 U1443 ( .A(n2636), .B(n2896), .C(n4392), .Y(n3422) );
  AOI22X1 U1444 ( .A(n4400), .B(\data_in<15> ), .C(n4399), .D(\data_in<7> ), 
        .Y(n4392) );
  AOI21X1 U1445 ( .A(n368), .B(n362), .C(n2673), .Y(n4402) );
  OAI21X1 U1446 ( .A(n2635), .B(n2895), .C(n4390), .Y(n3421) );
  AOI22X1 U1447 ( .A(n4389), .B(\data_in<8> ), .C(n4388), .D(\data_in<0> ), 
        .Y(n4390) );
  OAI21X1 U1448 ( .A(n2635), .B(n2894), .C(n4387), .Y(n3420) );
  AOI22X1 U1449 ( .A(n4389), .B(\data_in<9> ), .C(n4388), .D(\data_in<1> ), 
        .Y(n4387) );
  OAI21X1 U1450 ( .A(n2635), .B(n2893), .C(n4386), .Y(n3419) );
  AOI22X1 U1451 ( .A(n4389), .B(\data_in<10> ), .C(n4388), .D(\data_in<2> ), 
        .Y(n4386) );
  OAI21X1 U1452 ( .A(n2635), .B(n2892), .C(n4385), .Y(n3418) );
  AOI22X1 U1453 ( .A(n4389), .B(\data_in<11> ), .C(n4388), .D(\data_in<3> ), 
        .Y(n4385) );
  OAI21X1 U1454 ( .A(n2635), .B(n2891), .C(n4384), .Y(n3417) );
  AOI22X1 U1455 ( .A(n4389), .B(\data_in<12> ), .C(n4388), .D(\data_in<4> ), 
        .Y(n4384) );
  OAI21X1 U1456 ( .A(n2635), .B(n2890), .C(n4383), .Y(n3416) );
  AOI22X1 U1457 ( .A(n4389), .B(\data_in<13> ), .C(n4388), .D(\data_in<5> ), 
        .Y(n4383) );
  OAI21X1 U1458 ( .A(n2635), .B(n2889), .C(n4382), .Y(n3415) );
  AOI22X1 U1459 ( .A(n4389), .B(\data_in<14> ), .C(n4388), .D(\data_in<6> ), 
        .Y(n4382) );
  OAI21X1 U1460 ( .A(n2635), .B(n2888), .C(n4381), .Y(n3414) );
  AOI22X1 U1461 ( .A(n4389), .B(\data_in<15> ), .C(n4388), .D(\data_in<7> ), 
        .Y(n4381) );
  AOI21X1 U1462 ( .A(n362), .B(n364), .C(n2673), .Y(n4391) );
  OAI21X1 U1463 ( .A(n2634), .B(n2887), .C(n4379), .Y(n3413) );
  AOI22X1 U1464 ( .A(n4378), .B(\data_in<8> ), .C(n4377), .D(\data_in<0> ), 
        .Y(n4379) );
  OAI21X1 U1465 ( .A(n2634), .B(n2886), .C(n4376), .Y(n3412) );
  AOI22X1 U1466 ( .A(n4378), .B(\data_in<9> ), .C(n4377), .D(\data_in<1> ), 
        .Y(n4376) );
  OAI21X1 U1467 ( .A(n2634), .B(n2885), .C(n4375), .Y(n3411) );
  AOI22X1 U1468 ( .A(n4378), .B(\data_in<10> ), .C(n4377), .D(\data_in<2> ), 
        .Y(n4375) );
  OAI21X1 U1469 ( .A(n2634), .B(n2884), .C(n4374), .Y(n3410) );
  AOI22X1 U1470 ( .A(n4378), .B(\data_in<11> ), .C(n4377), .D(\data_in<3> ), 
        .Y(n4374) );
  OAI21X1 U1471 ( .A(n2634), .B(n2883), .C(n4373), .Y(n3409) );
  AOI22X1 U1472 ( .A(n4378), .B(\data_in<12> ), .C(n4377), .D(\data_in<4> ), 
        .Y(n4373) );
  OAI21X1 U1473 ( .A(n2634), .B(n2882), .C(n4372), .Y(n3408) );
  AOI22X1 U1474 ( .A(n4378), .B(\data_in<13> ), .C(n4377), .D(\data_in<5> ), 
        .Y(n4372) );
  OAI21X1 U1475 ( .A(n2634), .B(n2881), .C(n4371), .Y(n3407) );
  AOI22X1 U1476 ( .A(n4378), .B(\data_in<14> ), .C(n4377), .D(\data_in<6> ), 
        .Y(n4371) );
  OAI21X1 U1477 ( .A(n2634), .B(n2880), .C(n4370), .Y(n3406) );
  AOI22X1 U1478 ( .A(n4378), .B(\data_in<15> ), .C(n4377), .D(\data_in<7> ), 
        .Y(n4370) );
  AOI21X1 U1479 ( .A(n364), .B(n358), .C(n2673), .Y(n4380) );
  OAI21X1 U1480 ( .A(n2633), .B(n2879), .C(n4368), .Y(n3405) );
  AOI22X1 U1481 ( .A(n4367), .B(\data_in<8> ), .C(n4366), .D(\data_in<0> ), 
        .Y(n4368) );
  OAI21X1 U1482 ( .A(n2633), .B(n2878), .C(n4365), .Y(n3404) );
  AOI22X1 U1483 ( .A(n4367), .B(\data_in<9> ), .C(n4366), .D(\data_in<1> ), 
        .Y(n4365) );
  OAI21X1 U1484 ( .A(n2633), .B(n2877), .C(n4364), .Y(n3403) );
  AOI22X1 U1485 ( .A(n4367), .B(\data_in<10> ), .C(n4366), .D(\data_in<2> ), 
        .Y(n4364) );
  OAI21X1 U1486 ( .A(n2633), .B(n2876), .C(n4363), .Y(n3402) );
  AOI22X1 U1487 ( .A(n4367), .B(\data_in<11> ), .C(n4366), .D(\data_in<3> ), 
        .Y(n4363) );
  OAI21X1 U1488 ( .A(n2633), .B(n2875), .C(n4362), .Y(n3401) );
  AOI22X1 U1489 ( .A(n4367), .B(\data_in<12> ), .C(n4366), .D(\data_in<4> ), 
        .Y(n4362) );
  OAI21X1 U1490 ( .A(n2633), .B(n2874), .C(n4361), .Y(n3400) );
  AOI22X1 U1491 ( .A(n4367), .B(\data_in<13> ), .C(n4366), .D(\data_in<5> ), 
        .Y(n4361) );
  OAI21X1 U1492 ( .A(n2633), .B(n2873), .C(n4360), .Y(n3399) );
  AOI22X1 U1493 ( .A(n4367), .B(\data_in<14> ), .C(n4366), .D(\data_in<6> ), 
        .Y(n4360) );
  OAI21X1 U1494 ( .A(n2633), .B(n2872), .C(n4359), .Y(n3398) );
  AOI22X1 U1495 ( .A(n4367), .B(\data_in<15> ), .C(n4366), .D(\data_in<7> ), 
        .Y(n4359) );
  AOI21X1 U1496 ( .A(n358), .B(n360), .C(n2673), .Y(n4369) );
  OAI21X1 U1497 ( .A(n2632), .B(n2871), .C(n4357), .Y(n3397) );
  AOI22X1 U1498 ( .A(n4356), .B(\data_in<8> ), .C(n4355), .D(\data_in<0> ), 
        .Y(n4357) );
  OAI21X1 U1499 ( .A(n2632), .B(n2870), .C(n4354), .Y(n3396) );
  AOI22X1 U1500 ( .A(n4356), .B(\data_in<9> ), .C(n4355), .D(\data_in<1> ), 
        .Y(n4354) );
  OAI21X1 U1501 ( .A(n2632), .B(n2869), .C(n4353), .Y(n3395) );
  AOI22X1 U1502 ( .A(n4356), .B(\data_in<10> ), .C(n4355), .D(\data_in<2> ), 
        .Y(n4353) );
  OAI21X1 U1503 ( .A(n2632), .B(n2868), .C(n4352), .Y(n3394) );
  AOI22X1 U1504 ( .A(n4356), .B(\data_in<11> ), .C(n4355), .D(\data_in<3> ), 
        .Y(n4352) );
  OAI21X1 U1505 ( .A(n2632), .B(n2867), .C(n4351), .Y(n3393) );
  AOI22X1 U1506 ( .A(n4356), .B(\data_in<12> ), .C(n4355), .D(\data_in<4> ), 
        .Y(n4351) );
  OAI21X1 U1507 ( .A(n2632), .B(n2866), .C(n4350), .Y(n3392) );
  AOI22X1 U1508 ( .A(n4356), .B(\data_in<13> ), .C(n4355), .D(\data_in<5> ), 
        .Y(n4350) );
  OAI21X1 U1509 ( .A(n2632), .B(n2865), .C(n4349), .Y(n3391) );
  AOI22X1 U1510 ( .A(n4356), .B(\data_in<14> ), .C(n4355), .D(\data_in<6> ), 
        .Y(n4349) );
  OAI21X1 U1511 ( .A(n2632), .B(n2864), .C(n4348), .Y(n3390) );
  AOI22X1 U1512 ( .A(n4356), .B(\data_in<15> ), .C(n4355), .D(\data_in<7> ), 
        .Y(n4348) );
  AOI21X1 U1513 ( .A(n360), .B(n386), .C(n2673), .Y(n4358) );
  OAI21X1 U1514 ( .A(n2631), .B(n2863), .C(n4346), .Y(n3389) );
  AOI22X1 U1515 ( .A(n4345), .B(\data_in<8> ), .C(n4344), .D(\data_in<0> ), 
        .Y(n4346) );
  OAI21X1 U1516 ( .A(n2631), .B(n2862), .C(n4343), .Y(n3388) );
  AOI22X1 U1517 ( .A(n4345), .B(\data_in<9> ), .C(n4344), .D(\data_in<1> ), 
        .Y(n4343) );
  OAI21X1 U1518 ( .A(n2631), .B(n2861), .C(n4342), .Y(n3387) );
  AOI22X1 U1519 ( .A(n4345), .B(\data_in<10> ), .C(n4344), .D(\data_in<2> ), 
        .Y(n4342) );
  OAI21X1 U1520 ( .A(n2631), .B(n2860), .C(n4341), .Y(n3386) );
  AOI22X1 U1521 ( .A(n4345), .B(\data_in<11> ), .C(n4344), .D(\data_in<3> ), 
        .Y(n4341) );
  OAI21X1 U1522 ( .A(n2631), .B(n2859), .C(n4340), .Y(n3385) );
  AOI22X1 U1523 ( .A(n4345), .B(\data_in<12> ), .C(n4344), .D(\data_in<4> ), 
        .Y(n4340) );
  OAI21X1 U1524 ( .A(n2631), .B(n2858), .C(n4339), .Y(n3384) );
  AOI22X1 U1525 ( .A(n4345), .B(\data_in<13> ), .C(n4344), .D(\data_in<5> ), 
        .Y(n4339) );
  OAI21X1 U1526 ( .A(n2631), .B(n2857), .C(n4338), .Y(n3383) );
  AOI22X1 U1527 ( .A(n4345), .B(\data_in<14> ), .C(n4344), .D(\data_in<6> ), 
        .Y(n4338) );
  OAI21X1 U1528 ( .A(n2631), .B(n2856), .C(n4337), .Y(n3382) );
  AOI22X1 U1529 ( .A(n4345), .B(\data_in<15> ), .C(n4344), .D(\data_in<7> ), 
        .Y(n4337) );
  AOI21X1 U1530 ( .A(n386), .B(n387), .C(n2673), .Y(n4347) );
  OAI21X1 U1531 ( .A(n2630), .B(n2855), .C(n4335), .Y(n3381) );
  AOI22X1 U1532 ( .A(n4334), .B(\data_in<8> ), .C(n4333), .D(\data_in<0> ), 
        .Y(n4335) );
  OAI21X1 U1533 ( .A(n2630), .B(n2854), .C(n4332), .Y(n3380) );
  AOI22X1 U1534 ( .A(n4334), .B(\data_in<9> ), .C(n4333), .D(\data_in<1> ), 
        .Y(n4332) );
  OAI21X1 U1535 ( .A(n2630), .B(n2853), .C(n4331), .Y(n3379) );
  AOI22X1 U1536 ( .A(n4334), .B(\data_in<10> ), .C(n4333), .D(\data_in<2> ), 
        .Y(n4331) );
  OAI21X1 U1537 ( .A(n2630), .B(n2852), .C(n4330), .Y(n3378) );
  AOI22X1 U1538 ( .A(n4334), .B(\data_in<11> ), .C(n4333), .D(\data_in<3> ), 
        .Y(n4330) );
  OAI21X1 U1539 ( .A(n2630), .B(n2851), .C(n4329), .Y(n3377) );
  AOI22X1 U1540 ( .A(n4334), .B(\data_in<12> ), .C(n4333), .D(\data_in<4> ), 
        .Y(n4329) );
  OAI21X1 U1541 ( .A(n2630), .B(n2850), .C(n4328), .Y(n3376) );
  AOI22X1 U1542 ( .A(n4334), .B(\data_in<13> ), .C(n4333), .D(\data_in<5> ), 
        .Y(n4328) );
  OAI21X1 U1543 ( .A(n2630), .B(n2849), .C(n4327), .Y(n3375) );
  AOI22X1 U1544 ( .A(n4334), .B(\data_in<14> ), .C(n4333), .D(\data_in<6> ), 
        .Y(n4327) );
  OAI21X1 U1545 ( .A(n2630), .B(n2848), .C(n4326), .Y(n3374) );
  AOI22X1 U1546 ( .A(n4334), .B(\data_in<15> ), .C(n4333), .D(\data_in<7> ), 
        .Y(n4326) );
  AOI21X1 U1547 ( .A(n387), .B(n382), .C(n2673), .Y(n4336) );
  OAI21X1 U1548 ( .A(n2629), .B(n2847), .C(n4324), .Y(n3373) );
  AOI22X1 U1549 ( .A(n4323), .B(\data_in<8> ), .C(n4322), .D(\data_in<0> ), 
        .Y(n4324) );
  OAI21X1 U1550 ( .A(n2629), .B(n2846), .C(n4321), .Y(n3372) );
  AOI22X1 U1551 ( .A(n4323), .B(\data_in<9> ), .C(n4322), .D(\data_in<1> ), 
        .Y(n4321) );
  OAI21X1 U1552 ( .A(n2629), .B(n2845), .C(n4320), .Y(n3371) );
  AOI22X1 U1553 ( .A(n4323), .B(\data_in<10> ), .C(n4322), .D(\data_in<2> ), 
        .Y(n4320) );
  OAI21X1 U1554 ( .A(n2629), .B(n2844), .C(n4319), .Y(n3370) );
  AOI22X1 U1555 ( .A(n4323), .B(\data_in<11> ), .C(n4322), .D(\data_in<3> ), 
        .Y(n4319) );
  OAI21X1 U1556 ( .A(n2629), .B(n2843), .C(n4318), .Y(n3369) );
  AOI22X1 U1557 ( .A(n4323), .B(\data_in<12> ), .C(n4322), .D(\data_in<4> ), 
        .Y(n4318) );
  OAI21X1 U1558 ( .A(n2629), .B(n2842), .C(n4317), .Y(n3368) );
  AOI22X1 U1559 ( .A(n4323), .B(\data_in<13> ), .C(n4322), .D(\data_in<5> ), 
        .Y(n4317) );
  OAI21X1 U1560 ( .A(n2629), .B(n2841), .C(n4316), .Y(n3367) );
  AOI22X1 U1561 ( .A(n4323), .B(\data_in<14> ), .C(n4322), .D(\data_in<6> ), 
        .Y(n4316) );
  OAI21X1 U1562 ( .A(n2629), .B(n2840), .C(n4315), .Y(n3366) );
  AOI22X1 U1563 ( .A(n4323), .B(\data_in<15> ), .C(n4322), .D(\data_in<7> ), 
        .Y(n4315) );
  AOI21X1 U1564 ( .A(n382), .B(n383), .C(n2673), .Y(n4325) );
  OAI21X1 U1565 ( .A(n2628), .B(n2839), .C(n4313), .Y(n3365) );
  AOI22X1 U1566 ( .A(n4312), .B(\data_in<8> ), .C(n4311), .D(\data_in<0> ), 
        .Y(n4313) );
  OAI21X1 U1567 ( .A(n2628), .B(n2838), .C(n4310), .Y(n3364) );
  AOI22X1 U1568 ( .A(n4312), .B(\data_in<9> ), .C(n4311), .D(\data_in<1> ), 
        .Y(n4310) );
  OAI21X1 U1569 ( .A(n2628), .B(n2837), .C(n4309), .Y(n3363) );
  AOI22X1 U1570 ( .A(n4312), .B(\data_in<10> ), .C(n4311), .D(\data_in<2> ), 
        .Y(n4309) );
  OAI21X1 U1571 ( .A(n2628), .B(n2836), .C(n4308), .Y(n3362) );
  AOI22X1 U1572 ( .A(n4312), .B(\data_in<11> ), .C(n4311), .D(\data_in<3> ), 
        .Y(n4308) );
  OAI21X1 U1573 ( .A(n2628), .B(n2835), .C(n4307), .Y(n3361) );
  AOI22X1 U1574 ( .A(n4312), .B(\data_in<12> ), .C(n4311), .D(\data_in<4> ), 
        .Y(n4307) );
  OAI21X1 U1575 ( .A(n2628), .B(n2834), .C(n4306), .Y(n3360) );
  AOI22X1 U1576 ( .A(n4312), .B(\data_in<13> ), .C(n4311), .D(\data_in<5> ), 
        .Y(n4306) );
  OAI21X1 U1577 ( .A(n2628), .B(n2833), .C(n4305), .Y(n3359) );
  AOI22X1 U1578 ( .A(n4312), .B(\data_in<14> ), .C(n4311), .D(\data_in<6> ), 
        .Y(n4305) );
  OAI21X1 U1579 ( .A(n2628), .B(n2832), .C(n4304), .Y(n3358) );
  AOI22X1 U1580 ( .A(n4312), .B(\data_in<15> ), .C(n4311), .D(\data_in<7> ), 
        .Y(n4304) );
  AOI21X1 U1581 ( .A(n383), .B(n378), .C(n2673), .Y(n4314) );
  OAI21X1 U1582 ( .A(n2627), .B(n2831), .C(n4302), .Y(n3357) );
  AOI22X1 U1583 ( .A(n4301), .B(\data_in<8> ), .C(n4300), .D(\data_in<0> ), 
        .Y(n4302) );
  OAI21X1 U1584 ( .A(n2627), .B(n2830), .C(n4299), .Y(n3356) );
  AOI22X1 U1585 ( .A(n4301), .B(\data_in<9> ), .C(n4300), .D(\data_in<1> ), 
        .Y(n4299) );
  OAI21X1 U1586 ( .A(n2627), .B(n2829), .C(n4298), .Y(n3355) );
  AOI22X1 U1587 ( .A(n4301), .B(\data_in<10> ), .C(n4300), .D(\data_in<2> ), 
        .Y(n4298) );
  OAI21X1 U1588 ( .A(n2627), .B(n2828), .C(n4297), .Y(n3354) );
  AOI22X1 U1589 ( .A(n4301), .B(\data_in<11> ), .C(n4300), .D(\data_in<3> ), 
        .Y(n4297) );
  OAI21X1 U1590 ( .A(n2627), .B(n2827), .C(n4296), .Y(n3353) );
  AOI22X1 U1591 ( .A(n4301), .B(\data_in<12> ), .C(n4300), .D(\data_in<4> ), 
        .Y(n4296) );
  OAI21X1 U1592 ( .A(n2627), .B(n2826), .C(n4295), .Y(n3352) );
  AOI22X1 U1593 ( .A(n4301), .B(\data_in<13> ), .C(n4300), .D(\data_in<5> ), 
        .Y(n4295) );
  OAI21X1 U1594 ( .A(n2627), .B(n2825), .C(n4294), .Y(n3351) );
  AOI22X1 U1595 ( .A(n4301), .B(\data_in<14> ), .C(n4300), .D(\data_in<6> ), 
        .Y(n4294) );
  OAI21X1 U1596 ( .A(n2627), .B(n2824), .C(n4293), .Y(n3350) );
  AOI22X1 U1597 ( .A(n4301), .B(\data_in<15> ), .C(n4300), .D(\data_in<7> ), 
        .Y(n4293) );
  AOI21X1 U1598 ( .A(n378), .B(n379), .C(n2673), .Y(n4303) );
  OAI21X1 U1599 ( .A(n2626), .B(n2823), .C(n4291), .Y(n3349) );
  AOI22X1 U1600 ( .A(n4290), .B(\data_in<8> ), .C(n4289), .D(\data_in<0> ), 
        .Y(n4291) );
  OAI21X1 U1601 ( .A(n2626), .B(n2822), .C(n4288), .Y(n3348) );
  AOI22X1 U1602 ( .A(n4290), .B(\data_in<9> ), .C(n4289), .D(\data_in<1> ), 
        .Y(n4288) );
  OAI21X1 U1603 ( .A(n2626), .B(n2821), .C(n4287), .Y(n3347) );
  AOI22X1 U1604 ( .A(n4290), .B(\data_in<10> ), .C(n4289), .D(\data_in<2> ), 
        .Y(n4287) );
  OAI21X1 U1605 ( .A(n2626), .B(n2820), .C(n4286), .Y(n3346) );
  AOI22X1 U1606 ( .A(n4290), .B(\data_in<11> ), .C(n4289), .D(\data_in<3> ), 
        .Y(n4286) );
  OAI21X1 U1607 ( .A(n2626), .B(n2819), .C(n4285), .Y(n3345) );
  AOI22X1 U1608 ( .A(n4290), .B(\data_in<12> ), .C(n4289), .D(\data_in<4> ), 
        .Y(n4285) );
  OAI21X1 U1609 ( .A(n2626), .B(n2818), .C(n4284), .Y(n3344) );
  AOI22X1 U1610 ( .A(n4290), .B(\data_in<13> ), .C(n4289), .D(\data_in<5> ), 
        .Y(n4284) );
  OAI21X1 U1611 ( .A(n2626), .B(n2817), .C(n4283), .Y(n3343) );
  AOI22X1 U1612 ( .A(n4290), .B(\data_in<14> ), .C(n4289), .D(\data_in<6> ), 
        .Y(n4283) );
  OAI21X1 U1613 ( .A(n2626), .B(n2816), .C(n4282), .Y(n3342) );
  AOI22X1 U1614 ( .A(n4290), .B(\data_in<15> ), .C(n4289), .D(\data_in<7> ), 
        .Y(n4282) );
  AOI21X1 U1615 ( .A(n379), .B(n374), .C(n2673), .Y(n4292) );
  OAI21X1 U1616 ( .A(n2625), .B(n2815), .C(n4280), .Y(n3341) );
  AOI22X1 U1617 ( .A(n4279), .B(\data_in<8> ), .C(n4278), .D(\data_in<0> ), 
        .Y(n4280) );
  OAI21X1 U1618 ( .A(n2625), .B(n2814), .C(n4277), .Y(n3340) );
  AOI22X1 U1619 ( .A(n4279), .B(\data_in<9> ), .C(n4278), .D(\data_in<1> ), 
        .Y(n4277) );
  OAI21X1 U1620 ( .A(n2625), .B(n2813), .C(n4276), .Y(n3339) );
  AOI22X1 U1621 ( .A(n4279), .B(\data_in<10> ), .C(n4278), .D(\data_in<2> ), 
        .Y(n4276) );
  OAI21X1 U1622 ( .A(n2625), .B(n2812), .C(n4275), .Y(n3338) );
  AOI22X1 U1623 ( .A(n4279), .B(\data_in<11> ), .C(n4278), .D(\data_in<3> ), 
        .Y(n4275) );
  OAI21X1 U1624 ( .A(n2625), .B(n2811), .C(n4274), .Y(n3337) );
  AOI22X1 U1625 ( .A(n4279), .B(\data_in<12> ), .C(n4278), .D(\data_in<4> ), 
        .Y(n4274) );
  OAI21X1 U1626 ( .A(n2625), .B(n2810), .C(n4273), .Y(n3336) );
  AOI22X1 U1627 ( .A(n4279), .B(\data_in<13> ), .C(n4278), .D(\data_in<5> ), 
        .Y(n4273) );
  OAI21X1 U1628 ( .A(n2625), .B(n2809), .C(n4272), .Y(n3335) );
  AOI22X1 U1629 ( .A(n4279), .B(\data_in<14> ), .C(n4278), .D(\data_in<6> ), 
        .Y(n4272) );
  OAI21X1 U1630 ( .A(n2625), .B(n2808), .C(n4271), .Y(n3334) );
  AOI22X1 U1631 ( .A(n4279), .B(\data_in<15> ), .C(n4278), .D(\data_in<7> ), 
        .Y(n4271) );
  AOI21X1 U1632 ( .A(n374), .B(n375), .C(n2673), .Y(n4281) );
  OAI21X1 U1633 ( .A(n2624), .B(n2807), .C(n4269), .Y(n3333) );
  AOI22X1 U1634 ( .A(n4268), .B(\data_in<8> ), .C(n4267), .D(\data_in<0> ), 
        .Y(n4269) );
  OAI21X1 U1635 ( .A(n2624), .B(n2806), .C(n4266), .Y(n3332) );
  AOI22X1 U1636 ( .A(n4268), .B(\data_in<9> ), .C(n4267), .D(\data_in<1> ), 
        .Y(n4266) );
  OAI21X1 U1637 ( .A(n2624), .B(n2805), .C(n4265), .Y(n3331) );
  AOI22X1 U1638 ( .A(n4268), .B(\data_in<10> ), .C(n4267), .D(\data_in<2> ), 
        .Y(n4265) );
  OAI21X1 U1639 ( .A(n2624), .B(n2804), .C(n4264), .Y(n3330) );
  AOI22X1 U1640 ( .A(n4268), .B(\data_in<11> ), .C(n4267), .D(\data_in<3> ), 
        .Y(n4264) );
  OAI21X1 U1641 ( .A(n2624), .B(n2803), .C(n4263), .Y(n3329) );
  AOI22X1 U1642 ( .A(n4268), .B(\data_in<12> ), .C(n4267), .D(\data_in<4> ), 
        .Y(n4263) );
  OAI21X1 U1643 ( .A(n2624), .B(n2802), .C(n4262), .Y(n3328) );
  AOI22X1 U1644 ( .A(n4268), .B(\data_in<13> ), .C(n4267), .D(\data_in<5> ), 
        .Y(n4262) );
  OAI21X1 U1645 ( .A(n2624), .B(n2801), .C(n4261), .Y(n3327) );
  AOI22X1 U1646 ( .A(n4268), .B(\data_in<14> ), .C(n4267), .D(\data_in<6> ), 
        .Y(n4261) );
  OAI21X1 U1647 ( .A(n2624), .B(n2800), .C(n4260), .Y(n3326) );
  AOI22X1 U1648 ( .A(n4268), .B(\data_in<15> ), .C(n4267), .D(\data_in<7> ), 
        .Y(n4260) );
  AOI21X1 U1649 ( .A(n375), .B(n402), .C(n2673), .Y(n4270) );
  OAI21X1 U1650 ( .A(n2623), .B(n2799), .C(n4258), .Y(n3325) );
  AOI22X1 U1651 ( .A(n4257), .B(\data_in<8> ), .C(n4256), .D(\data_in<0> ), 
        .Y(n4258) );
  OAI21X1 U1652 ( .A(n2623), .B(n2798), .C(n4255), .Y(n3324) );
  AOI22X1 U1653 ( .A(n4257), .B(\data_in<9> ), .C(n4256), .D(\data_in<1> ), 
        .Y(n4255) );
  OAI21X1 U1654 ( .A(n2623), .B(n2797), .C(n4254), .Y(n3323) );
  AOI22X1 U1655 ( .A(n4257), .B(\data_in<10> ), .C(n4256), .D(\data_in<2> ), 
        .Y(n4254) );
  OAI21X1 U1656 ( .A(n2623), .B(n2796), .C(n4253), .Y(n3322) );
  AOI22X1 U1657 ( .A(n4257), .B(\data_in<11> ), .C(n4256), .D(\data_in<3> ), 
        .Y(n4253) );
  OAI21X1 U1658 ( .A(n2623), .B(n2795), .C(n4252), .Y(n3321) );
  AOI22X1 U1659 ( .A(n4257), .B(\data_in<12> ), .C(n4256), .D(\data_in<4> ), 
        .Y(n4252) );
  OAI21X1 U1660 ( .A(n2623), .B(n2794), .C(n4251), .Y(n3320) );
  AOI22X1 U1661 ( .A(n4257), .B(\data_in<13> ), .C(n4256), .D(\data_in<5> ), 
        .Y(n4251) );
  OAI21X1 U1662 ( .A(n2623), .B(n2793), .C(n4250), .Y(n3319) );
  AOI22X1 U1663 ( .A(n4257), .B(\data_in<14> ), .C(n4256), .D(\data_in<6> ), 
        .Y(n4250) );
  OAI21X1 U1664 ( .A(n2623), .B(n2792), .C(n4249), .Y(n3318) );
  AOI22X1 U1665 ( .A(n4257), .B(\data_in<15> ), .C(n4256), .D(\data_in<7> ), 
        .Y(n4249) );
  AOI21X1 U1666 ( .A(n402), .B(n403), .C(n2672), .Y(n4259) );
  OAI21X1 U1667 ( .A(n2622), .B(n2791), .C(n4247), .Y(n3317) );
  AOI22X1 U1668 ( .A(n4246), .B(\data_in<8> ), .C(n4245), .D(\data_in<0> ), 
        .Y(n4247) );
  OAI21X1 U1669 ( .A(n2622), .B(n2790), .C(n4244), .Y(n3316) );
  AOI22X1 U1670 ( .A(n4246), .B(\data_in<9> ), .C(n4245), .D(\data_in<1> ), 
        .Y(n4244) );
  OAI21X1 U1671 ( .A(n2622), .B(n2789), .C(n4243), .Y(n3315) );
  AOI22X1 U1672 ( .A(n4246), .B(\data_in<10> ), .C(n4245), .D(\data_in<2> ), 
        .Y(n4243) );
  OAI21X1 U1673 ( .A(n2622), .B(n2788), .C(n4242), .Y(n3314) );
  AOI22X1 U1674 ( .A(n4246), .B(\data_in<11> ), .C(n4245), .D(\data_in<3> ), 
        .Y(n4242) );
  OAI21X1 U1675 ( .A(n2622), .B(n2787), .C(n4241), .Y(n3313) );
  AOI22X1 U1676 ( .A(n4246), .B(\data_in<12> ), .C(n4245), .D(\data_in<4> ), 
        .Y(n4241) );
  OAI21X1 U1677 ( .A(n2622), .B(n2786), .C(n4240), .Y(n3312) );
  AOI22X1 U1678 ( .A(n4246), .B(\data_in<13> ), .C(n4245), .D(\data_in<5> ), 
        .Y(n4240) );
  OAI21X1 U1679 ( .A(n2622), .B(n2785), .C(n4239), .Y(n3311) );
  AOI22X1 U1680 ( .A(n4246), .B(\data_in<14> ), .C(n4245), .D(\data_in<6> ), 
        .Y(n4239) );
  OAI21X1 U1681 ( .A(n2622), .B(n2784), .C(n4238), .Y(n3310) );
  AOI22X1 U1682 ( .A(n4246), .B(\data_in<15> ), .C(n4245), .D(\data_in<7> ), 
        .Y(n4238) );
  AOI21X1 U1683 ( .A(n403), .B(n398), .C(n2672), .Y(n4248) );
  OAI21X1 U1684 ( .A(n2621), .B(n2783), .C(n4236), .Y(n3309) );
  AOI22X1 U1685 ( .A(n4235), .B(\data_in<8> ), .C(n4234), .D(\data_in<0> ), 
        .Y(n4236) );
  OAI21X1 U1686 ( .A(n2621), .B(n2782), .C(n4233), .Y(n3308) );
  AOI22X1 U1687 ( .A(n4235), .B(\data_in<9> ), .C(n4234), .D(\data_in<1> ), 
        .Y(n4233) );
  OAI21X1 U1688 ( .A(n2621), .B(n2781), .C(n4232), .Y(n3307) );
  AOI22X1 U1689 ( .A(n4235), .B(\data_in<10> ), .C(n4234), .D(\data_in<2> ), 
        .Y(n4232) );
  OAI21X1 U1690 ( .A(n2621), .B(n2780), .C(n4231), .Y(n3306) );
  AOI22X1 U1691 ( .A(n4235), .B(\data_in<11> ), .C(n4234), .D(\data_in<3> ), 
        .Y(n4231) );
  OAI21X1 U1692 ( .A(n2621), .B(n2779), .C(n4230), .Y(n3305) );
  AOI22X1 U1693 ( .A(n4235), .B(\data_in<12> ), .C(n4234), .D(\data_in<4> ), 
        .Y(n4230) );
  OAI21X1 U1694 ( .A(n2621), .B(n2778), .C(n4229), .Y(n3304) );
  AOI22X1 U1695 ( .A(n4235), .B(\data_in<13> ), .C(n4234), .D(\data_in<5> ), 
        .Y(n4229) );
  OAI21X1 U1696 ( .A(n2621), .B(n2777), .C(n4228), .Y(n3303) );
  AOI22X1 U1697 ( .A(n4235), .B(\data_in<14> ), .C(n4234), .D(\data_in<6> ), 
        .Y(n4228) );
  OAI21X1 U1698 ( .A(n2621), .B(n2776), .C(n4227), .Y(n3302) );
  AOI22X1 U1699 ( .A(n4235), .B(\data_in<15> ), .C(n4234), .D(\data_in<7> ), 
        .Y(n4227) );
  AOI21X1 U1700 ( .A(n398), .B(n399), .C(n2672), .Y(n4237) );
  OAI21X1 U1701 ( .A(n2620), .B(n2775), .C(n4225), .Y(n3301) );
  AOI22X1 U1702 ( .A(n4224), .B(\data_in<8> ), .C(n4223), .D(\data_in<0> ), 
        .Y(n4225) );
  OAI21X1 U1703 ( .A(n2620), .B(n2774), .C(n4222), .Y(n3300) );
  AOI22X1 U1704 ( .A(n4224), .B(\data_in<9> ), .C(n4223), .D(\data_in<1> ), 
        .Y(n4222) );
  OAI21X1 U1705 ( .A(n2620), .B(n2773), .C(n4221), .Y(n3299) );
  AOI22X1 U1706 ( .A(n4224), .B(\data_in<10> ), .C(n4223), .D(\data_in<2> ), 
        .Y(n4221) );
  OAI21X1 U1707 ( .A(n2620), .B(n2772), .C(n4220), .Y(n3298) );
  AOI22X1 U1708 ( .A(n4224), .B(\data_in<11> ), .C(n4223), .D(\data_in<3> ), 
        .Y(n4220) );
  OAI21X1 U1709 ( .A(n2620), .B(n2771), .C(n4219), .Y(n3297) );
  AOI22X1 U1710 ( .A(n4224), .B(\data_in<12> ), .C(n4223), .D(\data_in<4> ), 
        .Y(n4219) );
  OAI21X1 U1711 ( .A(n2620), .B(n2770), .C(n4218), .Y(n3296) );
  AOI22X1 U1712 ( .A(n4224), .B(\data_in<13> ), .C(n4223), .D(\data_in<5> ), 
        .Y(n4218) );
  OAI21X1 U1713 ( .A(n2620), .B(n2769), .C(n4217), .Y(n3295) );
  AOI22X1 U1714 ( .A(n4224), .B(\data_in<14> ), .C(n4223), .D(\data_in<6> ), 
        .Y(n4217) );
  OAI21X1 U1715 ( .A(n2620), .B(n2768), .C(n4216), .Y(n3294) );
  AOI22X1 U1716 ( .A(n4224), .B(\data_in<15> ), .C(n4223), .D(\data_in<7> ), 
        .Y(n4216) );
  AOI21X1 U1717 ( .A(n399), .B(n394), .C(n2672), .Y(n4226) );
  OAI21X1 U1718 ( .A(n2619), .B(n2767), .C(n4214), .Y(n3293) );
  AOI22X1 U1719 ( .A(n4213), .B(\data_in<8> ), .C(n4212), .D(\data_in<0> ), 
        .Y(n4214) );
  OAI21X1 U1720 ( .A(n2619), .B(n2766), .C(n4211), .Y(n3292) );
  AOI22X1 U1721 ( .A(n4213), .B(\data_in<9> ), .C(n4212), .D(\data_in<1> ), 
        .Y(n4211) );
  OAI21X1 U1722 ( .A(n2619), .B(n2765), .C(n4210), .Y(n3291) );
  AOI22X1 U1723 ( .A(n4213), .B(\data_in<10> ), .C(n4212), .D(\data_in<2> ), 
        .Y(n4210) );
  OAI21X1 U1724 ( .A(n2619), .B(n2764), .C(n4209), .Y(n3290) );
  AOI22X1 U1725 ( .A(n4213), .B(\data_in<11> ), .C(n4212), .D(\data_in<3> ), 
        .Y(n4209) );
  OAI21X1 U1726 ( .A(n2619), .B(n2763), .C(n4208), .Y(n3289) );
  AOI22X1 U1727 ( .A(n4213), .B(\data_in<12> ), .C(n4212), .D(\data_in<4> ), 
        .Y(n4208) );
  OAI21X1 U1728 ( .A(n2619), .B(n2762), .C(n4207), .Y(n3288) );
  AOI22X1 U1729 ( .A(n4213), .B(\data_in<13> ), .C(n4212), .D(\data_in<5> ), 
        .Y(n4207) );
  OAI21X1 U1730 ( .A(n2619), .B(n2761), .C(n4206), .Y(n3287) );
  AOI22X1 U1731 ( .A(n4213), .B(\data_in<14> ), .C(n4212), .D(\data_in<6> ), 
        .Y(n4206) );
  OAI21X1 U1732 ( .A(n2619), .B(n2760), .C(n4205), .Y(n3286) );
  AOI22X1 U1733 ( .A(n4213), .B(\data_in<15> ), .C(n4212), .D(\data_in<7> ), 
        .Y(n4205) );
  AOI21X1 U1734 ( .A(n394), .B(n395), .C(n2672), .Y(n4215) );
  OAI21X1 U1735 ( .A(n2618), .B(n2759), .C(n4203), .Y(n3285) );
  AOI22X1 U1736 ( .A(n4202), .B(\data_in<8> ), .C(n4201), .D(\data_in<0> ), 
        .Y(n4203) );
  OAI21X1 U1737 ( .A(n2618), .B(n2758), .C(n4200), .Y(n3284) );
  AOI22X1 U1738 ( .A(n4202), .B(\data_in<9> ), .C(n4201), .D(\data_in<1> ), 
        .Y(n4200) );
  OAI21X1 U1739 ( .A(n2618), .B(n2757), .C(n4199), .Y(n3283) );
  AOI22X1 U1740 ( .A(n4202), .B(\data_in<10> ), .C(n4201), .D(\data_in<2> ), 
        .Y(n4199) );
  OAI21X1 U1741 ( .A(n2618), .B(n2756), .C(n4198), .Y(n3282) );
  AOI22X1 U1742 ( .A(n4202), .B(\data_in<11> ), .C(n4201), .D(\data_in<3> ), 
        .Y(n4198) );
  OAI21X1 U1743 ( .A(n2618), .B(n2755), .C(n4197), .Y(n3281) );
  AOI22X1 U1744 ( .A(n4202), .B(\data_in<12> ), .C(n4201), .D(\data_in<4> ), 
        .Y(n4197) );
  OAI21X1 U1745 ( .A(n2618), .B(n2754), .C(n4196), .Y(n3280) );
  AOI22X1 U1746 ( .A(n4202), .B(\data_in<13> ), .C(n4201), .D(\data_in<5> ), 
        .Y(n4196) );
  OAI21X1 U1747 ( .A(n2618), .B(n2753), .C(n4195), .Y(n3279) );
  AOI22X1 U1748 ( .A(n4202), .B(\data_in<14> ), .C(n4201), .D(\data_in<6> ), 
        .Y(n4195) );
  OAI21X1 U1749 ( .A(n2618), .B(n2752), .C(n4194), .Y(n3278) );
  AOI22X1 U1750 ( .A(n4202), .B(\data_in<15> ), .C(n4201), .D(\data_in<7> ), 
        .Y(n4194) );
  AOI21X1 U1751 ( .A(n395), .B(n390), .C(n2672), .Y(n4204) );
  OAI21X1 U1752 ( .A(n2617), .B(n2751), .C(n4192), .Y(n3277) );
  AOI22X1 U1753 ( .A(n4191), .B(\data_in<8> ), .C(n4190), .D(\data_in<0> ), 
        .Y(n4192) );
  OAI21X1 U1754 ( .A(n2617), .B(n2750), .C(n4189), .Y(n3276) );
  AOI22X1 U1755 ( .A(n4191), .B(\data_in<9> ), .C(n4190), .D(\data_in<1> ), 
        .Y(n4189) );
  OAI21X1 U1756 ( .A(n2617), .B(n2749), .C(n4188), .Y(n3275) );
  AOI22X1 U1757 ( .A(n4191), .B(\data_in<10> ), .C(n4190), .D(\data_in<2> ), 
        .Y(n4188) );
  OAI21X1 U1758 ( .A(n2617), .B(n2748), .C(n4187), .Y(n3274) );
  AOI22X1 U1759 ( .A(n4191), .B(\data_in<11> ), .C(n4190), .D(\data_in<3> ), 
        .Y(n4187) );
  OAI21X1 U1760 ( .A(n2617), .B(n2747), .C(n4186), .Y(n3273) );
  AOI22X1 U1761 ( .A(n4191), .B(\data_in<12> ), .C(n4190), .D(\data_in<4> ), 
        .Y(n4186) );
  OAI21X1 U1762 ( .A(n2617), .B(n2746), .C(n4185), .Y(n3272) );
  AOI22X1 U1763 ( .A(n4191), .B(\data_in<13> ), .C(n4190), .D(\data_in<5> ), 
        .Y(n4185) );
  OAI21X1 U1764 ( .A(n2617), .B(n2745), .C(n4184), .Y(n3271) );
  AOI22X1 U1765 ( .A(n4191), .B(\data_in<14> ), .C(n4190), .D(\data_in<6> ), 
        .Y(n4184) );
  OAI21X1 U1766 ( .A(n2617), .B(n2744), .C(n4183), .Y(n3270) );
  AOI22X1 U1767 ( .A(n4191), .B(\data_in<15> ), .C(n4190), .D(\data_in<7> ), 
        .Y(n4183) );
  AOI21X1 U1768 ( .A(n390), .B(n392), .C(n2672), .Y(n4193) );
  OAI21X1 U1769 ( .A(n2616), .B(n2743), .C(n4181), .Y(n3269) );
  AOI22X1 U1770 ( .A(n4180), .B(\data_in<8> ), .C(n4179), .D(\data_in<0> ), 
        .Y(n4181) );
  OAI21X1 U1771 ( .A(n2616), .B(n2742), .C(n4178), .Y(n3268) );
  AOI22X1 U1772 ( .A(n4180), .B(\data_in<9> ), .C(n4179), .D(\data_in<1> ), 
        .Y(n4178) );
  OAI21X1 U1773 ( .A(n2616), .B(n2741), .C(n4177), .Y(n3267) );
  AOI22X1 U1774 ( .A(n4180), .B(\data_in<10> ), .C(n4179), .D(\data_in<2> ), 
        .Y(n4177) );
  OAI21X1 U1775 ( .A(n2616), .B(n2740), .C(n4176), .Y(n3266) );
  AOI22X1 U1776 ( .A(n4180), .B(\data_in<11> ), .C(n4179), .D(\data_in<3> ), 
        .Y(n4176) );
  OAI21X1 U1777 ( .A(n2616), .B(n2739), .C(n4175), .Y(n3265) );
  AOI22X1 U1778 ( .A(n4180), .B(\data_in<12> ), .C(n4179), .D(\data_in<4> ), 
        .Y(n4175) );
  OAI21X1 U1779 ( .A(n2616), .B(n2738), .C(n4174), .Y(n3264) );
  AOI22X1 U1780 ( .A(n4180), .B(\data_in<13> ), .C(n4179), .D(\data_in<5> ), 
        .Y(n4174) );
  OAI21X1 U1781 ( .A(n2616), .B(n2737), .C(n4173), .Y(n3263) );
  AOI22X1 U1782 ( .A(n4180), .B(\data_in<14> ), .C(n4179), .D(\data_in<6> ), 
        .Y(n4173) );
  OAI21X1 U1783 ( .A(n2616), .B(n2736), .C(n4172), .Y(n3262) );
  AOI22X1 U1784 ( .A(n4180), .B(\data_in<15> ), .C(n4179), .D(\data_in<7> ), 
        .Y(n4172) );
  AOI21X1 U1785 ( .A(n392), .B(n412), .C(n2672), .Y(n4182) );
  OAI21X1 U1786 ( .A(n2615), .B(n2735), .C(n4170), .Y(n3261) );
  AOI22X1 U1787 ( .A(n4169), .B(\data_in<8> ), .C(n4168), .D(\data_in<0> ), 
        .Y(n4170) );
  OAI21X1 U1788 ( .A(n2615), .B(n2734), .C(n4167), .Y(n3260) );
  AOI22X1 U1789 ( .A(n4169), .B(\data_in<9> ), .C(n4168), .D(\data_in<1> ), 
        .Y(n4167) );
  OAI21X1 U1790 ( .A(n2615), .B(n2733), .C(n4166), .Y(n3259) );
  AOI22X1 U1791 ( .A(n4169), .B(\data_in<10> ), .C(n4168), .D(\data_in<2> ), 
        .Y(n4166) );
  OAI21X1 U1792 ( .A(n2615), .B(n2732), .C(n4165), .Y(n3258) );
  AOI22X1 U1793 ( .A(n4169), .B(\data_in<11> ), .C(n4168), .D(\data_in<3> ), 
        .Y(n4165) );
  OAI21X1 U1794 ( .A(n2615), .B(n2731), .C(n4164), .Y(n3257) );
  AOI22X1 U1795 ( .A(n4169), .B(\data_in<12> ), .C(n4168), .D(\data_in<4> ), 
        .Y(n4164) );
  OAI21X1 U1796 ( .A(n2615), .B(n2730), .C(n4163), .Y(n3256) );
  AOI22X1 U1797 ( .A(n4169), .B(\data_in<13> ), .C(n4168), .D(\data_in<5> ), 
        .Y(n4163) );
  OAI21X1 U1798 ( .A(n2615), .B(n2729), .C(n4162), .Y(n3255) );
  AOI22X1 U1799 ( .A(n4169), .B(\data_in<14> ), .C(n4168), .D(\data_in<6> ), 
        .Y(n4162) );
  OAI21X1 U1800 ( .A(n2615), .B(n2728), .C(n4161), .Y(n3254) );
  AOI22X1 U1801 ( .A(n4169), .B(\data_in<15> ), .C(n4168), .D(\data_in<7> ), 
        .Y(n4161) );
  AOI21X1 U1802 ( .A(n412), .B(n414), .C(n2672), .Y(n4171) );
  OAI21X1 U1803 ( .A(n2614), .B(n2727), .C(n4159), .Y(n3253) );
  AOI22X1 U1804 ( .A(n4158), .B(\data_in<8> ), .C(n4157), .D(\data_in<0> ), 
        .Y(n4159) );
  OAI21X1 U1805 ( .A(n2614), .B(n2726), .C(n4156), .Y(n3252) );
  AOI22X1 U1806 ( .A(n4158), .B(\data_in<9> ), .C(n4157), .D(\data_in<1> ), 
        .Y(n4156) );
  OAI21X1 U1807 ( .A(n2614), .B(n2725), .C(n4155), .Y(n3251) );
  AOI22X1 U1808 ( .A(n4158), .B(\data_in<10> ), .C(n4157), .D(\data_in<2> ), 
        .Y(n4155) );
  OAI21X1 U1809 ( .A(n2614), .B(n2724), .C(n4154), .Y(n3250) );
  AOI22X1 U1810 ( .A(n4158), .B(\data_in<11> ), .C(n4157), .D(\data_in<3> ), 
        .Y(n4154) );
  OAI21X1 U1811 ( .A(n2614), .B(n2723), .C(n4153), .Y(n3249) );
  AOI22X1 U1812 ( .A(n4158), .B(\data_in<12> ), .C(n4157), .D(\data_in<4> ), 
        .Y(n4153) );
  OAI21X1 U1813 ( .A(n2614), .B(n2722), .C(n4152), .Y(n3248) );
  AOI22X1 U1814 ( .A(n4158), .B(\data_in<13> ), .C(n4157), .D(\data_in<5> ), 
        .Y(n4152) );
  OAI21X1 U1815 ( .A(n2614), .B(n2721), .C(n4151), .Y(n3247) );
  AOI22X1 U1816 ( .A(n4158), .B(\data_in<14> ), .C(n4157), .D(\data_in<6> ), 
        .Y(n4151) );
  OAI21X1 U1817 ( .A(n2614), .B(n2720), .C(n4150), .Y(n3246) );
  AOI22X1 U1818 ( .A(n4158), .B(\data_in<15> ), .C(n4157), .D(\data_in<7> ), 
        .Y(n4150) );
  AOI21X1 U1819 ( .A(n414), .B(n408), .C(n2672), .Y(n4160) );
  OAI21X1 U1820 ( .A(n2613), .B(n2719), .C(n4148), .Y(n3245) );
  AOI22X1 U1821 ( .A(n4147), .B(\data_in<8> ), .C(n4146), .D(\data_in<0> ), 
        .Y(n4148) );
  OAI21X1 U1822 ( .A(n2613), .B(n2718), .C(n4145), .Y(n3244) );
  AOI22X1 U1823 ( .A(n4147), .B(\data_in<9> ), .C(n4146), .D(\data_in<1> ), 
        .Y(n4145) );
  OAI21X1 U1824 ( .A(n2613), .B(n2717), .C(n4144), .Y(n3243) );
  AOI22X1 U1825 ( .A(n4147), .B(\data_in<10> ), .C(n4146), .D(\data_in<2> ), 
        .Y(n4144) );
  OAI21X1 U1826 ( .A(n2613), .B(n2716), .C(n4143), .Y(n3242) );
  AOI22X1 U1827 ( .A(n4147), .B(\data_in<11> ), .C(n4146), .D(\data_in<3> ), 
        .Y(n4143) );
  OAI21X1 U1828 ( .A(n2613), .B(n2715), .C(n4142), .Y(n3241) );
  AOI22X1 U1829 ( .A(n4147), .B(\data_in<12> ), .C(n4146), .D(\data_in<4> ), 
        .Y(n4142) );
  OAI21X1 U1830 ( .A(n2613), .B(n2714), .C(n4141), .Y(n3240) );
  AOI22X1 U1831 ( .A(n4147), .B(\data_in<13> ), .C(n4146), .D(\data_in<5> ), 
        .Y(n4141) );
  OAI21X1 U1832 ( .A(n2613), .B(n2713), .C(n4140), .Y(n3239) );
  AOI22X1 U1833 ( .A(n4147), .B(\data_in<14> ), .C(n4146), .D(\data_in<6> ), 
        .Y(n4140) );
  OAI21X1 U1834 ( .A(n2613), .B(n2712), .C(n4139), .Y(n3238) );
  AOI22X1 U1835 ( .A(n4147), .B(\data_in<15> ), .C(n4146), .D(\data_in<7> ), 
        .Y(n4139) );
  AOI21X1 U1836 ( .A(n408), .B(n410), .C(n2672), .Y(n4149) );
  OAI21X1 U1837 ( .A(n2612), .B(n2711), .C(n4137), .Y(n3237) );
  AOI22X1 U1838 ( .A(n4136), .B(\data_in<8> ), .C(n4135), .D(\data_in<0> ), 
        .Y(n4137) );
  OAI21X1 U1839 ( .A(n2612), .B(n2710), .C(n4134), .Y(n3236) );
  AOI22X1 U1840 ( .A(n4136), .B(\data_in<9> ), .C(n4135), .D(\data_in<1> ), 
        .Y(n4134) );
  OAI21X1 U1841 ( .A(n2612), .B(n2709), .C(n4133), .Y(n3235) );
  AOI22X1 U1842 ( .A(n4136), .B(\data_in<10> ), .C(n4135), .D(\data_in<2> ), 
        .Y(n4133) );
  OAI21X1 U1843 ( .A(n2612), .B(n2708), .C(n4132), .Y(n3234) );
  AOI22X1 U1844 ( .A(n4136), .B(\data_in<11> ), .C(n4135), .D(\data_in<3> ), 
        .Y(n4132) );
  OAI21X1 U1845 ( .A(n2612), .B(n2707), .C(n4131), .Y(n3233) );
  AOI22X1 U1846 ( .A(n4136), .B(\data_in<12> ), .C(n4135), .D(\data_in<4> ), 
        .Y(n4131) );
  OAI21X1 U1847 ( .A(n2612), .B(n2706), .C(n4130), .Y(n3232) );
  AOI22X1 U1848 ( .A(n4136), .B(\data_in<13> ), .C(n4135), .D(\data_in<5> ), 
        .Y(n4130) );
  OAI21X1 U1849 ( .A(n2612), .B(n2705), .C(n4129), .Y(n3231) );
  AOI22X1 U1850 ( .A(n4136), .B(\data_in<14> ), .C(n4135), .D(\data_in<6> ), 
        .Y(n4129) );
  OAI21X1 U1851 ( .A(n2612), .B(n2704), .C(n4128), .Y(n3230) );
  AOI22X1 U1852 ( .A(n4136), .B(\data_in<15> ), .C(n4135), .D(\data_in<7> ), 
        .Y(n4128) );
  AOI21X1 U1853 ( .A(n410), .B(n406), .C(n2672), .Y(n4138) );
  OAI21X1 U1854 ( .A(n2611), .B(n2703), .C(n4126), .Y(n3229) );
  AOI22X1 U1855 ( .A(n4125), .B(\data_in<8> ), .C(n4124), .D(\data_in<0> ), 
        .Y(n4126) );
  OAI21X1 U1856 ( .A(n2611), .B(n2702), .C(n4123), .Y(n3228) );
  AOI22X1 U1857 ( .A(n4125), .B(\data_in<9> ), .C(n4124), .D(\data_in<1> ), 
        .Y(n4123) );
  OAI21X1 U1858 ( .A(n2611), .B(n2701), .C(n4122), .Y(n3227) );
  AOI22X1 U1859 ( .A(n4125), .B(\data_in<10> ), .C(n4124), .D(\data_in<2> ), 
        .Y(n4122) );
  OAI21X1 U1860 ( .A(n2611), .B(n2700), .C(n4121), .Y(n3226) );
  AOI22X1 U1861 ( .A(n4125), .B(\data_in<11> ), .C(n4124), .D(\data_in<3> ), 
        .Y(n4121) );
  OAI21X1 U1862 ( .A(n2611), .B(n2699), .C(n4120), .Y(n3225) );
  AOI22X1 U1863 ( .A(n4125), .B(\data_in<12> ), .C(n4124), .D(\data_in<4> ), 
        .Y(n4120) );
  OAI21X1 U1864 ( .A(n2611), .B(n2698), .C(n4119), .Y(n3224) );
  AOI22X1 U1865 ( .A(n4125), .B(\data_in<13> ), .C(n4124), .D(\data_in<5> ), 
        .Y(n4119) );
  OAI21X1 U1866 ( .A(n2611), .B(n2697), .C(n4118), .Y(n3223) );
  AOI22X1 U1867 ( .A(n4125), .B(\data_in<14> ), .C(n4124), .D(\data_in<6> ), 
        .Y(n4118) );
  OAI21X1 U1868 ( .A(n2611), .B(n2696), .C(n4117), .Y(n3222) );
  AOI22X1 U1869 ( .A(n4125), .B(\data_in<15> ), .C(n4124), .D(\data_in<7> ), 
        .Y(n4117) );
  AOI21X1 U1870 ( .A(n406), .B(n478), .C(n2672), .Y(n4127) );
  OAI21X1 U1871 ( .A(n2610), .B(n2695), .C(n4115), .Y(n3221) );
  AOI22X1 U1872 ( .A(n4114), .B(\data_in<8> ), .C(n4113), .D(\data_in<0> ), 
        .Y(n4115) );
  OAI21X1 U1873 ( .A(n2610), .B(n2694), .C(n4112), .Y(n3220) );
  AOI22X1 U1874 ( .A(n4114), .B(\data_in<9> ), .C(n4113), .D(\data_in<1> ), 
        .Y(n4112) );
  OAI21X1 U1875 ( .A(n2610), .B(n2693), .C(n4111), .Y(n3219) );
  AOI22X1 U1876 ( .A(n4114), .B(\data_in<10> ), .C(n4113), .D(\data_in<2> ), 
        .Y(n4111) );
  OAI21X1 U1877 ( .A(n2610), .B(n2692), .C(n4110), .Y(n3218) );
  AOI22X1 U1878 ( .A(n4114), .B(\data_in<11> ), .C(n4113), .D(\data_in<3> ), 
        .Y(n4110) );
  OAI21X1 U1879 ( .A(n2610), .B(n2691), .C(n4109), .Y(n3217) );
  AOI22X1 U1880 ( .A(n4114), .B(\data_in<12> ), .C(n4113), .D(\data_in<4> ), 
        .Y(n4109) );
  OAI21X1 U1881 ( .A(n2610), .B(n2690), .C(n4108), .Y(n3216) );
  AOI22X1 U1882 ( .A(n4114), .B(\data_in<13> ), .C(n4113), .D(\data_in<5> ), 
        .Y(n4108) );
  OAI21X1 U1883 ( .A(n2610), .B(n2689), .C(n4107), .Y(n3215) );
  AOI22X1 U1884 ( .A(n4114), .B(\data_in<14> ), .C(n4113), .D(\data_in<6> ), 
        .Y(n4107) );
  OAI21X1 U1885 ( .A(n2610), .B(n2688), .C(n4106), .Y(n3214) );
  AOI22X1 U1886 ( .A(n4114), .B(\data_in<15> ), .C(n4113), .D(\data_in<7> ), 
        .Y(n4106) );
  OAI21X1 U1887 ( .A(n2672), .B(n478), .C(n354), .Y(n4116) );
  OAI21X1 U1888 ( .A(n353), .B(n2687), .C(n4105), .Y(n3213) );
  NAND2X1 U1889 ( .A(n353), .B(\data_in<8> ), .Y(n4105) );
  OAI21X1 U1890 ( .A(n353), .B(n2686), .C(n4104), .Y(n3212) );
  NAND2X1 U1891 ( .A(n353), .B(\data_in<9> ), .Y(n4104) );
  OAI21X1 U1892 ( .A(n353), .B(n2685), .C(n4103), .Y(n3211) );
  NAND2X1 U1893 ( .A(n353), .B(\data_in<10> ), .Y(n4103) );
  OAI21X1 U1894 ( .A(n353), .B(n2684), .C(n4102), .Y(n3210) );
  NAND2X1 U1895 ( .A(n353), .B(\data_in<11> ), .Y(n4102) );
  OAI21X1 U1896 ( .A(n353), .B(n2683), .C(n4101), .Y(n3209) );
  NAND2X1 U1897 ( .A(n353), .B(\data_in<12> ), .Y(n4101) );
  OAI21X1 U1898 ( .A(n353), .B(n2682), .C(n4100), .Y(n3208) );
  NAND2X1 U1899 ( .A(n353), .B(\data_in<13> ), .Y(n4100) );
  OAI21X1 U1900 ( .A(n353), .B(n2681), .C(n4099), .Y(n3207) );
  NAND2X1 U1901 ( .A(n353), .B(\data_in<14> ), .Y(n4099) );
  OAI21X1 U1902 ( .A(n353), .B(n2680), .C(n4098), .Y(n3206) );
  NAND2X1 U1903 ( .A(n353), .B(\data_in<15> ), .Y(n4098) );
  NAND3X1 U1905 ( .A(enable), .B(n2679), .C(wr), .Y(n4777) );
  AOI21X1 U1906 ( .A(n4097), .B(n4096), .C(n2609), .Y(n4802) );
  NOR3X1 U1907 ( .A(n4094), .B(n201), .C(n258), .Y(n4096) );
  AOI22X1 U1909 ( .A(\mem<55><7> ), .B(n473), .C(\mem<54><7> ), .D(n475), .Y(
        n4089) );
  AOI22X1 U1910 ( .A(\mem<53><7> ), .B(n469), .C(\mem<52><7> ), .D(n471), .Y(
        n4090) );
  AOI22X1 U1911 ( .A(\mem<51><7> ), .B(n465), .C(\mem<50><7> ), .D(n467), .Y(
        n4092) );
  AOI22X1 U1912 ( .A(\mem<49><7> ), .B(n461), .C(\mem<48><7> ), .D(n463), .Y(
        n4093) );
  AOI22X1 U1914 ( .A(\mem<63><7> ), .B(n356), .C(\mem<62><7> ), .D(n459), .Y(
        n4084) );
  AOI22X1 U1915 ( .A(\mem<61><7> ), .B(n456), .C(\mem<60><7> ), .D(n457), .Y(
        n4085) );
  AOI22X1 U1916 ( .A(\mem<59><7> ), .B(n452), .C(\mem<58><7> ), .D(n453), .Y(
        n4087) );
  AOI22X1 U1917 ( .A(\mem<57><7> ), .B(n448), .C(\mem<56><7> ), .D(n449), .Y(
        n4088) );
  AOI22X1 U1919 ( .A(\mem<39><7> ), .B(n443), .C(\mem<38><7> ), .D(n446), .Y(
        n4079) );
  AOI22X1 U1920 ( .A(\mem<37><7> ), .B(n439), .C(\mem<36><7> ), .D(n442), .Y(
        n4080) );
  AOI22X1 U1921 ( .A(\mem<35><7> ), .B(n435), .C(\mem<34><7> ), .D(n437), .Y(
        n4082) );
  AOI22X1 U1922 ( .A(\mem<33><7> ), .B(n431), .C(\mem<32><7> ), .D(n433), .Y(
        n4083) );
  AOI22X1 U1924 ( .A(\mem<47><7> ), .B(n427), .C(\mem<46><7> ), .D(n429), .Y(
        n4074) );
  AOI22X1 U1925 ( .A(\mem<45><7> ), .B(n423), .C(\mem<44><7> ), .D(n425), .Y(
        n4075) );
  AOI22X1 U1926 ( .A(\mem<43><7> ), .B(n419), .C(\mem<42><7> ), .D(n421), .Y(
        n4077) );
  AOI22X1 U1927 ( .A(\mem<41><7> ), .B(n415), .C(\mem<40><7> ), .D(n417), .Y(
        n4078) );
  NOR3X1 U1928 ( .A(n4073), .B(n226), .C(n256), .Y(n4097) );
  AOI22X1 U1930 ( .A(\mem<7><7> ), .B(n3192), .C(\mem<6><7> ), .D(n413), .Y(
        n4068) );
  AOI22X1 U1931 ( .A(\mem<5><7> ), .B(n3193), .C(\mem<4><7> ), .D(n409), .Y(
        n4069) );
  AOI22X1 U1932 ( .A(\mem<3><7> ), .B(n3194), .C(\mem<2><7> ), .D(n477), .Y(
        n4071) );
  AOI22X1 U1933 ( .A(\mem<1><7> ), .B(n351), .C(n4067), .D(\mem<0><7> ), .Y(
        n4072) );
  AOI22X1 U1935 ( .A(\mem<15><7> ), .B(n401), .C(\mem<14><7> ), .D(n404), .Y(
        n4062) );
  AOI22X1 U1936 ( .A(\mem<13><7> ), .B(n397), .C(\mem<12><7> ), .D(n400), .Y(
        n4063) );
  AOI22X1 U1937 ( .A(\mem<11><7> ), .B(n393), .C(\mem<10><7> ), .D(n396), .Y(
        n4065) );
  AOI22X1 U1938 ( .A(\mem<9><7> ), .B(n389), .C(\mem<8><7> ), .D(n391), .Y(
        n4066) );
  AOI22X1 U1940 ( .A(\mem<23><7> ), .B(n385), .C(\mem<22><7> ), .D(n388), .Y(
        n4057) );
  AOI22X1 U1941 ( .A(\mem<21><7> ), .B(n381), .C(\mem<20><7> ), .D(n384), .Y(
        n4058) );
  AOI22X1 U1942 ( .A(\mem<19><7> ), .B(n377), .C(\mem<18><7> ), .D(n380), .Y(
        n4060) );
  AOI22X1 U1943 ( .A(\mem<17><7> ), .B(n373), .C(\mem<16><7> ), .D(n376), .Y(
        n4061) );
  AOI22X1 U1945 ( .A(\mem<31><7> ), .B(n369), .C(\mem<30><7> ), .D(n371), .Y(
        n4052) );
  AOI22X1 U1946 ( .A(\mem<29><7> ), .B(n365), .C(\mem<28><7> ), .D(n367), .Y(
        n4053) );
  AOI22X1 U1947 ( .A(\mem<27><7> ), .B(n361), .C(\mem<26><7> ), .D(n363), .Y(
        n4055) );
  AOI22X1 U1948 ( .A(\mem<25><7> ), .B(n357), .C(\mem<24><7> ), .D(n359), .Y(
        n4056) );
  AOI21X1 U1949 ( .A(n4051), .B(n4050), .C(n2609), .Y(n4803) );
  NOR3X1 U1950 ( .A(n4049), .B(n176), .C(n254), .Y(n4050) );
  AOI22X1 U1952 ( .A(\mem<55><6> ), .B(n473), .C(\mem<54><6> ), .D(n475), .Y(
        n4044) );
  AOI22X1 U1953 ( .A(\mem<53><6> ), .B(n469), .C(\mem<52><6> ), .D(n471), .Y(
        n4045) );
  AOI22X1 U1954 ( .A(\mem<51><6> ), .B(n465), .C(\mem<50><6> ), .D(n467), .Y(
        n4047) );
  AOI22X1 U1955 ( .A(\mem<49><6> ), .B(n461), .C(\mem<48><6> ), .D(n463), .Y(
        n4048) );
  AOI22X1 U1957 ( .A(\mem<63><6> ), .B(n356), .C(\mem<62><6> ), .D(n459), .Y(
        n4039) );
  AOI22X1 U1958 ( .A(\mem<61><6> ), .B(n456), .C(\mem<60><6> ), .D(n457), .Y(
        n4040) );
  AOI22X1 U1959 ( .A(\mem<59><6> ), .B(n452), .C(\mem<58><6> ), .D(n453), .Y(
        n4042) );
  AOI22X1 U1960 ( .A(\mem<57><6> ), .B(n448), .C(\mem<56><6> ), .D(n449), .Y(
        n4043) );
  AOI22X1 U1962 ( .A(\mem<39><6> ), .B(n443), .C(\mem<38><6> ), .D(n446), .Y(
        n4034) );
  AOI22X1 U1963 ( .A(\mem<37><6> ), .B(n439), .C(\mem<36><6> ), .D(n442), .Y(
        n4035) );
  AOI22X1 U1964 ( .A(\mem<35><6> ), .B(n435), .C(\mem<34><6> ), .D(n437), .Y(
        n4037) );
  AOI22X1 U1965 ( .A(\mem<33><6> ), .B(n431), .C(\mem<32><6> ), .D(n433), .Y(
        n4038) );
  AOI22X1 U1967 ( .A(\mem<47><6> ), .B(n427), .C(\mem<46><6> ), .D(n429), .Y(
        n4029) );
  AOI22X1 U1968 ( .A(\mem<45><6> ), .B(n423), .C(\mem<44><6> ), .D(n425), .Y(
        n4030) );
  AOI22X1 U1969 ( .A(\mem<43><6> ), .B(n419), .C(\mem<42><6> ), .D(n421), .Y(
        n4032) );
  AOI22X1 U1970 ( .A(\mem<41><6> ), .B(n415), .C(\mem<40><6> ), .D(n417), .Y(
        n4033) );
  NOR3X1 U1971 ( .A(n4028), .B(n224), .C(n252), .Y(n4051) );
  AOI22X1 U1973 ( .A(\mem<7><6> ), .B(n3192), .C(\mem<6><6> ), .D(n413), .Y(
        n4023) );
  AOI22X1 U1974 ( .A(\mem<5><6> ), .B(n3193), .C(\mem<4><6> ), .D(n409), .Y(
        n4024) );
  AOI22X1 U1975 ( .A(\mem<3><6> ), .B(n3194), .C(\mem<2><6> ), .D(n477), .Y(
        n4026) );
  AOI22X1 U1976 ( .A(\mem<1><6> ), .B(n351), .C(n4067), .D(\mem<0><6> ), .Y(
        n4027) );
  AOI22X1 U1978 ( .A(\mem<15><6> ), .B(n401), .C(\mem<14><6> ), .D(n404), .Y(
        n4018) );
  AOI22X1 U1979 ( .A(\mem<13><6> ), .B(n397), .C(\mem<12><6> ), .D(n400), .Y(
        n4019) );
  AOI22X1 U1980 ( .A(\mem<11><6> ), .B(n393), .C(\mem<10><6> ), .D(n396), .Y(
        n4021) );
  AOI22X1 U1981 ( .A(\mem<9><6> ), .B(n389), .C(\mem<8><6> ), .D(n391), .Y(
        n4022) );
  AOI22X1 U1983 ( .A(\mem<23><6> ), .B(n385), .C(\mem<22><6> ), .D(n388), .Y(
        n4013) );
  AOI22X1 U1984 ( .A(\mem<21><6> ), .B(n381), .C(\mem<20><6> ), .D(n384), .Y(
        n4014) );
  AOI22X1 U1985 ( .A(\mem<19><6> ), .B(n377), .C(\mem<18><6> ), .D(n380), .Y(
        n4016) );
  AOI22X1 U1986 ( .A(\mem<17><6> ), .B(n373), .C(\mem<16><6> ), .D(n376), .Y(
        n4017) );
  AOI22X1 U1988 ( .A(\mem<31><6> ), .B(n369), .C(\mem<30><6> ), .D(n371), .Y(
        n4008) );
  AOI22X1 U1989 ( .A(\mem<29><6> ), .B(n365), .C(\mem<28><6> ), .D(n367), .Y(
        n4009) );
  AOI22X1 U1990 ( .A(\mem<27><6> ), .B(n361), .C(\mem<26><6> ), .D(n363), .Y(
        n4011) );
  AOI22X1 U1991 ( .A(\mem<25><6> ), .B(n357), .C(\mem<24><6> ), .D(n359), .Y(
        n4012) );
  AOI21X1 U1992 ( .A(n4007), .B(n4006), .C(n2609), .Y(n4804) );
  NOR3X1 U1993 ( .A(n4005), .B(n151), .C(n250), .Y(n4006) );
  AOI22X1 U1995 ( .A(\mem<55><5> ), .B(n473), .C(\mem<54><5> ), .D(n475), .Y(
        n4000) );
  AOI22X1 U1996 ( .A(\mem<53><5> ), .B(n469), .C(\mem<52><5> ), .D(n471), .Y(
        n4001) );
  AOI22X1 U1997 ( .A(\mem<51><5> ), .B(n465), .C(\mem<50><5> ), .D(n467), .Y(
        n4003) );
  AOI22X1 U1998 ( .A(\mem<49><5> ), .B(n461), .C(\mem<48><5> ), .D(n463), .Y(
        n4004) );
  AOI22X1 U2000 ( .A(\mem<63><5> ), .B(n356), .C(\mem<62><5> ), .D(n459), .Y(
        n3995) );
  AOI22X1 U2001 ( .A(\mem<61><5> ), .B(n456), .C(\mem<60><5> ), .D(n457), .Y(
        n3996) );
  AOI22X1 U2002 ( .A(\mem<59><5> ), .B(n452), .C(\mem<58><5> ), .D(n453), .Y(
        n3998) );
  AOI22X1 U2003 ( .A(\mem<57><5> ), .B(n448), .C(\mem<56><5> ), .D(n449), .Y(
        n3999) );
  AOI22X1 U2005 ( .A(\mem<39><5> ), .B(n443), .C(\mem<38><5> ), .D(n446), .Y(
        n3990) );
  AOI22X1 U2006 ( .A(\mem<37><5> ), .B(n439), .C(\mem<36><5> ), .D(n442), .Y(
        n3991) );
  AOI22X1 U2007 ( .A(\mem<35><5> ), .B(n435), .C(\mem<34><5> ), .D(n437), .Y(
        n3993) );
  AOI22X1 U2008 ( .A(\mem<33><5> ), .B(n431), .C(\mem<32><5> ), .D(n433), .Y(
        n3994) );
  AOI22X1 U2010 ( .A(\mem<47><5> ), .B(n427), .C(\mem<46><5> ), .D(n429), .Y(
        n3985) );
  AOI22X1 U2011 ( .A(\mem<45><5> ), .B(n423), .C(\mem<44><5> ), .D(n425), .Y(
        n3986) );
  AOI22X1 U2012 ( .A(\mem<43><5> ), .B(n419), .C(\mem<42><5> ), .D(n421), .Y(
        n3988) );
  AOI22X1 U2013 ( .A(\mem<41><5> ), .B(n415), .C(\mem<40><5> ), .D(n417), .Y(
        n3989) );
  NOR3X1 U2014 ( .A(n3984), .B(n222), .C(n248), .Y(n4007) );
  AOI22X1 U2016 ( .A(\mem<7><5> ), .B(n3192), .C(\mem<6><5> ), .D(n413), .Y(
        n3979) );
  AOI22X1 U2017 ( .A(\mem<5><5> ), .B(n3193), .C(\mem<4><5> ), .D(n409), .Y(
        n3980) );
  AOI22X1 U2018 ( .A(\mem<3><5> ), .B(n3194), .C(\mem<2><5> ), .D(n477), .Y(
        n3982) );
  AOI22X1 U2019 ( .A(\mem<1><5> ), .B(n351), .C(n4067), .D(\mem<0><5> ), .Y(
        n3983) );
  AOI22X1 U2021 ( .A(\mem<15><5> ), .B(n401), .C(\mem<14><5> ), .D(n404), .Y(
        n3974) );
  AOI22X1 U2022 ( .A(\mem<13><5> ), .B(n397), .C(\mem<12><5> ), .D(n400), .Y(
        n3975) );
  AOI22X1 U2023 ( .A(\mem<11><5> ), .B(n393), .C(\mem<10><5> ), .D(n396), .Y(
        n3977) );
  AOI22X1 U2024 ( .A(\mem<9><5> ), .B(n389), .C(\mem<8><5> ), .D(n391), .Y(
        n3978) );
  AOI22X1 U2026 ( .A(\mem<23><5> ), .B(n385), .C(\mem<22><5> ), .D(n388), .Y(
        n3969) );
  AOI22X1 U2027 ( .A(\mem<21><5> ), .B(n381), .C(\mem<20><5> ), .D(n384), .Y(
        n3970) );
  AOI22X1 U2028 ( .A(\mem<19><5> ), .B(n377), .C(\mem<18><5> ), .D(n380), .Y(
        n3972) );
  AOI22X1 U2029 ( .A(\mem<17><5> ), .B(n373), .C(\mem<16><5> ), .D(n376), .Y(
        n3973) );
  AOI22X1 U2031 ( .A(\mem<31><5> ), .B(n369), .C(\mem<30><5> ), .D(n371), .Y(
        n3964) );
  AOI22X1 U2032 ( .A(\mem<29><5> ), .B(n365), .C(\mem<28><5> ), .D(n367), .Y(
        n3965) );
  AOI22X1 U2033 ( .A(\mem<27><5> ), .B(n361), .C(\mem<26><5> ), .D(n363), .Y(
        n3967) );
  AOI22X1 U2034 ( .A(\mem<25><5> ), .B(n357), .C(\mem<24><5> ), .D(n359), .Y(
        n3968) );
  AOI21X1 U2035 ( .A(n3963), .B(n3962), .C(n2609), .Y(n4805) );
  NOR3X1 U2036 ( .A(n3961), .B(n126), .C(n246), .Y(n3962) );
  AOI22X1 U2038 ( .A(\mem<55><4> ), .B(n473), .C(\mem<54><4> ), .D(n475), .Y(
        n3956) );
  AOI22X1 U2039 ( .A(\mem<53><4> ), .B(n469), .C(\mem<52><4> ), .D(n471), .Y(
        n3957) );
  AOI22X1 U2040 ( .A(\mem<51><4> ), .B(n465), .C(\mem<50><4> ), .D(n467), .Y(
        n3959) );
  AOI22X1 U2041 ( .A(\mem<49><4> ), .B(n461), .C(\mem<48><4> ), .D(n463), .Y(
        n3960) );
  AOI22X1 U2043 ( .A(\mem<63><4> ), .B(n356), .C(\mem<62><4> ), .D(n459), .Y(
        n3951) );
  AOI22X1 U2044 ( .A(\mem<61><4> ), .B(n456), .C(\mem<60><4> ), .D(n457), .Y(
        n3952) );
  AOI22X1 U2045 ( .A(\mem<59><4> ), .B(n452), .C(\mem<58><4> ), .D(n453), .Y(
        n3954) );
  AOI22X1 U2046 ( .A(\mem<57><4> ), .B(n448), .C(\mem<56><4> ), .D(n449), .Y(
        n3955) );
  AOI22X1 U2048 ( .A(\mem<39><4> ), .B(n443), .C(\mem<38><4> ), .D(n446), .Y(
        n3946) );
  AOI22X1 U2049 ( .A(\mem<37><4> ), .B(n439), .C(\mem<36><4> ), .D(n442), .Y(
        n3947) );
  AOI22X1 U2050 ( .A(\mem<35><4> ), .B(n435), .C(\mem<34><4> ), .D(n437), .Y(
        n3949) );
  AOI22X1 U2051 ( .A(\mem<33><4> ), .B(n431), .C(\mem<32><4> ), .D(n433), .Y(
        n3950) );
  AOI22X1 U2053 ( .A(\mem<47><4> ), .B(n427), .C(\mem<46><4> ), .D(n429), .Y(
        n3941) );
  AOI22X1 U2054 ( .A(\mem<45><4> ), .B(n423), .C(\mem<44><4> ), .D(n425), .Y(
        n3942) );
  AOI22X1 U2055 ( .A(\mem<43><4> ), .B(n419), .C(\mem<42><4> ), .D(n421), .Y(
        n3944) );
  AOI22X1 U2056 ( .A(\mem<41><4> ), .B(n415), .C(\mem<40><4> ), .D(n417), .Y(
        n3945) );
  NOR3X1 U2057 ( .A(n3940), .B(n220), .C(n244), .Y(n3963) );
  AOI22X1 U2059 ( .A(\mem<7><4> ), .B(n3192), .C(\mem<6><4> ), .D(n413), .Y(
        n3935) );
  AOI22X1 U2060 ( .A(\mem<5><4> ), .B(n3193), .C(\mem<4><4> ), .D(n409), .Y(
        n3936) );
  AOI22X1 U2061 ( .A(\mem<3><4> ), .B(n3194), .C(\mem<2><4> ), .D(n477), .Y(
        n3938) );
  AOI22X1 U2062 ( .A(\mem<1><4> ), .B(n351), .C(n4067), .D(\mem<0><4> ), .Y(
        n3939) );
  AOI22X1 U2064 ( .A(\mem<15><4> ), .B(n401), .C(\mem<14><4> ), .D(n404), .Y(
        n3930) );
  AOI22X1 U2065 ( .A(\mem<13><4> ), .B(n397), .C(\mem<12><4> ), .D(n400), .Y(
        n3931) );
  AOI22X1 U2066 ( .A(\mem<11><4> ), .B(n393), .C(\mem<10><4> ), .D(n396), .Y(
        n3933) );
  AOI22X1 U2067 ( .A(\mem<9><4> ), .B(n389), .C(\mem<8><4> ), .D(n391), .Y(
        n3934) );
  AOI22X1 U2069 ( .A(\mem<23><4> ), .B(n385), .C(\mem<22><4> ), .D(n388), .Y(
        n3925) );
  AOI22X1 U2070 ( .A(\mem<21><4> ), .B(n381), .C(\mem<20><4> ), .D(n384), .Y(
        n3926) );
  AOI22X1 U2071 ( .A(\mem<19><4> ), .B(n377), .C(\mem<18><4> ), .D(n380), .Y(
        n3928) );
  AOI22X1 U2072 ( .A(\mem<17><4> ), .B(n373), .C(\mem<16><4> ), .D(n376), .Y(
        n3929) );
  AOI22X1 U2074 ( .A(\mem<31><4> ), .B(n369), .C(\mem<30><4> ), .D(n371), .Y(
        n3920) );
  AOI22X1 U2075 ( .A(\mem<29><4> ), .B(n365), .C(\mem<28><4> ), .D(n367), .Y(
        n3921) );
  AOI22X1 U2076 ( .A(\mem<27><4> ), .B(n361), .C(\mem<26><4> ), .D(n363), .Y(
        n3923) );
  AOI22X1 U2077 ( .A(\mem<25><4> ), .B(n357), .C(\mem<24><4> ), .D(n359), .Y(
        n3924) );
  AOI21X1 U2078 ( .A(n3919), .B(n3918), .C(n2609), .Y(n4806) );
  NOR3X1 U2079 ( .A(n3917), .B(n101), .C(n242), .Y(n3918) );
  AOI22X1 U2081 ( .A(\mem<55><3> ), .B(n473), .C(\mem<54><3> ), .D(n475), .Y(
        n3912) );
  AOI22X1 U2082 ( .A(\mem<53><3> ), .B(n469), .C(\mem<52><3> ), .D(n471), .Y(
        n3913) );
  AOI22X1 U2083 ( .A(\mem<51><3> ), .B(n465), .C(\mem<50><3> ), .D(n467), .Y(
        n3915) );
  AOI22X1 U2084 ( .A(\mem<49><3> ), .B(n461), .C(\mem<48><3> ), .D(n463), .Y(
        n3916) );
  AOI22X1 U2086 ( .A(\mem<63><3> ), .B(n356), .C(\mem<62><3> ), .D(n459), .Y(
        n3907) );
  AOI22X1 U2087 ( .A(\mem<61><3> ), .B(n456), .C(\mem<60><3> ), .D(n457), .Y(
        n3908) );
  AOI22X1 U2088 ( .A(\mem<59><3> ), .B(n452), .C(\mem<58><3> ), .D(n453), .Y(
        n3910) );
  AOI22X1 U2089 ( .A(\mem<57><3> ), .B(n448), .C(\mem<56><3> ), .D(n449), .Y(
        n3911) );
  AOI22X1 U2091 ( .A(\mem<39><3> ), .B(n443), .C(\mem<38><3> ), .D(n446), .Y(
        n3902) );
  AOI22X1 U2092 ( .A(\mem<37><3> ), .B(n439), .C(\mem<36><3> ), .D(n442), .Y(
        n3903) );
  AOI22X1 U2093 ( .A(\mem<35><3> ), .B(n435), .C(\mem<34><3> ), .D(n437), .Y(
        n3905) );
  AOI22X1 U2094 ( .A(\mem<33><3> ), .B(n431), .C(\mem<32><3> ), .D(n433), .Y(
        n3906) );
  AOI22X1 U2096 ( .A(\mem<47><3> ), .B(n427), .C(\mem<46><3> ), .D(n429), .Y(
        n3897) );
  AOI22X1 U2097 ( .A(\mem<45><3> ), .B(n423), .C(\mem<44><3> ), .D(n425), .Y(
        n3898) );
  AOI22X1 U2098 ( .A(\mem<43><3> ), .B(n419), .C(\mem<42><3> ), .D(n421), .Y(
        n3900) );
  AOI22X1 U2099 ( .A(\mem<41><3> ), .B(n415), .C(\mem<40><3> ), .D(n417), .Y(
        n3901) );
  NOR3X1 U2100 ( .A(n3896), .B(n218), .C(n240), .Y(n3919) );
  AOI22X1 U2102 ( .A(\mem<7><3> ), .B(n3192), .C(\mem<6><3> ), .D(n413), .Y(
        n3891) );
  AOI22X1 U2103 ( .A(\mem<5><3> ), .B(n3193), .C(\mem<4><3> ), .D(n409), .Y(
        n3892) );
  AOI22X1 U2104 ( .A(\mem<3><3> ), .B(n3194), .C(\mem<2><3> ), .D(n477), .Y(
        n3894) );
  AOI22X1 U2105 ( .A(\mem<1><3> ), .B(n351), .C(n4067), .D(\mem<0><3> ), .Y(
        n3895) );
  AOI22X1 U2107 ( .A(\mem<15><3> ), .B(n401), .C(\mem<14><3> ), .D(n404), .Y(
        n3886) );
  AOI22X1 U2108 ( .A(\mem<13><3> ), .B(n397), .C(\mem<12><3> ), .D(n400), .Y(
        n3887) );
  AOI22X1 U2109 ( .A(\mem<11><3> ), .B(n393), .C(\mem<10><3> ), .D(n396), .Y(
        n3889) );
  AOI22X1 U2110 ( .A(\mem<9><3> ), .B(n389), .C(\mem<8><3> ), .D(n391), .Y(
        n3890) );
  AOI22X1 U2112 ( .A(\mem<23><3> ), .B(n385), .C(\mem<22><3> ), .D(n388), .Y(
        n3881) );
  AOI22X1 U2113 ( .A(\mem<21><3> ), .B(n381), .C(\mem<20><3> ), .D(n384), .Y(
        n3882) );
  AOI22X1 U2114 ( .A(\mem<19><3> ), .B(n377), .C(\mem<18><3> ), .D(n380), .Y(
        n3884) );
  AOI22X1 U2115 ( .A(\mem<17><3> ), .B(n373), .C(\mem<16><3> ), .D(n376), .Y(
        n3885) );
  AOI22X1 U2117 ( .A(\mem<31><3> ), .B(n369), .C(\mem<30><3> ), .D(n371), .Y(
        n3876) );
  AOI22X1 U2118 ( .A(\mem<29><3> ), .B(n365), .C(\mem<28><3> ), .D(n367), .Y(
        n3877) );
  AOI22X1 U2119 ( .A(\mem<27><3> ), .B(n361), .C(\mem<26><3> ), .D(n363), .Y(
        n3879) );
  AOI22X1 U2120 ( .A(\mem<25><3> ), .B(n357), .C(\mem<24><3> ), .D(n359), .Y(
        n3880) );
  AOI21X1 U2121 ( .A(n3875), .B(n3874), .C(n2609), .Y(n4807) );
  NOR3X1 U2122 ( .A(n3873), .B(n76), .C(n238), .Y(n3874) );
  AOI22X1 U2124 ( .A(\mem<55><2> ), .B(n473), .C(\mem<54><2> ), .D(n475), .Y(
        n3868) );
  AOI22X1 U2125 ( .A(\mem<53><2> ), .B(n469), .C(\mem<52><2> ), .D(n471), .Y(
        n3869) );
  AOI22X1 U2126 ( .A(\mem<51><2> ), .B(n465), .C(\mem<50><2> ), .D(n467), .Y(
        n3871) );
  AOI22X1 U2127 ( .A(\mem<49><2> ), .B(n461), .C(\mem<48><2> ), .D(n463), .Y(
        n3872) );
  AOI22X1 U2129 ( .A(\mem<63><2> ), .B(n356), .C(\mem<62><2> ), .D(n459), .Y(
        n3863) );
  AOI22X1 U2130 ( .A(\mem<61><2> ), .B(n456), .C(\mem<60><2> ), .D(n457), .Y(
        n3864) );
  AOI22X1 U2131 ( .A(\mem<59><2> ), .B(n452), .C(\mem<58><2> ), .D(n453), .Y(
        n3866) );
  AOI22X1 U2132 ( .A(\mem<57><2> ), .B(n448), .C(\mem<56><2> ), .D(n449), .Y(
        n3867) );
  AOI22X1 U2134 ( .A(\mem<39><2> ), .B(n443), .C(\mem<38><2> ), .D(n446), .Y(
        n3858) );
  AOI22X1 U2135 ( .A(\mem<37><2> ), .B(n439), .C(\mem<36><2> ), .D(n442), .Y(
        n3859) );
  AOI22X1 U2136 ( .A(\mem<35><2> ), .B(n435), .C(\mem<34><2> ), .D(n437), .Y(
        n3861) );
  AOI22X1 U2137 ( .A(\mem<33><2> ), .B(n431), .C(\mem<32><2> ), .D(n433), .Y(
        n3862) );
  AOI22X1 U2139 ( .A(\mem<47><2> ), .B(n427), .C(\mem<46><2> ), .D(n429), .Y(
        n3853) );
  AOI22X1 U2140 ( .A(\mem<45><2> ), .B(n423), .C(\mem<44><2> ), .D(n425), .Y(
        n3854) );
  AOI22X1 U2141 ( .A(\mem<43><2> ), .B(n419), .C(\mem<42><2> ), .D(n421), .Y(
        n3856) );
  AOI22X1 U2142 ( .A(\mem<41><2> ), .B(n415), .C(\mem<40><2> ), .D(n417), .Y(
        n3857) );
  NOR3X1 U2143 ( .A(n3852), .B(n216), .C(n236), .Y(n3875) );
  AOI22X1 U2145 ( .A(\mem<7><2> ), .B(n3192), .C(\mem<6><2> ), .D(n413), .Y(
        n3847) );
  AOI22X1 U2146 ( .A(\mem<5><2> ), .B(n3193), .C(\mem<4><2> ), .D(n409), .Y(
        n3848) );
  AOI22X1 U2147 ( .A(\mem<3><2> ), .B(n3194), .C(\mem<2><2> ), .D(n477), .Y(
        n3850) );
  AOI22X1 U2148 ( .A(\mem<1><2> ), .B(n351), .C(n4067), .D(\mem<0><2> ), .Y(
        n3851) );
  AOI22X1 U2150 ( .A(\mem<15><2> ), .B(n401), .C(\mem<14><2> ), .D(n404), .Y(
        n3842) );
  AOI22X1 U2151 ( .A(\mem<13><2> ), .B(n397), .C(\mem<12><2> ), .D(n400), .Y(
        n3843) );
  AOI22X1 U2152 ( .A(\mem<11><2> ), .B(n393), .C(\mem<10><2> ), .D(n396), .Y(
        n3845) );
  AOI22X1 U2153 ( .A(\mem<9><2> ), .B(n389), .C(\mem<8><2> ), .D(n391), .Y(
        n3846) );
  AOI22X1 U2155 ( .A(\mem<23><2> ), .B(n385), .C(\mem<22><2> ), .D(n388), .Y(
        n3837) );
  AOI22X1 U2156 ( .A(\mem<21><2> ), .B(n381), .C(\mem<20><2> ), .D(n384), .Y(
        n3838) );
  AOI22X1 U2157 ( .A(\mem<19><2> ), .B(n377), .C(\mem<18><2> ), .D(n380), .Y(
        n3840) );
  AOI22X1 U2158 ( .A(\mem<17><2> ), .B(n373), .C(\mem<16><2> ), .D(n376), .Y(
        n3841) );
  AOI22X1 U2160 ( .A(\mem<31><2> ), .B(n369), .C(\mem<30><2> ), .D(n371), .Y(
        n3832) );
  AOI22X1 U2161 ( .A(\mem<29><2> ), .B(n365), .C(\mem<28><2> ), .D(n367), .Y(
        n3833) );
  AOI22X1 U2162 ( .A(\mem<27><2> ), .B(n361), .C(\mem<26><2> ), .D(n363), .Y(
        n3835) );
  AOI22X1 U2163 ( .A(\mem<25><2> ), .B(n357), .C(\mem<24><2> ), .D(n359), .Y(
        n3836) );
  AOI21X1 U2164 ( .A(n3831), .B(n3830), .C(n2609), .Y(n4808) );
  NOR3X1 U2165 ( .A(n3829), .B(n51), .C(n234), .Y(n3830) );
  AOI22X1 U2167 ( .A(\mem<55><1> ), .B(n473), .C(\mem<54><1> ), .D(n475), .Y(
        n3824) );
  AOI22X1 U2168 ( .A(\mem<53><1> ), .B(n469), .C(\mem<52><1> ), .D(n471), .Y(
        n3825) );
  AOI22X1 U2169 ( .A(\mem<51><1> ), .B(n465), .C(\mem<50><1> ), .D(n467), .Y(
        n3827) );
  AOI22X1 U2170 ( .A(\mem<49><1> ), .B(n461), .C(\mem<48><1> ), .D(n463), .Y(
        n3828) );
  AOI22X1 U2172 ( .A(\mem<63><1> ), .B(n356), .C(\mem<62><1> ), .D(n459), .Y(
        n3819) );
  AOI22X1 U2173 ( .A(\mem<61><1> ), .B(n456), .C(\mem<60><1> ), .D(n457), .Y(
        n3820) );
  AOI22X1 U2174 ( .A(\mem<59><1> ), .B(n452), .C(\mem<58><1> ), .D(n453), .Y(
        n3822) );
  AOI22X1 U2175 ( .A(\mem<57><1> ), .B(n448), .C(\mem<56><1> ), .D(n449), .Y(
        n3823) );
  AOI22X1 U2177 ( .A(\mem<39><1> ), .B(n443), .C(\mem<38><1> ), .D(n446), .Y(
        n3814) );
  AOI22X1 U2178 ( .A(\mem<37><1> ), .B(n439), .C(\mem<36><1> ), .D(n442), .Y(
        n3815) );
  AOI22X1 U2179 ( .A(\mem<35><1> ), .B(n435), .C(\mem<34><1> ), .D(n437), .Y(
        n3817) );
  AOI22X1 U2180 ( .A(\mem<33><1> ), .B(n431), .C(\mem<32><1> ), .D(n433), .Y(
        n3818) );
  AOI22X1 U2182 ( .A(\mem<47><1> ), .B(n427), .C(\mem<46><1> ), .D(n429), .Y(
        n3809) );
  AOI22X1 U2183 ( .A(\mem<45><1> ), .B(n423), .C(\mem<44><1> ), .D(n425), .Y(
        n3810) );
  AOI22X1 U2184 ( .A(\mem<43><1> ), .B(n419), .C(\mem<42><1> ), .D(n421), .Y(
        n3812) );
  AOI22X1 U2185 ( .A(\mem<41><1> ), .B(n415), .C(\mem<40><1> ), .D(n417), .Y(
        n3813) );
  NOR3X1 U2186 ( .A(n3808), .B(n214), .C(n232), .Y(n3831) );
  AOI22X1 U2188 ( .A(\mem<7><1> ), .B(n3192), .C(\mem<6><1> ), .D(n413), .Y(
        n3803) );
  AOI22X1 U2189 ( .A(\mem<5><1> ), .B(n3193), .C(\mem<4><1> ), .D(n409), .Y(
        n3804) );
  AOI22X1 U2190 ( .A(\mem<3><1> ), .B(n3194), .C(\mem<2><1> ), .D(n477), .Y(
        n3806) );
  AOI22X1 U2191 ( .A(\mem<1><1> ), .B(n351), .C(n4067), .D(\mem<0><1> ), .Y(
        n3807) );
  AOI22X1 U2193 ( .A(\mem<15><1> ), .B(n401), .C(\mem<14><1> ), .D(n404), .Y(
        n3798) );
  AOI22X1 U2194 ( .A(\mem<13><1> ), .B(n397), .C(\mem<12><1> ), .D(n400), .Y(
        n3799) );
  AOI22X1 U2195 ( .A(\mem<11><1> ), .B(n393), .C(\mem<10><1> ), .D(n396), .Y(
        n3801) );
  AOI22X1 U2196 ( .A(\mem<9><1> ), .B(n389), .C(\mem<8><1> ), .D(n391), .Y(
        n3802) );
  AOI22X1 U2198 ( .A(\mem<23><1> ), .B(n385), .C(\mem<22><1> ), .D(n388), .Y(
        n3793) );
  AOI22X1 U2199 ( .A(\mem<21><1> ), .B(n381), .C(\mem<20><1> ), .D(n384), .Y(
        n3794) );
  AOI22X1 U2200 ( .A(\mem<19><1> ), .B(n377), .C(\mem<18><1> ), .D(n380), .Y(
        n3796) );
  AOI22X1 U2201 ( .A(\mem<17><1> ), .B(n373), .C(\mem<16><1> ), .D(n376), .Y(
        n3797) );
  AOI22X1 U2203 ( .A(\mem<31><1> ), .B(n369), .C(\mem<30><1> ), .D(n371), .Y(
        n3788) );
  AOI22X1 U2204 ( .A(\mem<29><1> ), .B(n365), .C(\mem<28><1> ), .D(n367), .Y(
        n3789) );
  AOI22X1 U2205 ( .A(\mem<27><1> ), .B(n361), .C(\mem<26><1> ), .D(n363), .Y(
        n3791) );
  AOI22X1 U2206 ( .A(\mem<25><1> ), .B(n357), .C(\mem<24><1> ), .D(n359), .Y(
        n3792) );
  AOI21X1 U2207 ( .A(n3787), .B(n3786), .C(n2609), .Y(n4809) );
  NAND2X1 U2208 ( .A(enable), .B(n3205), .Y(n4095) );
  NOR3X1 U2209 ( .A(n3785), .B(n26), .C(n230), .Y(n3786) );
  AOI22X1 U2211 ( .A(\mem<55><0> ), .B(n473), .C(\mem<54><0> ), .D(n475), .Y(
        n3780) );
  AOI22X1 U2214 ( .A(\mem<53><0> ), .B(n469), .C(\mem<52><0> ), .D(n471), .Y(
        n3781) );
  AOI22X1 U2217 ( .A(\mem<51><0> ), .B(n465), .C(\mem<50><0> ), .D(n467), .Y(
        n3783) );
  AOI22X1 U2220 ( .A(\mem<49><0> ), .B(n461), .C(\mem<48><0> ), .D(n463), .Y(
        n3784) );
  AOI22X1 U2224 ( .A(\mem<63><0> ), .B(n356), .C(\mem<62><0> ), .D(n459), .Y(
        n3768) );
  AOI22X1 U2227 ( .A(\mem<61><0> ), .B(n456), .C(\mem<60><0> ), .D(n457), .Y(
        n3769) );
  AOI22X1 U2230 ( .A(\mem<59><0> ), .B(n452), .C(\mem<58><0> ), .D(n453), .Y(
        n3771) );
  AOI22X1 U2233 ( .A(\mem<57><0> ), .B(n448), .C(\mem<56><0> ), .D(n449), .Y(
        n3772) );
  NAND3X1 U2235 ( .A(n3766), .B(N182), .C(n3765), .Y(n3767) );
  AOI22X1 U2239 ( .A(\mem<39><0> ), .B(n443), .C(\mem<38><0> ), .D(n446), .Y(
        n3760) );
  AOI22X1 U2242 ( .A(\mem<37><0> ), .B(n439), .C(\mem<36><0> ), .D(n442), .Y(
        n3761) );
  AOI22X1 U2245 ( .A(\mem<35><0> ), .B(n435), .C(\mem<34><0> ), .D(n437), .Y(
        n3763) );
  AOI22X1 U2248 ( .A(\mem<33><0> ), .B(n431), .C(\mem<32><0> ), .D(n433), .Y(
        n3764) );
  AOI22X1 U2252 ( .A(\mem<47><0> ), .B(n427), .C(\mem<46><0> ), .D(n429), .Y(
        n3755) );
  AOI22X1 U2255 ( .A(\mem<45><0> ), .B(n423), .C(\mem<44><0> ), .D(n425), .Y(
        n3756) );
  AOI22X1 U2258 ( .A(\mem<43><0> ), .B(n419), .C(\mem<42><0> ), .D(n421), .Y(
        n3758) );
  AOI22X1 U2261 ( .A(\mem<41><0> ), .B(n415), .C(\mem<40><0> ), .D(n417), .Y(
        n3759) );
  NAND3X1 U2263 ( .A(n3766), .B(N182), .C(n276), .Y(n3754) );
  NAND3X1 U2266 ( .A(n3766), .B(N182), .C(n274), .Y(n3753) );
  NOR3X1 U2268 ( .A(n3752), .B(n212), .C(n228), .Y(n3787) );
  AOI22X1 U2270 ( .A(\mem<7><0> ), .B(n3192), .C(\mem<6><0> ), .D(n413), .Y(
        n3747) );
  AOI22X1 U2273 ( .A(\mem<5><0> ), .B(n3193), .C(\mem<4><0> ), .D(n409), .Y(
        n3748) );
  AOI22X1 U2276 ( .A(\mem<3><0> ), .B(n3194), .C(\mem<2><0> ), .D(n477), .Y(
        n3750) );
  AOI22X1 U2279 ( .A(\mem<1><0> ), .B(n351), .C(n4067), .D(\mem<0><0> ), .Y(
        n3751) );
  NOR3X1 U2280 ( .A(n3746), .B(n1), .C(n3745), .Y(n4067) );
  NAND3X1 U2281 ( .A(\addr<8> ), .B(\addr<7> ), .C(\addr<9> ), .Y(n3743) );
  NAND3X1 U2282 ( .A(\addr<15> ), .B(\addr<14> ), .C(\addr<6> ), .Y(n3744) );
  NAND3X1 U2284 ( .A(N181), .B(N180), .C(N182), .Y(n3742) );
  NAND3X1 U2285 ( .A(\addr<13> ), .B(\addr<11> ), .C(\addr<12> ), .Y(n3746) );
  AOI22X1 U2288 ( .A(\mem<15><0> ), .B(n401), .C(\mem<14><0> ), .D(n404), .Y(
        n3737) );
  AOI22X1 U2291 ( .A(\mem<13><0> ), .B(n397), .C(\mem<12><0> ), .D(n400), .Y(
        n3738) );
  AOI22X1 U2294 ( .A(\mem<11><0> ), .B(n393), .C(\mem<10><0> ), .D(n396), .Y(
        n3740) );
  AOI22X1 U2297 ( .A(\mem<9><0> ), .B(n389), .C(\mem<8><0> ), .D(n391), .Y(
        n3741) );
  AOI22X1 U2302 ( .A(\mem<23><0> ), .B(n385), .C(\mem<22><0> ), .D(n388), .Y(
        n3731) );
  AOI22X1 U2305 ( .A(\mem<21><0> ), .B(n381), .C(\mem<20><0> ), .D(n384), .Y(
        n3732) );
  AOI22X1 U2308 ( .A(\mem<19><0> ), .B(n377), .C(\mem<18><0> ), .D(n380), .Y(
        n3734) );
  AOI22X1 U2311 ( .A(\mem<17><0> ), .B(n373), .C(\mem<16><0> ), .D(n376), .Y(
        n3735) );
  NOR2X1 U2314 ( .A(N182), .B(N181), .Y(n3736) );
  AOI22X1 U2317 ( .A(\mem<31><0> ), .B(n369), .C(\mem<30><0> ), .D(n371), .Y(
        n3726) );
  NOR3X1 U2319 ( .A(n2677), .B(N178), .C(n2675), .Y(n3779) );
  NOR3X1 U2321 ( .A(n2676), .B(N177), .C(n2677), .Y(n3778) );
  AOI22X1 U2322 ( .A(\mem<29><0> ), .B(n365), .C(\mem<28><0> ), .D(n367), .Y(
        n3727) );
  NOR3X1 U2324 ( .A(n2676), .B(N179), .C(n2675), .Y(n3777) );
  NOR3X1 U2326 ( .A(N177), .B(N178), .C(n2677), .Y(n3776) );
  AOI22X1 U2327 ( .A(\mem<27><0> ), .B(n361), .C(\mem<26><0> ), .D(n363), .Y(
        n3729) );
  NOR3X1 U2329 ( .A(N178), .B(N179), .C(n2675), .Y(n3775) );
  NOR3X1 U2331 ( .A(N177), .B(N179), .C(n2676), .Y(n3774) );
  AOI22X1 U2332 ( .A(\mem<25><0> ), .B(n357), .C(\mem<24><0> ), .D(n359), .Y(
        n3730) );
  NAND3X1 U2334 ( .A(N179), .B(N178), .C(N177), .Y(n4789) );
  NAND3X1 U2335 ( .A(n3766), .B(N181), .C(n3724), .Y(n3725) );
  NOR2X1 U2336 ( .A(N182), .B(N180), .Y(n3724) );
  NOR3X1 U2338 ( .A(N178), .B(N179), .C(N177), .Y(n3773) );
  NAND3X1 U2339 ( .A(n3766), .B(N181), .C(n3722), .Y(n3723) );
  NOR2X1 U2340 ( .A(N182), .B(n2678), .Y(n3722) );
  NOR3X1 U2341 ( .A(n3202), .B(\addr<6> ), .C(\addr<15> ), .Y(n3720) );
  NOR3X1 U2342 ( .A(\addr<8> ), .B(\addr<9> ), .C(\addr<7> ), .Y(n3719) );
  NOR3X1 U2343 ( .A(n3203), .B(\addr<11> ), .C(\addr<10> ), .Y(n3721) );
  NOR3X1 U2344 ( .A(\addr<13> ), .B(\addr<14> ), .C(\addr<12> ), .Y(n3718) );
  INVX1 U3 ( .A(n3718), .Y(n3203) );
  INVX1 U4 ( .A(n2609), .Y(n3204) );
  BUFX2 U5 ( .A(n4116), .Y(n2610) );
  OR2X1 U6 ( .A(n13), .B(n14), .Y(n12) );
  OR2X1 U7 ( .A(n23), .B(n24), .Y(n22) );
  OR2X1 U8 ( .A(n38), .B(n39), .Y(n37) );
  OR2X1 U9 ( .A(n48), .B(n49), .Y(n47) );
  OR2X1 U10 ( .A(n63), .B(n64), .Y(n62) );
  OR2X1 U11 ( .A(n73), .B(n74), .Y(n72) );
  OR2X1 U12 ( .A(n88), .B(n89), .Y(n87) );
  OR2X1 U13 ( .A(n98), .B(n99), .Y(n97) );
  OR2X1 U14 ( .A(n113), .B(n114), .Y(n112) );
  OR2X1 U15 ( .A(n123), .B(n124), .Y(n122) );
  OR2X1 U16 ( .A(n138), .B(n139), .Y(n137) );
  OR2X1 U17 ( .A(n148), .B(n149), .Y(n147) );
  OR2X1 U18 ( .A(n163), .B(n164), .Y(n162) );
  OR2X1 U19 ( .A(n173), .B(n174), .Y(n172) );
  OR2X1 U20 ( .A(n188), .B(n189), .Y(n187) );
  OR2X1 U21 ( .A(n198), .B(n199), .Y(n197) );
  INVX1 U22 ( .A(n412), .Y(n3192) );
  INVX1 U23 ( .A(n408), .Y(n3193) );
  INVX1 U24 ( .A(n406), .Y(n3194) );
  AND2X1 U25 ( .A(n2674), .B(n4790), .Y(n4801) );
  AND2X1 U26 ( .A(n4801), .B(n355), .Y(n4799) );
  AND2X1 U27 ( .A(n356), .B(n4801), .Y(n4798) );
  AND2X1 U28 ( .A(n2671), .B(n460), .Y(n4786) );
  AND2X1 U29 ( .A(n459), .B(n2671), .Y(n4785) );
  AND2X1 U30 ( .A(n2670), .B(n455), .Y(n4774) );
  AND2X1 U31 ( .A(n456), .B(n2670), .Y(n4773) );
  AND2X1 U32 ( .A(n2669), .B(n458), .Y(n4763) );
  AND2X1 U33 ( .A(n457), .B(n2669), .Y(n4762) );
  AND2X1 U34 ( .A(n2668), .B(n451), .Y(n4752) );
  AND2X1 U35 ( .A(n452), .B(n2668), .Y(n4751) );
  AND2X1 U36 ( .A(n2667), .B(n454), .Y(n4741) );
  AND2X1 U37 ( .A(n453), .B(n2667), .Y(n4740) );
  AND2X1 U38 ( .A(n2666), .B(n447), .Y(n4730) );
  AND2X1 U39 ( .A(n448), .B(n2666), .Y(n4729) );
  AND2X1 U40 ( .A(n2665), .B(n450), .Y(n4719) );
  AND2X1 U41 ( .A(n449), .B(n2665), .Y(n4718) );
  AND2X1 U42 ( .A(n2664), .B(n474), .Y(n4708) );
  AND2X1 U43 ( .A(n473), .B(n2664), .Y(n4707) );
  AND2X1 U44 ( .A(n2663), .B(n476), .Y(n4697) );
  AND2X1 U45 ( .A(n475), .B(n2663), .Y(n4696) );
  AND2X1 U46 ( .A(n2662), .B(n470), .Y(n4686) );
  AND2X1 U47 ( .A(n469), .B(n2662), .Y(n4685) );
  AND2X1 U48 ( .A(n2661), .B(n472), .Y(n4675) );
  AND2X1 U49 ( .A(n471), .B(n2661), .Y(n4674) );
  AND2X1 U50 ( .A(n2660), .B(n466), .Y(n4664) );
  AND2X1 U51 ( .A(n465), .B(n2660), .Y(n4663) );
  AND2X1 U52 ( .A(n2659), .B(n468), .Y(n4653) );
  AND2X1 U53 ( .A(n467), .B(n2659), .Y(n4652) );
  AND2X1 U54 ( .A(n2658), .B(n462), .Y(n4642) );
  AND2X1 U55 ( .A(n461), .B(n2658), .Y(n4641) );
  AND2X1 U56 ( .A(n2657), .B(n464), .Y(n4631) );
  AND2X1 U57 ( .A(n463), .B(n2657), .Y(n4630) );
  AND2X1 U58 ( .A(n2656), .B(n428), .Y(n4620) );
  AND2X1 U59 ( .A(n427), .B(n2656), .Y(n4619) );
  AND2X1 U60 ( .A(n2655), .B(n430), .Y(n4609) );
  AND2X1 U61 ( .A(n429), .B(n2655), .Y(n4608) );
  AND2X1 U62 ( .A(n2654), .B(n424), .Y(n4598) );
  AND2X1 U63 ( .A(n423), .B(n2654), .Y(n4597) );
  AND2X1 U64 ( .A(n2653), .B(n426), .Y(n4587) );
  AND2X1 U65 ( .A(n425), .B(n2653), .Y(n4586) );
  AND2X1 U66 ( .A(n2652), .B(n420), .Y(n4576) );
  AND2X1 U67 ( .A(n419), .B(n2652), .Y(n4575) );
  AND2X1 U68 ( .A(n2651), .B(n422), .Y(n4565) );
  AND2X1 U69 ( .A(n421), .B(n2651), .Y(n4564) );
  AND2X1 U70 ( .A(n2650), .B(n416), .Y(n4554) );
  AND2X1 U71 ( .A(n415), .B(n2650), .Y(n4553) );
  AND2X1 U72 ( .A(n2649), .B(n418), .Y(n4543) );
  AND2X1 U73 ( .A(n417), .B(n2649), .Y(n4542) );
  AND2X1 U74 ( .A(n2648), .B(n444), .Y(n4532) );
  AND2X1 U75 ( .A(n443), .B(n2648), .Y(n4531) );
  AND2X1 U76 ( .A(n2647), .B(n445), .Y(n4521) );
  AND2X1 U77 ( .A(n446), .B(n2647), .Y(n4520) );
  AND2X1 U78 ( .A(n2646), .B(n440), .Y(n4510) );
  AND2X1 U79 ( .A(n439), .B(n2646), .Y(n4509) );
  AND2X1 U80 ( .A(n2645), .B(n441), .Y(n4499) );
  AND2X1 U81 ( .A(n442), .B(n2645), .Y(n4498) );
  AND2X1 U82 ( .A(n2644), .B(n436), .Y(n4488) );
  AND2X1 U83 ( .A(n435), .B(n2644), .Y(n4487) );
  AND2X1 U84 ( .A(n2643), .B(n438), .Y(n4477) );
  AND2X1 U85 ( .A(n437), .B(n2643), .Y(n4476) );
  AND2X1 U86 ( .A(n2642), .B(n432), .Y(n4466) );
  AND2X1 U87 ( .A(n431), .B(n2642), .Y(n4465) );
  AND2X1 U88 ( .A(n2641), .B(n434), .Y(n4455) );
  AND2X1 U89 ( .A(n433), .B(n2641), .Y(n4454) );
  AND2X1 U90 ( .A(n2640), .B(n370), .Y(n4444) );
  AND2X1 U91 ( .A(n369), .B(n2640), .Y(n4443) );
  AND2X1 U92 ( .A(n2639), .B(n372), .Y(n4433) );
  AND2X1 U93 ( .A(n371), .B(n2639), .Y(n4432) );
  AND2X1 U94 ( .A(n2638), .B(n366), .Y(n4422) );
  AND2X1 U95 ( .A(n365), .B(n2638), .Y(n4421) );
  AND2X1 U96 ( .A(n2637), .B(n368), .Y(n4411) );
  AND2X1 U97 ( .A(n367), .B(n2637), .Y(n4410) );
  AND2X1 U98 ( .A(n2636), .B(n362), .Y(n4400) );
  AND2X1 U99 ( .A(n361), .B(n2636), .Y(n4399) );
  AND2X1 U100 ( .A(n2635), .B(n364), .Y(n4389) );
  AND2X1 U101 ( .A(n363), .B(n2635), .Y(n4388) );
  AND2X1 U102 ( .A(n2634), .B(n358), .Y(n4378) );
  AND2X1 U103 ( .A(n357), .B(n2634), .Y(n4377) );
  AND2X1 U104 ( .A(n2633), .B(n360), .Y(n4367) );
  AND2X1 U105 ( .A(n359), .B(n2633), .Y(n4366) );
  AND2X1 U106 ( .A(n2632), .B(n386), .Y(n4356) );
  AND2X1 U107 ( .A(n385), .B(n2632), .Y(n4355) );
  AND2X1 U108 ( .A(n2631), .B(n387), .Y(n4345) );
  AND2X1 U109 ( .A(n388), .B(n2631), .Y(n4344) );
  AND2X1 U110 ( .A(n2630), .B(n382), .Y(n4334) );
  AND2X1 U111 ( .A(n381), .B(n2630), .Y(n4333) );
  AND2X1 U112 ( .A(n2629), .B(n383), .Y(n4323) );
  AND2X1 U113 ( .A(n384), .B(n2629), .Y(n4322) );
  AND2X1 U114 ( .A(n2628), .B(n378), .Y(n4312) );
  AND2X1 U115 ( .A(n377), .B(n2628), .Y(n4311) );
  AND2X1 U116 ( .A(n2627), .B(n379), .Y(n4301) );
  AND2X1 U117 ( .A(n380), .B(n2627), .Y(n4300) );
  AND2X1 U118 ( .A(n2626), .B(n374), .Y(n4290) );
  AND2X1 U119 ( .A(n373), .B(n2626), .Y(n4289) );
  AND2X1 U120 ( .A(n2625), .B(n375), .Y(n4279) );
  AND2X1 U121 ( .A(n376), .B(n2625), .Y(n4278) );
  AND2X1 U122 ( .A(n2624), .B(n402), .Y(n4268) );
  AND2X1 U123 ( .A(n401), .B(n2624), .Y(n4267) );
  AND2X1 U124 ( .A(n2623), .B(n403), .Y(n4257) );
  AND2X1 U125 ( .A(n404), .B(n2623), .Y(n4256) );
  AND2X1 U126 ( .A(n2622), .B(n398), .Y(n4246) );
  AND2X1 U127 ( .A(n397), .B(n2622), .Y(n4245) );
  AND2X1 U128 ( .A(n2621), .B(n399), .Y(n4235) );
  AND2X1 U129 ( .A(n400), .B(n2621), .Y(n4234) );
  AND2X1 U130 ( .A(n2620), .B(n394), .Y(n4224) );
  AND2X1 U131 ( .A(n393), .B(n2620), .Y(n4223) );
  AND2X1 U134 ( .A(n2619), .B(n395), .Y(n4213) );
  AND2X1 U139 ( .A(n396), .B(n2619), .Y(n4212) );
  AND2X1 U144 ( .A(n2618), .B(n390), .Y(n4202) );
  AND2X1 U149 ( .A(n389), .B(n2618), .Y(n4201) );
  AND2X1 U154 ( .A(n2617), .B(n392), .Y(n4191) );
  AND2X1 U159 ( .A(n391), .B(n2617), .Y(n4190) );
  AND2X1 U164 ( .A(n2616), .B(n412), .Y(n4180) );
  AND2X1 U169 ( .A(n3192), .B(n2616), .Y(n4179) );
  AND2X1 U174 ( .A(n2615), .B(n414), .Y(n4169) );
  AND2X1 U179 ( .A(n413), .B(n2615), .Y(n4168) );
  AND2X1 U184 ( .A(n2614), .B(n408), .Y(n4158) );
  AND2X1 U189 ( .A(n3193), .B(n2614), .Y(n4157) );
  AND2X1 U194 ( .A(n2613), .B(n410), .Y(n4147) );
  AND2X1 U199 ( .A(n409), .B(n2613), .Y(n4146) );
  AND2X1 U202 ( .A(n2612), .B(n406), .Y(n4136) );
  AND2X1 U203 ( .A(n3194), .B(n2612), .Y(n4135) );
  AND2X1 U204 ( .A(n2611), .B(n478), .Y(n4125) );
  AND2X1 U205 ( .A(n477), .B(n2611), .Y(n4124) );
  AND2X1 U206 ( .A(n2610), .B(n352), .Y(n4114) );
  AND2X1 U207 ( .A(n351), .B(n2610), .Y(n4113) );
  AND2X1 U210 ( .A(N192), .B(n3204), .Y(\data_out<8> ) );
  AND2X1 U211 ( .A(N191), .B(n3204), .Y(\data_out<9> ) );
  AND2X1 U217 ( .A(N190), .B(n3204), .Y(\data_out<10> ) );
  AND2X1 U220 ( .A(N189), .B(n3204), .Y(\data_out<11> ) );
  AND2X1 U221 ( .A(N188), .B(n3204), .Y(\data_out<12> ) );
  AND2X1 U222 ( .A(N187), .B(n3204), .Y(\data_out<13> ) );
  AND2X1 U223 ( .A(N186), .B(n3204), .Y(\data_out<14> ) );
  AND2X1 U224 ( .A(N185), .B(n3204), .Y(\data_out<15> ) );
  INVX1 U225 ( .A(n2608), .Y(n2588) );
  INVX1 U226 ( .A(n2608), .Y(n2587) );
  INVX1 U227 ( .A(n2608), .Y(n2586) );
  INVX1 U228 ( .A(n2608), .Y(n2585) );
  INVX1 U229 ( .A(n3719), .Y(n3202) );
  INVX1 U230 ( .A(n2588), .Y(n2596) );
  INVX1 U231 ( .A(n2588), .Y(n2597) );
  INVX1 U232 ( .A(n2587), .Y(n2600) );
  INVX1 U233 ( .A(n2587), .Y(n2599) );
  INVX1 U234 ( .A(n2588), .Y(n2598) );
  INVX1 U235 ( .A(n2587), .Y(n2601) );
  INVX1 U236 ( .A(n2586), .Y(n2602) );
  INVX1 U237 ( .A(n2586), .Y(n2603) );
  INVX1 U238 ( .A(n2586), .Y(n2604) );
  INVX1 U239 ( .A(n2585), .Y(n2605) );
  INVX1 U240 ( .A(n2585), .Y(n2606) );
  INVX1 U241 ( .A(n2585), .Y(n2607) );
  OR2X1 U242 ( .A(n263), .B(n208), .Y(n206) );
  OR2X1 U243 ( .A(n262), .B(n2678), .Y(n208) );
  OR2X1 U244 ( .A(n263), .B(n211), .Y(n209) );
  OR2X1 U245 ( .A(n6), .B(n11), .Y(n3752) );
  OR2X1 U246 ( .A(n10), .B(n7), .Y(n6) );
  OR2X1 U247 ( .A(n16), .B(n21), .Y(n3785) );
  OR2X1 U248 ( .A(n20), .B(n17), .Y(n16) );
  OR2X1 U249 ( .A(n28), .B(n29), .Y(n27) );
  OR2X1 U250 ( .A(n31), .B(n36), .Y(n3808) );
  OR2X1 U251 ( .A(n35), .B(n32), .Y(n31) );
  OR2X1 U252 ( .A(n41), .B(n46), .Y(n3829) );
  OR2X1 U253 ( .A(n45), .B(n42), .Y(n41) );
  OR2X1 U254 ( .A(n53), .B(n54), .Y(n52) );
  OR2X1 U255 ( .A(n56), .B(n61), .Y(n3852) );
  OR2X1 U256 ( .A(n60), .B(n57), .Y(n56) );
  OR2X1 U257 ( .A(n66), .B(n71), .Y(n3873) );
  OR2X1 U258 ( .A(n70), .B(n67), .Y(n66) );
  OR2X1 U259 ( .A(n78), .B(n79), .Y(n77) );
  OR2X1 U260 ( .A(n81), .B(n86), .Y(n3896) );
  OR2X1 U261 ( .A(n85), .B(n82), .Y(n81) );
  OR2X1 U262 ( .A(n91), .B(n96), .Y(n3917) );
  OR2X1 U263 ( .A(n95), .B(n92), .Y(n91) );
  OR2X1 U264 ( .A(n103), .B(n104), .Y(n102) );
  OR2X1 U265 ( .A(n106), .B(n111), .Y(n3940) );
  OR2X1 U266 ( .A(n110), .B(n107), .Y(n106) );
  OR2X1 U267 ( .A(n116), .B(n121), .Y(n3961) );
  OR2X1 U268 ( .A(n120), .B(n117), .Y(n116) );
  OR2X1 U269 ( .A(n128), .B(n129), .Y(n127) );
  OR2X1 U270 ( .A(n131), .B(n136), .Y(n3984) );
  OR2X1 U271 ( .A(n135), .B(n132), .Y(n131) );
  OR2X1 U272 ( .A(n141), .B(n146), .Y(n4005) );
  OR2X1 U273 ( .A(n145), .B(n142), .Y(n141) );
  OR2X1 U274 ( .A(n153), .B(n154), .Y(n152) );
  OR2X1 U275 ( .A(n156), .B(n161), .Y(n4028) );
  OR2X1 U276 ( .A(n160), .B(n157), .Y(n156) );
  OR2X1 U277 ( .A(n166), .B(n171), .Y(n4049) );
  OR2X1 U278 ( .A(n170), .B(n167), .Y(n166) );
  OR2X1 U279 ( .A(n178), .B(n179), .Y(n177) );
  OR2X1 U280 ( .A(n181), .B(n186), .Y(n4073) );
  OR2X1 U281 ( .A(n185), .B(n182), .Y(n181) );
  OR2X1 U282 ( .A(n191), .B(n196), .Y(n4094) );
  OR2X1 U283 ( .A(n195), .B(n192), .Y(n191) );
  OR2X1 U284 ( .A(n203), .B(n204), .Y(n202) );
  BUFX2 U285 ( .A(n4095), .Y(n2609) );
  INVX1 U286 ( .A(wr), .Y(n3205) );
  INVX1 U287 ( .A(\mem<63><0> ), .Y(n3191) );
  INVX1 U288 ( .A(\mem<63><1> ), .Y(n3190) );
  INVX1 U289 ( .A(\mem<63><2> ), .Y(n3189) );
  INVX1 U290 ( .A(\mem<63><3> ), .Y(n3188) );
  INVX1 U291 ( .A(\mem<63><4> ), .Y(n3187) );
  INVX1 U292 ( .A(\mem<63><5> ), .Y(n3186) );
  INVX1 U293 ( .A(\mem<63><6> ), .Y(n3185) );
  INVX1 U294 ( .A(\mem<63><7> ), .Y(n3184) );
  INVX1 U295 ( .A(\mem<62><0> ), .Y(n3183) );
  INVX1 U296 ( .A(\mem<62><1> ), .Y(n3182) );
  INVX1 U297 ( .A(\mem<62><2> ), .Y(n3181) );
  INVX1 U298 ( .A(\mem<62><3> ), .Y(n3180) );
  INVX1 U299 ( .A(\mem<62><4> ), .Y(n3179) );
  INVX1 U300 ( .A(\mem<62><5> ), .Y(n3178) );
  INVX1 U301 ( .A(\mem<62><6> ), .Y(n3177) );
  INVX1 U302 ( .A(\mem<62><7> ), .Y(n3176) );
  INVX1 U303 ( .A(\mem<61><0> ), .Y(n3175) );
  INVX1 U304 ( .A(\mem<61><1> ), .Y(n3174) );
  INVX1 U305 ( .A(\mem<61><2> ), .Y(n3173) );
  INVX1 U306 ( .A(\mem<61><3> ), .Y(n3172) );
  INVX1 U307 ( .A(\mem<61><4> ), .Y(n3171) );
  INVX1 U308 ( .A(\mem<61><5> ), .Y(n3170) );
  INVX1 U309 ( .A(\mem<61><6> ), .Y(n3169) );
  INVX1 U310 ( .A(\mem<61><7> ), .Y(n3168) );
  INVX1 U311 ( .A(\mem<60><0> ), .Y(n3167) );
  INVX1 U312 ( .A(\mem<60><1> ), .Y(n3166) );
  INVX1 U313 ( .A(\mem<60><2> ), .Y(n3165) );
  INVX1 U314 ( .A(\mem<60><3> ), .Y(n3164) );
  INVX1 U315 ( .A(\mem<60><4> ), .Y(n3163) );
  INVX1 U316 ( .A(\mem<60><5> ), .Y(n3162) );
  INVX1 U317 ( .A(\mem<60><6> ), .Y(n3161) );
  INVX1 U318 ( .A(\mem<60><7> ), .Y(n3160) );
  INVX1 U319 ( .A(\mem<59><0> ), .Y(n3159) );
  INVX1 U320 ( .A(\mem<59><1> ), .Y(n3158) );
  INVX1 U321 ( .A(\mem<59><2> ), .Y(n3157) );
  INVX1 U322 ( .A(\mem<59><3> ), .Y(n3156) );
  INVX1 U323 ( .A(\mem<59><4> ), .Y(n3155) );
  INVX1 U324 ( .A(\mem<59><5> ), .Y(n3154) );
  INVX1 U325 ( .A(\mem<59><6> ), .Y(n3153) );
  INVX1 U326 ( .A(\mem<59><7> ), .Y(n3152) );
  INVX1 U327 ( .A(\mem<58><0> ), .Y(n3151) );
  INVX1 U328 ( .A(\mem<58><1> ), .Y(n3150) );
  INVX1 U329 ( .A(\mem<58><2> ), .Y(n3149) );
  INVX1 U330 ( .A(\mem<58><3> ), .Y(n3148) );
  INVX1 U331 ( .A(\mem<58><4> ), .Y(n3147) );
  INVX1 U332 ( .A(\mem<58><5> ), .Y(n3146) );
  INVX1 U333 ( .A(\mem<58><6> ), .Y(n3145) );
  INVX1 U334 ( .A(\mem<58><7> ), .Y(n3144) );
  INVX1 U335 ( .A(\mem<57><0> ), .Y(n3143) );
  INVX1 U336 ( .A(\mem<57><1> ), .Y(n3142) );
  INVX1 U337 ( .A(\mem<57><2> ), .Y(n3141) );
  INVX1 U338 ( .A(\mem<57><3> ), .Y(n3140) );
  INVX1 U339 ( .A(\mem<57><4> ), .Y(n3139) );
  INVX1 U340 ( .A(\mem<57><5> ), .Y(n3138) );
  INVX1 U341 ( .A(\mem<57><6> ), .Y(n3137) );
  INVX1 U342 ( .A(\mem<57><7> ), .Y(n3136) );
  INVX1 U343 ( .A(\mem<56><0> ), .Y(n3135) );
  INVX1 U344 ( .A(\mem<56><1> ), .Y(n3134) );
  INVX1 U345 ( .A(\mem<56><2> ), .Y(n3133) );
  INVX1 U346 ( .A(\mem<56><3> ), .Y(n3132) );
  INVX1 U347 ( .A(\mem<56><4> ), .Y(n3131) );
  INVX1 U348 ( .A(\mem<56><5> ), .Y(n3130) );
  INVX1 U349 ( .A(\mem<56><6> ), .Y(n3129) );
  INVX1 U350 ( .A(\mem<56><7> ), .Y(n3128) );
  INVX1 U351 ( .A(\mem<55><0> ), .Y(n3127) );
  INVX1 U352 ( .A(\mem<55><1> ), .Y(n3126) );
  INVX1 U353 ( .A(\mem<55><2> ), .Y(n3125) );
  INVX1 U354 ( .A(\mem<55><3> ), .Y(n3124) );
  INVX1 U355 ( .A(\mem<55><4> ), .Y(n3123) );
  INVX1 U356 ( .A(\mem<55><5> ), .Y(n3122) );
  INVX1 U357 ( .A(\mem<55><6> ), .Y(n3121) );
  INVX1 U358 ( .A(\mem<55><7> ), .Y(n3120) );
  INVX1 U359 ( .A(\mem<54><0> ), .Y(n3119) );
  INVX1 U360 ( .A(\mem<54><1> ), .Y(n3118) );
  INVX1 U361 ( .A(\mem<54><2> ), .Y(n3117) );
  INVX1 U362 ( .A(\mem<54><3> ), .Y(n3116) );
  INVX1 U363 ( .A(\mem<54><4> ), .Y(n3115) );
  INVX1 U364 ( .A(\mem<54><5> ), .Y(n3114) );
  INVX1 U365 ( .A(\mem<54><6> ), .Y(n3113) );
  INVX1 U366 ( .A(\mem<54><7> ), .Y(n3112) );
  INVX1 U367 ( .A(\mem<53><0> ), .Y(n3111) );
  INVX1 U368 ( .A(\mem<53><1> ), .Y(n3110) );
  INVX1 U369 ( .A(\mem<53><2> ), .Y(n3109) );
  INVX1 U370 ( .A(\mem<53><3> ), .Y(n3108) );
  INVX1 U371 ( .A(\mem<53><4> ), .Y(n3107) );
  INVX1 U372 ( .A(\mem<53><5> ), .Y(n3106) );
  INVX1 U373 ( .A(\mem<53><6> ), .Y(n3105) );
  INVX1 U374 ( .A(\mem<53><7> ), .Y(n3104) );
  INVX1 U375 ( .A(\mem<52><0> ), .Y(n3103) );
  INVX1 U376 ( .A(\mem<52><1> ), .Y(n3102) );
  INVX1 U377 ( .A(\mem<52><2> ), .Y(n3101) );
  INVX1 U378 ( .A(\mem<52><3> ), .Y(n3100) );
  INVX1 U379 ( .A(\mem<52><4> ), .Y(n3099) );
  INVX1 U380 ( .A(\mem<52><5> ), .Y(n3098) );
  INVX1 U381 ( .A(\mem<52><6> ), .Y(n3097) );
  INVX1 U382 ( .A(\mem<52><7> ), .Y(n3096) );
  INVX1 U383 ( .A(\mem<51><0> ), .Y(n3095) );
  INVX1 U384 ( .A(\mem<51><1> ), .Y(n3094) );
  INVX1 U385 ( .A(\mem<51><2> ), .Y(n3093) );
  INVX1 U386 ( .A(\mem<51><3> ), .Y(n3092) );
  INVX1 U387 ( .A(\mem<51><4> ), .Y(n3091) );
  INVX1 U388 ( .A(\mem<51><5> ), .Y(n3090) );
  INVX1 U389 ( .A(\mem<51><6> ), .Y(n3089) );
  INVX1 U390 ( .A(\mem<51><7> ), .Y(n3088) );
  INVX1 U391 ( .A(\mem<50><0> ), .Y(n3087) );
  INVX1 U392 ( .A(\mem<50><1> ), .Y(n3086) );
  INVX1 U393 ( .A(\mem<50><2> ), .Y(n3085) );
  INVX1 U394 ( .A(\mem<50><3> ), .Y(n3084) );
  INVX1 U395 ( .A(\mem<50><4> ), .Y(n3083) );
  INVX1 U396 ( .A(\mem<50><5> ), .Y(n3082) );
  INVX1 U397 ( .A(\mem<50><6> ), .Y(n3081) );
  INVX1 U398 ( .A(\mem<50><7> ), .Y(n3080) );
  INVX1 U399 ( .A(\mem<49><0> ), .Y(n3079) );
  INVX1 U400 ( .A(\mem<49><1> ), .Y(n3078) );
  INVX1 U401 ( .A(\mem<49><2> ), .Y(n3077) );
  INVX1 U402 ( .A(\mem<49><3> ), .Y(n3076) );
  INVX1 U403 ( .A(\mem<49><4> ), .Y(n3075) );
  INVX1 U404 ( .A(\mem<49><5> ), .Y(n3074) );
  INVX1 U405 ( .A(\mem<49><6> ), .Y(n3073) );
  INVX1 U406 ( .A(\mem<49><7> ), .Y(n3072) );
  INVX1 U407 ( .A(\mem<48><0> ), .Y(n3071) );
  INVX1 U408 ( .A(\mem<48><1> ), .Y(n3070) );
  INVX1 U409 ( .A(\mem<48><2> ), .Y(n3069) );
  INVX1 U410 ( .A(\mem<48><3> ), .Y(n3068) );
  INVX1 U411 ( .A(\mem<48><4> ), .Y(n3067) );
  INVX1 U412 ( .A(\mem<48><5> ), .Y(n3066) );
  INVX1 U413 ( .A(\mem<48><6> ), .Y(n3065) );
  INVX1 U414 ( .A(\mem<48><7> ), .Y(n3064) );
  INVX1 U415 ( .A(\mem<47><0> ), .Y(n3063) );
  INVX1 U416 ( .A(\mem<47><1> ), .Y(n3062) );
  INVX1 U417 ( .A(\mem<47><2> ), .Y(n3061) );
  INVX1 U418 ( .A(\mem<47><3> ), .Y(n3060) );
  INVX1 U419 ( .A(\mem<47><4> ), .Y(n3059) );
  INVX1 U420 ( .A(\mem<47><5> ), .Y(n3058) );
  INVX1 U421 ( .A(\mem<47><6> ), .Y(n3057) );
  INVX1 U422 ( .A(\mem<47><7> ), .Y(n3056) );
  INVX1 U423 ( .A(\mem<46><0> ), .Y(n3055) );
  INVX1 U424 ( .A(\mem<46><1> ), .Y(n3054) );
  INVX1 U425 ( .A(\mem<46><2> ), .Y(n3053) );
  INVX1 U426 ( .A(\mem<46><3> ), .Y(n3052) );
  INVX1 U427 ( .A(\mem<46><4> ), .Y(n3051) );
  INVX1 U428 ( .A(\mem<46><5> ), .Y(n3050) );
  INVX1 U429 ( .A(\mem<46><6> ), .Y(n3049) );
  INVX1 U430 ( .A(\mem<46><7> ), .Y(n3048) );
  INVX1 U431 ( .A(\mem<45><0> ), .Y(n3047) );
  INVX1 U432 ( .A(\mem<45><1> ), .Y(n3046) );
  INVX1 U433 ( .A(\mem<45><2> ), .Y(n3045) );
  INVX1 U434 ( .A(\mem<45><3> ), .Y(n3044) );
  INVX1 U435 ( .A(\mem<45><4> ), .Y(n3043) );
  INVX1 U436 ( .A(\mem<45><5> ), .Y(n3042) );
  INVX1 U437 ( .A(\mem<45><6> ), .Y(n3041) );
  INVX1 U438 ( .A(\mem<45><7> ), .Y(n3040) );
  INVX1 U439 ( .A(\mem<44><0> ), .Y(n3039) );
  INVX1 U440 ( .A(\mem<44><1> ), .Y(n3038) );
  INVX1 U441 ( .A(\mem<44><2> ), .Y(n3037) );
  INVX1 U442 ( .A(\mem<44><3> ), .Y(n3036) );
  INVX1 U443 ( .A(\mem<44><4> ), .Y(n3035) );
  INVX1 U444 ( .A(\mem<44><5> ), .Y(n3034) );
  INVX1 U445 ( .A(\mem<44><6> ), .Y(n3033) );
  INVX1 U446 ( .A(\mem<44><7> ), .Y(n3032) );
  INVX1 U447 ( .A(\mem<43><0> ), .Y(n3031) );
  INVX1 U448 ( .A(\mem<43><1> ), .Y(n3030) );
  INVX1 U449 ( .A(\mem<43><2> ), .Y(n3029) );
  INVX1 U450 ( .A(\mem<43><3> ), .Y(n3028) );
  INVX1 U451 ( .A(\mem<43><4> ), .Y(n3027) );
  INVX1 U452 ( .A(\mem<43><5> ), .Y(n3026) );
  INVX1 U453 ( .A(\mem<43><6> ), .Y(n3025) );
  INVX1 U454 ( .A(\mem<43><7> ), .Y(n3024) );
  INVX1 U455 ( .A(\mem<42><0> ), .Y(n3023) );
  INVX1 U456 ( .A(\mem<42><1> ), .Y(n3022) );
  INVX1 U457 ( .A(\mem<42><2> ), .Y(n3021) );
  INVX1 U458 ( .A(\mem<42><3> ), .Y(n3020) );
  INVX1 U459 ( .A(\mem<42><4> ), .Y(n3019) );
  INVX1 U460 ( .A(\mem<42><5> ), .Y(n3018) );
  INVX1 U461 ( .A(\mem<42><6> ), .Y(n3017) );
  INVX1 U462 ( .A(\mem<42><7> ), .Y(n3016) );
  INVX1 U463 ( .A(\mem<41><0> ), .Y(n3015) );
  INVX1 U464 ( .A(\mem<41><1> ), .Y(n3014) );
  INVX1 U465 ( .A(\mem<41><2> ), .Y(n3013) );
  INVX1 U466 ( .A(\mem<41><3> ), .Y(n3012) );
  INVX1 U467 ( .A(\mem<41><4> ), .Y(n3011) );
  INVX1 U468 ( .A(\mem<41><5> ), .Y(n3010) );
  INVX1 U469 ( .A(\mem<41><6> ), .Y(n3009) );
  INVX1 U470 ( .A(\mem<41><7> ), .Y(n3008) );
  INVX1 U471 ( .A(\mem<40><0> ), .Y(n3007) );
  INVX1 U472 ( .A(\mem<40><1> ), .Y(n3006) );
  INVX1 U473 ( .A(\mem<40><2> ), .Y(n3005) );
  INVX1 U474 ( .A(\mem<40><3> ), .Y(n3004) );
  INVX1 U475 ( .A(\mem<40><4> ), .Y(n3003) );
  INVX1 U476 ( .A(\mem<40><5> ), .Y(n3002) );
  INVX1 U477 ( .A(\mem<40><6> ), .Y(n3001) );
  INVX1 U478 ( .A(\mem<40><7> ), .Y(n3000) );
  INVX1 U479 ( .A(\mem<39><0> ), .Y(n2999) );
  INVX1 U480 ( .A(\mem<39><1> ), .Y(n2998) );
  INVX1 U481 ( .A(\mem<39><2> ), .Y(n2997) );
  INVX1 U482 ( .A(\mem<39><3> ), .Y(n2996) );
  INVX1 U483 ( .A(\mem<39><4> ), .Y(n2995) );
  INVX1 U484 ( .A(\mem<39><5> ), .Y(n2994) );
  INVX1 U485 ( .A(\mem<39><6> ), .Y(n2993) );
  INVX1 U486 ( .A(\mem<39><7> ), .Y(n2992) );
  INVX1 U487 ( .A(\mem<38><0> ), .Y(n2991) );
  INVX1 U488 ( .A(\mem<38><1> ), .Y(n2990) );
  INVX1 U489 ( .A(\mem<38><2> ), .Y(n2989) );
  INVX1 U490 ( .A(\mem<38><3> ), .Y(n2988) );
  INVX1 U491 ( .A(\mem<38><4> ), .Y(n2987) );
  INVX1 U492 ( .A(\mem<38><5> ), .Y(n2986) );
  INVX1 U493 ( .A(\mem<38><6> ), .Y(n2985) );
  INVX1 U494 ( .A(\mem<38><7> ), .Y(n2984) );
  INVX1 U495 ( .A(\mem<37><0> ), .Y(n2983) );
  INVX1 U496 ( .A(\mem<37><1> ), .Y(n2982) );
  INVX1 U497 ( .A(\mem<37><2> ), .Y(n2981) );
  INVX1 U498 ( .A(\mem<37><3> ), .Y(n2980) );
  INVX1 U499 ( .A(\mem<37><4> ), .Y(n2979) );
  INVX1 U500 ( .A(\mem<37><5> ), .Y(n2978) );
  INVX1 U501 ( .A(\mem<37><6> ), .Y(n2977) );
  INVX1 U502 ( .A(\mem<37><7> ), .Y(n2976) );
  INVX1 U503 ( .A(\mem<36><0> ), .Y(n2975) );
  INVX1 U504 ( .A(\mem<36><1> ), .Y(n2974) );
  INVX1 U505 ( .A(\mem<36><2> ), .Y(n2973) );
  INVX1 U506 ( .A(\mem<36><3> ), .Y(n2972) );
  INVX1 U507 ( .A(\mem<36><4> ), .Y(n2971) );
  INVX1 U508 ( .A(\mem<36><5> ), .Y(n2970) );
  INVX1 U509 ( .A(\mem<36><6> ), .Y(n2969) );
  INVX1 U510 ( .A(\mem<36><7> ), .Y(n2968) );
  INVX1 U511 ( .A(\mem<35><0> ), .Y(n2967) );
  INVX1 U512 ( .A(\mem<35><1> ), .Y(n2966) );
  INVX1 U513 ( .A(\mem<35><2> ), .Y(n2965) );
  INVX1 U514 ( .A(\mem<35><3> ), .Y(n2964) );
  INVX1 U515 ( .A(\mem<35><4> ), .Y(n2963) );
  INVX1 U516 ( .A(\mem<35><5> ), .Y(n2962) );
  INVX1 U517 ( .A(\mem<35><6> ), .Y(n2961) );
  INVX1 U518 ( .A(\mem<35><7> ), .Y(n2960) );
  INVX1 U519 ( .A(\mem<34><0> ), .Y(n2959) );
  INVX1 U520 ( .A(\mem<34><1> ), .Y(n2958) );
  INVX1 U521 ( .A(\mem<34><2> ), .Y(n2957) );
  INVX1 U522 ( .A(\mem<34><3> ), .Y(n2956) );
  INVX1 U523 ( .A(\mem<34><4> ), .Y(n2955) );
  INVX1 U524 ( .A(\mem<34><5> ), .Y(n2954) );
  INVX1 U525 ( .A(\mem<34><6> ), .Y(n2953) );
  INVX1 U526 ( .A(\mem<34><7> ), .Y(n2952) );
  INVX1 U527 ( .A(\mem<33><0> ), .Y(n2951) );
  INVX1 U528 ( .A(\mem<33><1> ), .Y(n2950) );
  INVX1 U529 ( .A(\mem<33><2> ), .Y(n2949) );
  INVX1 U530 ( .A(\mem<33><3> ), .Y(n2948) );
  INVX1 U531 ( .A(\mem<33><4> ), .Y(n2947) );
  INVX1 U532 ( .A(\mem<33><5> ), .Y(n2946) );
  INVX1 U533 ( .A(\mem<33><6> ), .Y(n2945) );
  INVX1 U534 ( .A(\mem<33><7> ), .Y(n2944) );
  INVX1 U535 ( .A(\mem<32><0> ), .Y(n2943) );
  INVX1 U536 ( .A(\mem<32><1> ), .Y(n2942) );
  INVX1 U537 ( .A(\mem<32><2> ), .Y(n2941) );
  INVX1 U538 ( .A(\mem<32><3> ), .Y(n2940) );
  INVX1 U539 ( .A(\mem<32><4> ), .Y(n2939) );
  INVX1 U540 ( .A(\mem<32><5> ), .Y(n2938) );
  INVX1 U541 ( .A(\mem<32><6> ), .Y(n2937) );
  INVX1 U542 ( .A(\mem<32><7> ), .Y(n2936) );
  INVX1 U543 ( .A(\mem<31><0> ), .Y(n2935) );
  INVX1 U544 ( .A(\mem<31><1> ), .Y(n2934) );
  INVX1 U545 ( .A(\mem<31><2> ), .Y(n2933) );
  INVX1 U546 ( .A(\mem<31><3> ), .Y(n2932) );
  INVX1 U547 ( .A(\mem<31><4> ), .Y(n2931) );
  INVX1 U548 ( .A(\mem<31><5> ), .Y(n2930) );
  INVX1 U549 ( .A(\mem<31><6> ), .Y(n2929) );
  INVX1 U550 ( .A(\mem<31><7> ), .Y(n2928) );
  INVX1 U551 ( .A(\mem<30><0> ), .Y(n2927) );
  INVX1 U552 ( .A(\mem<30><1> ), .Y(n2926) );
  INVX1 U553 ( .A(\mem<30><2> ), .Y(n2925) );
  INVX1 U554 ( .A(\mem<30><3> ), .Y(n2924) );
  INVX1 U555 ( .A(\mem<30><4> ), .Y(n2923) );
  INVX1 U556 ( .A(\mem<30><5> ), .Y(n2922) );
  INVX1 U557 ( .A(\mem<30><6> ), .Y(n2921) );
  INVX1 U558 ( .A(\mem<30><7> ), .Y(n2920) );
  INVX1 U559 ( .A(\mem<29><0> ), .Y(n2919) );
  INVX1 U560 ( .A(\mem<29><1> ), .Y(n2918) );
  INVX1 U561 ( .A(\mem<29><2> ), .Y(n2917) );
  INVX1 U562 ( .A(\mem<29><3> ), .Y(n2916) );
  INVX1 U563 ( .A(\mem<29><4> ), .Y(n2915) );
  INVX1 U564 ( .A(\mem<29><5> ), .Y(n2914) );
  INVX1 U565 ( .A(\mem<29><6> ), .Y(n2913) );
  INVX1 U566 ( .A(\mem<29><7> ), .Y(n2912) );
  INVX1 U567 ( .A(\mem<28><0> ), .Y(n2911) );
  INVX1 U568 ( .A(\mem<28><1> ), .Y(n2910) );
  INVX1 U569 ( .A(\mem<28><2> ), .Y(n2909) );
  INVX1 U570 ( .A(\mem<28><3> ), .Y(n2908) );
  INVX1 U571 ( .A(\mem<28><4> ), .Y(n2907) );
  INVX1 U572 ( .A(\mem<28><5> ), .Y(n2906) );
  INVX1 U573 ( .A(\mem<28><6> ), .Y(n2905) );
  INVX1 U574 ( .A(\mem<28><7> ), .Y(n2904) );
  INVX1 U575 ( .A(\mem<27><0> ), .Y(n2903) );
  INVX1 U576 ( .A(\mem<27><1> ), .Y(n2902) );
  INVX1 U577 ( .A(\mem<27><2> ), .Y(n2901) );
  INVX1 U578 ( .A(\mem<27><3> ), .Y(n2900) );
  INVX1 U579 ( .A(\mem<27><4> ), .Y(n2899) );
  INVX1 U580 ( .A(\mem<27><5> ), .Y(n2898) );
  INVX1 U581 ( .A(\mem<27><6> ), .Y(n2897) );
  INVX1 U582 ( .A(\mem<27><7> ), .Y(n2896) );
  INVX1 U583 ( .A(\mem<26><0> ), .Y(n2895) );
  INVX1 U584 ( .A(\mem<26><1> ), .Y(n2894) );
  INVX1 U585 ( .A(\mem<26><2> ), .Y(n2893) );
  INVX1 U586 ( .A(\mem<26><3> ), .Y(n2892) );
  INVX1 U587 ( .A(\mem<26><4> ), .Y(n2891) );
  INVX1 U588 ( .A(\mem<26><5> ), .Y(n2890) );
  INVX1 U589 ( .A(\mem<26><6> ), .Y(n2889) );
  INVX1 U590 ( .A(\mem<26><7> ), .Y(n2888) );
  INVX1 U591 ( .A(\mem<25><0> ), .Y(n2887) );
  INVX1 U592 ( .A(\mem<25><1> ), .Y(n2886) );
  INVX1 U593 ( .A(\mem<25><2> ), .Y(n2885) );
  INVX1 U594 ( .A(\mem<25><3> ), .Y(n2884) );
  INVX1 U595 ( .A(\mem<25><4> ), .Y(n2883) );
  INVX1 U596 ( .A(\mem<25><5> ), .Y(n2882) );
  INVX1 U597 ( .A(\mem<25><6> ), .Y(n2881) );
  INVX1 U598 ( .A(\mem<25><7> ), .Y(n2880) );
  INVX1 U599 ( .A(\mem<24><0> ), .Y(n2879) );
  INVX1 U600 ( .A(\mem<24><1> ), .Y(n2878) );
  INVX1 U601 ( .A(\mem<24><2> ), .Y(n2877) );
  INVX1 U602 ( .A(\mem<24><3> ), .Y(n2876) );
  INVX1 U603 ( .A(\mem<24><4> ), .Y(n2875) );
  INVX1 U604 ( .A(\mem<24><5> ), .Y(n2874) );
  INVX1 U605 ( .A(\mem<24><6> ), .Y(n2873) );
  INVX1 U606 ( .A(\mem<24><7> ), .Y(n2872) );
  INVX1 U607 ( .A(\mem<23><0> ), .Y(n2871) );
  INVX1 U608 ( .A(\mem<23><1> ), .Y(n2870) );
  INVX1 U609 ( .A(\mem<23><2> ), .Y(n2869) );
  INVX1 U610 ( .A(\mem<23><3> ), .Y(n2868) );
  INVX1 U611 ( .A(\mem<23><4> ), .Y(n2867) );
  INVX1 U612 ( .A(\mem<23><5> ), .Y(n2866) );
  INVX1 U613 ( .A(\mem<23><6> ), .Y(n2865) );
  INVX1 U614 ( .A(\mem<23><7> ), .Y(n2864) );
  INVX1 U615 ( .A(\mem<22><0> ), .Y(n2863) );
  INVX1 U616 ( .A(\mem<22><1> ), .Y(n2862) );
  INVX1 U617 ( .A(\mem<22><2> ), .Y(n2861) );
  INVX1 U618 ( .A(\mem<22><3> ), .Y(n2860) );
  INVX1 U619 ( .A(\mem<22><4> ), .Y(n2859) );
  INVX1 U620 ( .A(\mem<22><5> ), .Y(n2858) );
  INVX1 U621 ( .A(\mem<22><6> ), .Y(n2857) );
  INVX1 U622 ( .A(\mem<22><7> ), .Y(n2856) );
  INVX1 U623 ( .A(\mem<21><0> ), .Y(n2855) );
  INVX1 U624 ( .A(\mem<21><1> ), .Y(n2854) );
  INVX1 U625 ( .A(\mem<21><2> ), .Y(n2853) );
  INVX1 U626 ( .A(\mem<21><3> ), .Y(n2852) );
  INVX1 U627 ( .A(\mem<21><4> ), .Y(n2851) );
  INVX1 U628 ( .A(\mem<21><5> ), .Y(n2850) );
  INVX1 U629 ( .A(\mem<21><6> ), .Y(n2849) );
  INVX1 U630 ( .A(\mem<21><7> ), .Y(n2848) );
  INVX1 U631 ( .A(\mem<20><0> ), .Y(n2847) );
  INVX1 U632 ( .A(\mem<20><1> ), .Y(n2846) );
  INVX1 U633 ( .A(\mem<20><2> ), .Y(n2845) );
  INVX1 U634 ( .A(\mem<20><3> ), .Y(n2844) );
  INVX1 U635 ( .A(\mem<20><4> ), .Y(n2843) );
  INVX1 U636 ( .A(\mem<20><5> ), .Y(n2842) );
  INVX1 U637 ( .A(\mem<20><6> ), .Y(n2841) );
  INVX1 U638 ( .A(\mem<20><7> ), .Y(n2840) );
  INVX1 U639 ( .A(\mem<19><0> ), .Y(n2839) );
  INVX1 U640 ( .A(\mem<19><1> ), .Y(n2838) );
  INVX1 U641 ( .A(\mem<19><2> ), .Y(n2837) );
  INVX1 U642 ( .A(\mem<19><3> ), .Y(n2836) );
  INVX1 U643 ( .A(\mem<19><4> ), .Y(n2835) );
  INVX1 U644 ( .A(\mem<19><5> ), .Y(n2834) );
  INVX1 U645 ( .A(\mem<19><6> ), .Y(n2833) );
  INVX1 U646 ( .A(\mem<19><7> ), .Y(n2832) );
  INVX1 U647 ( .A(\mem<18><0> ), .Y(n2831) );
  INVX1 U648 ( .A(\mem<18><1> ), .Y(n2830) );
  INVX1 U649 ( .A(\mem<18><2> ), .Y(n2829) );
  INVX1 U650 ( .A(\mem<18><3> ), .Y(n2828) );
  INVX1 U651 ( .A(\mem<18><4> ), .Y(n2827) );
  INVX1 U652 ( .A(\mem<18><5> ), .Y(n2826) );
  INVX1 U653 ( .A(\mem<18><6> ), .Y(n2825) );
  INVX1 U654 ( .A(\mem<18><7> ), .Y(n2824) );
  INVX1 U655 ( .A(\mem<17><0> ), .Y(n2823) );
  INVX1 U656 ( .A(\mem<17><1> ), .Y(n2822) );
  INVX1 U657 ( .A(\mem<17><2> ), .Y(n2821) );
  INVX1 U658 ( .A(\mem<17><3> ), .Y(n2820) );
  INVX1 U659 ( .A(\mem<17><4> ), .Y(n2819) );
  INVX1 U660 ( .A(\mem<17><5> ), .Y(n2818) );
  INVX1 U661 ( .A(\mem<17><6> ), .Y(n2817) );
  INVX1 U662 ( .A(\mem<17><7> ), .Y(n2816) );
  INVX1 U663 ( .A(\mem<16><0> ), .Y(n2815) );
  INVX1 U664 ( .A(\mem<16><1> ), .Y(n2814) );
  INVX1 U665 ( .A(\mem<16><2> ), .Y(n2813) );
  INVX1 U666 ( .A(\mem<16><3> ), .Y(n2812) );
  INVX1 U667 ( .A(\mem<16><4> ), .Y(n2811) );
  INVX1 U668 ( .A(\mem<16><5> ), .Y(n2810) );
  INVX1 U669 ( .A(\mem<16><6> ), .Y(n2809) );
  INVX1 U670 ( .A(\mem<16><7> ), .Y(n2808) );
  INVX1 U671 ( .A(\mem<15><0> ), .Y(n2807) );
  INVX1 U672 ( .A(\mem<15><1> ), .Y(n2806) );
  INVX1 U673 ( .A(\mem<15><2> ), .Y(n2805) );
  INVX1 U674 ( .A(\mem<15><3> ), .Y(n2804) );
  INVX1 U675 ( .A(\mem<15><4> ), .Y(n2803) );
  INVX1 U676 ( .A(\mem<15><5> ), .Y(n2802) );
  INVX1 U677 ( .A(\mem<15><6> ), .Y(n2801) );
  INVX1 U678 ( .A(\mem<15><7> ), .Y(n2800) );
  INVX1 U679 ( .A(\mem<14><0> ), .Y(n2799) );
  INVX1 U680 ( .A(\mem<14><1> ), .Y(n2798) );
  INVX1 U681 ( .A(\mem<14><2> ), .Y(n2797) );
  INVX1 U682 ( .A(\mem<14><3> ), .Y(n2796) );
  INVX1 U683 ( .A(\mem<14><4> ), .Y(n2795) );
  INVX1 U684 ( .A(\mem<14><5> ), .Y(n2794) );
  INVX1 U685 ( .A(\mem<14><6> ), .Y(n2793) );
  INVX1 U686 ( .A(\mem<14><7> ), .Y(n2792) );
  INVX1 U687 ( .A(\mem<13><0> ), .Y(n2791) );
  INVX1 U688 ( .A(\mem<13><1> ), .Y(n2790) );
  INVX1 U689 ( .A(\mem<13><2> ), .Y(n2789) );
  INVX1 U690 ( .A(\mem<13><3> ), .Y(n2788) );
  INVX1 U691 ( .A(\mem<13><4> ), .Y(n2787) );
  INVX1 U692 ( .A(\mem<13><5> ), .Y(n2786) );
  INVX1 U693 ( .A(\mem<13><6> ), .Y(n2785) );
  INVX1 U694 ( .A(\mem<13><7> ), .Y(n2784) );
  INVX1 U695 ( .A(\mem<12><0> ), .Y(n2783) );
  INVX1 U696 ( .A(\mem<12><1> ), .Y(n2782) );
  INVX1 U697 ( .A(\mem<12><2> ), .Y(n2781) );
  INVX1 U698 ( .A(\mem<12><3> ), .Y(n2780) );
  INVX1 U699 ( .A(\mem<12><4> ), .Y(n2779) );
  INVX1 U700 ( .A(\mem<12><5> ), .Y(n2778) );
  INVX1 U701 ( .A(\mem<12><6> ), .Y(n2777) );
  INVX1 U702 ( .A(\mem<12><7> ), .Y(n2776) );
  INVX1 U703 ( .A(\mem<11><0> ), .Y(n2775) );
  INVX1 U704 ( .A(\mem<11><1> ), .Y(n2774) );
  INVX1 U705 ( .A(\mem<11><2> ), .Y(n2773) );
  INVX1 U706 ( .A(\mem<11><3> ), .Y(n2772) );
  INVX1 U707 ( .A(\mem<11><4> ), .Y(n2771) );
  INVX1 U708 ( .A(\mem<11><5> ), .Y(n2770) );
  INVX1 U709 ( .A(\mem<11><6> ), .Y(n2769) );
  INVX1 U710 ( .A(\mem<11><7> ), .Y(n2768) );
  INVX1 U711 ( .A(\mem<10><0> ), .Y(n2767) );
  INVX1 U712 ( .A(\mem<10><1> ), .Y(n2766) );
  INVX1 U713 ( .A(\mem<10><2> ), .Y(n2765) );
  INVX1 U714 ( .A(\mem<10><3> ), .Y(n2764) );
  INVX1 U715 ( .A(\mem<10><4> ), .Y(n2763) );
  INVX1 U716 ( .A(\mem<10><5> ), .Y(n2762) );
  INVX1 U717 ( .A(\mem<10><6> ), .Y(n2761) );
  INVX1 U718 ( .A(\mem<10><7> ), .Y(n2760) );
  INVX1 U719 ( .A(\mem<9><0> ), .Y(n2759) );
  INVX1 U720 ( .A(\mem<9><1> ), .Y(n2758) );
  INVX1 U721 ( .A(\mem<9><2> ), .Y(n2757) );
  INVX1 U722 ( .A(\mem<9><3> ), .Y(n2756) );
  INVX1 U723 ( .A(\mem<9><4> ), .Y(n2755) );
  INVX1 U724 ( .A(\mem<9><5> ), .Y(n2754) );
  INVX1 U725 ( .A(\mem<9><6> ), .Y(n2753) );
  INVX1 U726 ( .A(\mem<9><7> ), .Y(n2752) );
  INVX1 U727 ( .A(\mem<8><0> ), .Y(n2751) );
  INVX1 U728 ( .A(\mem<8><1> ), .Y(n2750) );
  INVX1 U729 ( .A(\mem<8><2> ), .Y(n2749) );
  INVX1 U730 ( .A(\mem<8><3> ), .Y(n2748) );
  INVX1 U731 ( .A(\mem<8><4> ), .Y(n2747) );
  INVX1 U732 ( .A(\mem<8><5> ), .Y(n2746) );
  INVX1 U733 ( .A(\mem<8><6> ), .Y(n2745) );
  INVX1 U734 ( .A(\mem<8><7> ), .Y(n2744) );
  INVX1 U735 ( .A(\mem<7><0> ), .Y(n2743) );
  INVX1 U736 ( .A(\mem<7><1> ), .Y(n2742) );
  INVX1 U737 ( .A(\mem<7><2> ), .Y(n2741) );
  INVX1 U738 ( .A(\mem<7><3> ), .Y(n2740) );
  INVX1 U739 ( .A(\mem<7><4> ), .Y(n2739) );
  INVX1 U740 ( .A(\mem<7><5> ), .Y(n2738) );
  INVX1 U741 ( .A(\mem<7><6> ), .Y(n2737) );
  INVX1 U742 ( .A(\mem<7><7> ), .Y(n2736) );
  INVX1 U743 ( .A(\mem<6><0> ), .Y(n2735) );
  INVX1 U744 ( .A(\mem<6><1> ), .Y(n2734) );
  INVX1 U745 ( .A(\mem<6><2> ), .Y(n2733) );
  INVX1 U746 ( .A(\mem<6><3> ), .Y(n2732) );
  INVX1 U747 ( .A(\mem<6><4> ), .Y(n2731) );
  INVX1 U748 ( .A(\mem<6><5> ), .Y(n2730) );
  INVX1 U749 ( .A(\mem<6><6> ), .Y(n2729) );
  INVX1 U750 ( .A(\mem<6><7> ), .Y(n2728) );
  INVX1 U751 ( .A(\mem<5><0> ), .Y(n2727) );
  INVX1 U752 ( .A(\mem<5><1> ), .Y(n2726) );
  INVX1 U753 ( .A(\mem<5><2> ), .Y(n2725) );
  INVX1 U754 ( .A(\mem<5><3> ), .Y(n2724) );
  INVX1 U755 ( .A(\mem<5><4> ), .Y(n2723) );
  INVX1 U756 ( .A(\mem<5><5> ), .Y(n2722) );
  INVX1 U757 ( .A(\mem<5><6> ), .Y(n2721) );
  INVX1 U758 ( .A(\mem<5><7> ), .Y(n2720) );
  INVX1 U759 ( .A(\mem<4><0> ), .Y(n2719) );
  INVX1 U760 ( .A(\mem<4><1> ), .Y(n2718) );
  INVX1 U761 ( .A(\mem<4><2> ), .Y(n2717) );
  INVX1 U762 ( .A(\mem<4><3> ), .Y(n2716) );
  INVX1 U763 ( .A(\mem<4><4> ), .Y(n2715) );
  INVX1 U764 ( .A(\mem<4><5> ), .Y(n2714) );
  INVX1 U765 ( .A(\mem<4><6> ), .Y(n2713) );
  INVX1 U766 ( .A(\mem<4><7> ), .Y(n2712) );
  INVX1 U767 ( .A(\mem<3><0> ), .Y(n2711) );
  INVX1 U768 ( .A(\mem<3><1> ), .Y(n2710) );
  INVX1 U769 ( .A(\mem<3><2> ), .Y(n2709) );
  INVX1 U770 ( .A(\mem<3><3> ), .Y(n2708) );
  INVX1 U771 ( .A(\mem<3><4> ), .Y(n2707) );
  INVX1 U772 ( .A(\mem<3><5> ), .Y(n2706) );
  INVX1 U773 ( .A(\mem<3><6> ), .Y(n2705) );
  INVX1 U774 ( .A(\mem<3><7> ), .Y(n2704) );
  INVX1 U775 ( .A(\mem<2><0> ), .Y(n2703) );
  INVX1 U776 ( .A(\mem<2><1> ), .Y(n2702) );
  INVX1 U777 ( .A(\mem<2><2> ), .Y(n2701) );
  INVX1 U778 ( .A(\mem<2><3> ), .Y(n2700) );
  INVX1 U779 ( .A(\mem<2><4> ), .Y(n2699) );
  INVX1 U780 ( .A(\mem<2><5> ), .Y(n2698) );
  INVX1 U781 ( .A(\mem<2><6> ), .Y(n2697) );
  INVX1 U782 ( .A(\mem<2><7> ), .Y(n2696) );
  INVX1 U783 ( .A(\mem<1><0> ), .Y(n2695) );
  INVX1 U784 ( .A(\mem<1><1> ), .Y(n2694) );
  INVX1 U785 ( .A(\mem<1><2> ), .Y(n2693) );
  INVX1 U786 ( .A(\mem<1><3> ), .Y(n2692) );
  INVX1 U787 ( .A(\mem<1><4> ), .Y(n2691) );
  INVX1 U788 ( .A(\mem<1><5> ), .Y(n2690) );
  INVX1 U789 ( .A(\mem<1><6> ), .Y(n2689) );
  INVX1 U790 ( .A(\mem<1><7> ), .Y(n2688) );
  INVX1 U791 ( .A(\mem<0><0> ), .Y(n2687) );
  INVX1 U792 ( .A(\mem<0><1> ), .Y(n2686) );
  INVX1 U793 ( .A(\mem<0><2> ), .Y(n2685) );
  INVX1 U794 ( .A(\mem<0><3> ), .Y(n2684) );
  INVX1 U795 ( .A(\mem<0><4> ), .Y(n2683) );
  INVX1 U796 ( .A(\mem<0><5> ), .Y(n2682) );
  INVX1 U797 ( .A(\mem<0><6> ), .Y(n2681) );
  INVX1 U798 ( .A(\mem<0><7> ), .Y(n2680) );
  INVX1 U799 ( .A(n2589), .Y(n2590) );
  INVX1 U800 ( .A(n2676), .Y(n2581) );
  INVX1 U801 ( .A(n2676), .Y(n2580) );
  INVX1 U802 ( .A(n2589), .Y(n2592) );
  INVX1 U803 ( .A(n2675), .Y(n2593) );
  INVX1 U804 ( .A(n2675), .Y(n2591) );
  INVX1 U805 ( .A(n2676), .Y(n2584) );
  INVX1 U806 ( .A(n2676), .Y(n2583) );
  INVX1 U807 ( .A(n2676), .Y(n2582) );
  INVX1 U808 ( .A(n2675), .Y(n2595) );
  INVX1 U809 ( .A(n2675), .Y(n2594) );
  INVX1 U810 ( .A(N179), .Y(n2677) );
  INVX1 U811 ( .A(N178), .Y(n2676) );
  INVX1 U812 ( .A(n2677), .Y(n2576) );
  INVX1 U813 ( .A(n2677), .Y(n2577) );
  INVX1 U814 ( .A(n2676), .Y(n2578) );
  INVX1 U815 ( .A(n2676), .Y(n2579) );
  INVX1 U816 ( .A(n2678), .Y(n2574) );
  INVX1 U1904 ( .A(n2678), .Y(n2573) );
  OR2X1 U1908 ( .A(n264), .B(N180), .Y(n211) );
  INVX1 U1913 ( .A(N177), .Y(n2675) );
  OR2X1 U1918 ( .A(n279), .B(n213), .Y(n212) );
  OR2X1 U1923 ( .A(n30), .B(n27), .Y(n26) );
  OR2X1 U1929 ( .A(n282), .B(n215), .Y(n214) );
  OR2X1 U1934 ( .A(n55), .B(n52), .Y(n51) );
  OR2X1 U1939 ( .A(n285), .B(n217), .Y(n216) );
  OR2X1 U1944 ( .A(n80), .B(n77), .Y(n76) );
  OR2X1 U1951 ( .A(n288), .B(n219), .Y(n218) );
  OR2X1 U1956 ( .A(n105), .B(n102), .Y(n101) );
  OR2X1 U1961 ( .A(n291), .B(n221), .Y(n220) );
  OR2X1 U1966 ( .A(n130), .B(n127), .Y(n126) );
  OR2X1 U1972 ( .A(n294), .B(n223), .Y(n222) );
  OR2X1 U1977 ( .A(n155), .B(n152), .Y(n151) );
  OR2X1 U1982 ( .A(n297), .B(n225), .Y(n224) );
  OR2X1 U1987 ( .A(n180), .B(n177), .Y(n176) );
  OR2X1 U1994 ( .A(n300), .B(n227), .Y(n226) );
  OR2X1 U1999 ( .A(n205), .B(n202), .Y(n201) );
  OR2X1 U2004 ( .A(n5), .B(n2), .Y(n1) );
  OR2X1 U2009 ( .A(n8), .B(n9), .Y(n7) );
  OR2X1 U2015 ( .A(n18), .B(n19), .Y(n17) );
  OR2X1 U2020 ( .A(n33), .B(n34), .Y(n32) );
  OR2X1 U2025 ( .A(n43), .B(n44), .Y(n42) );
  OR2X1 U2030 ( .A(n58), .B(n59), .Y(n57) );
  OR2X1 U2037 ( .A(n68), .B(n69), .Y(n67) );
  OR2X1 U2042 ( .A(n83), .B(n84), .Y(n82) );
  OR2X1 U2047 ( .A(n93), .B(n94), .Y(n92) );
  OR2X1 U2052 ( .A(n108), .B(n109), .Y(n107) );
  OR2X1 U2058 ( .A(n118), .B(n119), .Y(n117) );
  OR2X1 U2063 ( .A(n133), .B(n134), .Y(n132) );
  OR2X1 U2068 ( .A(n143), .B(n144), .Y(n142) );
  OR2X1 U2073 ( .A(n158), .B(n159), .Y(n157) );
  OR2X1 U2080 ( .A(n168), .B(n169), .Y(n167) );
  OR2X1 U2085 ( .A(n183), .B(n184), .Y(n182) );
  OR2X1 U2090 ( .A(n193), .B(n194), .Y(n192) );
  OR2X1 U2095 ( .A(n15), .B(n12), .Y(n11) );
  OR2X1 U2101 ( .A(n25), .B(n22), .Y(n21) );
  OR2X1 U2106 ( .A(n40), .B(n37), .Y(n36) );
  OR2X1 U2111 ( .A(n50), .B(n47), .Y(n46) );
  OR2X1 U2116 ( .A(n65), .B(n62), .Y(n61) );
  OR2X1 U2123 ( .A(n75), .B(n72), .Y(n71) );
  OR2X1 U2128 ( .A(n90), .B(n87), .Y(n86) );
  OR2X1 U2133 ( .A(n100), .B(n97), .Y(n96) );
  OR2X1 U2138 ( .A(n115), .B(n112), .Y(n111) );
  OR2X1 U2144 ( .A(n125), .B(n122), .Y(n121) );
  OR2X1 U2149 ( .A(n140), .B(n137), .Y(n136) );
  OR2X1 U2154 ( .A(n150), .B(n147), .Y(n146) );
  OR2X1 U2159 ( .A(n165), .B(n162), .Y(n161) );
  OR2X1 U2166 ( .A(n175), .B(n172), .Y(n171) );
  OR2X1 U2171 ( .A(n190), .B(n187), .Y(n186) );
  OR2X1 U2176 ( .A(n200), .B(n197), .Y(n196) );
  INVX1 U2181 ( .A(n2675), .Y(n2608) );
  INVX1 U2187 ( .A(n2674), .Y(n2673) );
  INVX1 U2192 ( .A(n2674), .Y(n2672) );
  INVX1 U2197 ( .A(N181), .Y(n2571) );
  INVX1 U2202 ( .A(n2571), .Y(n2572) );
  INVX1 U2210 ( .A(n2677), .Y(n2575) );
  INVX1 U2212 ( .A(N177), .Y(n2589) );
  OR2X1 U2213 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U2215 ( .A(n3195), .Y(n3) );
  INVX1 U2216 ( .A(n3200), .Y(n4) );
  INVX1 U2218 ( .A(\addr<10> ), .Y(n5) );
  INVX1 U2219 ( .A(n4789), .Y(n3195) );
  INVX1 U2221 ( .A(n3728), .Y(n8) );
  INVX1 U2222 ( .A(n3729), .Y(n9) );
  INVX1 U2223 ( .A(n3730), .Y(n10) );
  INVX1 U2225 ( .A(n3733), .Y(n13) );
  INVX1 U2226 ( .A(n3734), .Y(n14) );
  INVX1 U2228 ( .A(n3735), .Y(n15) );
  INVX1 U2229 ( .A(n3757), .Y(n18) );
  INVX1 U2231 ( .A(n3758), .Y(n19) );
  INVX1 U2232 ( .A(n3759), .Y(n20) );
  INVX1 U2234 ( .A(n3762), .Y(n23) );
  INVX1 U2236 ( .A(n3763), .Y(n24) );
  INVX1 U2237 ( .A(n3764), .Y(n25) );
  INVX1 U2238 ( .A(n3770), .Y(n28) );
  INVX1 U2240 ( .A(n3771), .Y(n29) );
  INVX1 U2241 ( .A(n3772), .Y(n30) );
  INVX1 U2243 ( .A(n3790), .Y(n33) );
  INVX1 U2244 ( .A(n3791), .Y(n34) );
  INVX1 U2246 ( .A(n3792), .Y(n35) );
  INVX1 U2247 ( .A(n3795), .Y(n38) );
  INVX1 U2249 ( .A(n3796), .Y(n39) );
  INVX1 U2250 ( .A(n3797), .Y(n40) );
  INVX1 U2251 ( .A(n3811), .Y(n43) );
  INVX1 U2253 ( .A(n3812), .Y(n44) );
  INVX1 U2254 ( .A(n3813), .Y(n45) );
  INVX1 U2256 ( .A(n3816), .Y(n48) );
  INVX1 U2257 ( .A(n3817), .Y(n49) );
  INVX1 U2259 ( .A(n3818), .Y(n50) );
  INVX1 U2260 ( .A(n3821), .Y(n53) );
  INVX1 U2262 ( .A(n3822), .Y(n54) );
  INVX1 U2264 ( .A(n3823), .Y(n55) );
  INVX1 U2265 ( .A(n3834), .Y(n58) );
  INVX1 U2267 ( .A(n3835), .Y(n59) );
  INVX1 U2269 ( .A(n3836), .Y(n60) );
  INVX1 U2271 ( .A(n3839), .Y(n63) );
  INVX1 U2272 ( .A(n3840), .Y(n64) );
  INVX1 U2274 ( .A(n3841), .Y(n65) );
  INVX1 U2275 ( .A(n3855), .Y(n68) );
  INVX1 U2277 ( .A(n3856), .Y(n69) );
  INVX1 U2278 ( .A(n3857), .Y(n70) );
  INVX1 U2283 ( .A(n3860), .Y(n73) );
  INVX1 U2286 ( .A(n3861), .Y(n74) );
  INVX1 U2287 ( .A(n3862), .Y(n75) );
  INVX1 U2289 ( .A(n3865), .Y(n78) );
  INVX1 U2290 ( .A(n3866), .Y(n79) );
  INVX1 U2292 ( .A(n3867), .Y(n80) );
  INVX1 U2293 ( .A(n3878), .Y(n83) );
  INVX1 U2295 ( .A(n3879), .Y(n84) );
  INVX1 U2296 ( .A(n3880), .Y(n85) );
  INVX1 U2298 ( .A(n3883), .Y(n88) );
  INVX1 U2299 ( .A(n3884), .Y(n89) );
  INVX1 U2300 ( .A(n3885), .Y(n90) );
  INVX1 U2301 ( .A(n3899), .Y(n93) );
  INVX1 U2303 ( .A(n3900), .Y(n94) );
  INVX1 U2304 ( .A(n3901), .Y(n95) );
  INVX1 U2306 ( .A(n3904), .Y(n98) );
  INVX1 U2307 ( .A(n3905), .Y(n99) );
  INVX1 U2309 ( .A(n3906), .Y(n100) );
  INVX1 U2310 ( .A(n3909), .Y(n103) );
  INVX1 U2312 ( .A(n3910), .Y(n104) );
  INVX1 U2313 ( .A(n3911), .Y(n105) );
  INVX1 U2315 ( .A(n3922), .Y(n108) );
  INVX1 U2316 ( .A(n3923), .Y(n109) );
  INVX1 U2318 ( .A(n3924), .Y(n110) );
  INVX1 U2320 ( .A(n3927), .Y(n113) );
  INVX1 U2323 ( .A(n3928), .Y(n114) );
  INVX1 U2325 ( .A(n3929), .Y(n115) );
  INVX1 U2328 ( .A(n3943), .Y(n118) );
  INVX1 U2330 ( .A(n3944), .Y(n119) );
  INVX1 U2333 ( .A(n3945), .Y(n120) );
  INVX1 U2337 ( .A(n3948), .Y(n123) );
  INVX1 U2345 ( .A(n3949), .Y(n124) );
  INVX1 U2346 ( .A(n3950), .Y(n125) );
  INVX1 U2347 ( .A(n3953), .Y(n128) );
  INVX1 U2348 ( .A(n3954), .Y(n129) );
  INVX1 U2349 ( .A(n3955), .Y(n130) );
  INVX1 U2350 ( .A(n3966), .Y(n133) );
  INVX1 U2351 ( .A(n3967), .Y(n134) );
  INVX1 U2352 ( .A(n3968), .Y(n135) );
  INVX1 U2353 ( .A(n3971), .Y(n138) );
  INVX1 U2354 ( .A(n3972), .Y(n139) );
  INVX1 U2355 ( .A(n3973), .Y(n140) );
  INVX1 U2356 ( .A(n3987), .Y(n143) );
  INVX1 U2357 ( .A(n3988), .Y(n144) );
  INVX1 U2358 ( .A(n3989), .Y(n145) );
  INVX1 U2359 ( .A(n3992), .Y(n148) );
  INVX1 U2360 ( .A(n3993), .Y(n149) );
  INVX1 U2361 ( .A(n3994), .Y(n150) );
  INVX1 U2362 ( .A(n3997), .Y(n153) );
  INVX1 U2363 ( .A(n3998), .Y(n154) );
  INVX1 U2364 ( .A(n3999), .Y(n155) );
  INVX1 U2365 ( .A(n4010), .Y(n158) );
  INVX1 U2366 ( .A(n4011), .Y(n159) );
  INVX1 U2367 ( .A(n4012), .Y(n160) );
  INVX1 U2368 ( .A(n4015), .Y(n163) );
  INVX1 U2369 ( .A(n4016), .Y(n164) );
  INVX1 U2370 ( .A(n4017), .Y(n165) );
  INVX1 U2371 ( .A(n4031), .Y(n168) );
  INVX1 U2372 ( .A(n4032), .Y(n169) );
  INVX1 U2373 ( .A(n4033), .Y(n170) );
  INVX1 U2374 ( .A(n4036), .Y(n173) );
  INVX1 U2375 ( .A(n4037), .Y(n174) );
  INVX1 U2376 ( .A(n4038), .Y(n175) );
  INVX1 U2377 ( .A(n4041), .Y(n178) );
  INVX1 U2378 ( .A(n4042), .Y(n179) );
  INVX1 U2379 ( .A(n4043), .Y(n180) );
  INVX1 U2380 ( .A(n4054), .Y(n183) );
  INVX1 U2381 ( .A(n4055), .Y(n184) );
  INVX1 U2382 ( .A(n4056), .Y(n185) );
  INVX1 U2383 ( .A(n4059), .Y(n188) );
  INVX1 U2384 ( .A(n4060), .Y(n189) );
  INVX1 U2385 ( .A(n4061), .Y(n190) );
  INVX1 U2386 ( .A(n4076), .Y(n193) );
  INVX1 U2387 ( .A(n4077), .Y(n194) );
  INVX1 U2388 ( .A(n4078), .Y(n195) );
  INVX1 U2389 ( .A(n4081), .Y(n198) );
  INVX1 U2390 ( .A(n4082), .Y(n199) );
  INVX1 U2391 ( .A(n4083), .Y(n200) );
  INVX1 U2392 ( .A(n4086), .Y(n203) );
  INVX1 U2393 ( .A(n4087), .Y(n204) );
  INVX1 U2394 ( .A(n4088), .Y(n205) );
  INVX1 U2395 ( .A(n206), .Y(n207) );
  INVX1 U2396 ( .A(n209), .Y(n210) );
  OR2X1 U2397 ( .A(n277), .B(n278), .Y(n213) );
  OR2X1 U2398 ( .A(n280), .B(n281), .Y(n215) );
  OR2X1 U2399 ( .A(n283), .B(n284), .Y(n217) );
  OR2X1 U2400 ( .A(n286), .B(n287), .Y(n219) );
  OR2X1 U2401 ( .A(n289), .B(n290), .Y(n221) );
  OR2X1 U2402 ( .A(n292), .B(n293), .Y(n223) );
  OR2X1 U2403 ( .A(n295), .B(n296), .Y(n225) );
  OR2X1 U2404 ( .A(n298), .B(n299), .Y(n227) );
  OR2X1 U2405 ( .A(n303), .B(n229), .Y(n228) );
  OR2X1 U2406 ( .A(n301), .B(n302), .Y(n229) );
  OR2X1 U2407 ( .A(n306), .B(n231), .Y(n230) );
  OR2X1 U2408 ( .A(n304), .B(n305), .Y(n231) );
  OR2X1 U2409 ( .A(n309), .B(n233), .Y(n232) );
  OR2X1 U2410 ( .A(n307), .B(n308), .Y(n233) );
  OR2X1 U2411 ( .A(n312), .B(n235), .Y(n234) );
  OR2X1 U2412 ( .A(n310), .B(n311), .Y(n235) );
  OR2X1 U2413 ( .A(n315), .B(n237), .Y(n236) );
  OR2X1 U2414 ( .A(n313), .B(n314), .Y(n237) );
  OR2X1 U2415 ( .A(n318), .B(n239), .Y(n238) );
  OR2X1 U2416 ( .A(n316), .B(n317), .Y(n239) );
  OR2X1 U2417 ( .A(n321), .B(n241), .Y(n240) );
  OR2X1 U2418 ( .A(n319), .B(n320), .Y(n241) );
  OR2X1 U2419 ( .A(n324), .B(n243), .Y(n242) );
  OR2X1 U2420 ( .A(n322), .B(n323), .Y(n243) );
  OR2X1 U2421 ( .A(n327), .B(n245), .Y(n244) );
  OR2X1 U2422 ( .A(n325), .B(n326), .Y(n245) );
  OR2X1 U2423 ( .A(n330), .B(n247), .Y(n246) );
  OR2X1 U2424 ( .A(n328), .B(n329), .Y(n247) );
  OR2X1 U2425 ( .A(n333), .B(n249), .Y(n248) );
  OR2X1 U2426 ( .A(n331), .B(n332), .Y(n249) );
  OR2X1 U2427 ( .A(n336), .B(n251), .Y(n250) );
  OR2X1 U2428 ( .A(n334), .B(n335), .Y(n251) );
  OR2X1 U2429 ( .A(n339), .B(n253), .Y(n252) );
  OR2X1 U2430 ( .A(n337), .B(n338), .Y(n253) );
  OR2X1 U2431 ( .A(n342), .B(n255), .Y(n254) );
  OR2X1 U2432 ( .A(n340), .B(n341), .Y(n255) );
  OR2X1 U2433 ( .A(n345), .B(n257), .Y(n256) );
  OR2X1 U2434 ( .A(n343), .B(n344), .Y(n257) );
  OR2X1 U2435 ( .A(n348), .B(n259), .Y(n258) );
  OR2X1 U2436 ( .A(n346), .B(n347), .Y(n259) );
  BUFX2 U2437 ( .A(n3723), .Y(n260) );
  INVX1 U2438 ( .A(n260), .Y(n3196) );
  BUFX2 U2439 ( .A(n3725), .Y(n261) );
  INVX1 U2440 ( .A(n261), .Y(n3201) );
  INVX1 U2441 ( .A(n3736), .Y(n262) );
  INVX1 U2442 ( .A(n3766), .Y(n263) );
  INVX1 U2443 ( .A(n3736), .Y(n264) );
  INVX1 U2444 ( .A(N180), .Y(n2678) );
  INVX1 U2445 ( .A(n3753), .Y(n3197) );
  INVX1 U2446 ( .A(n3754), .Y(n3199) );
  INVX1 U2447 ( .A(n3767), .Y(n3198) );
  AND2X1 U2448 ( .A(n3721), .B(n3720), .Y(n3766) );
  AND2X1 U2449 ( .A(n2678), .B(N181), .Y(n3765) );
  BUFX2 U2450 ( .A(n4809), .Y(\data_out<0> ) );
  BUFX2 U2451 ( .A(n4808), .Y(\data_out<1> ) );
  BUFX2 U2452 ( .A(n4807), .Y(\data_out<2> ) );
  BUFX2 U2453 ( .A(n4806), .Y(\data_out<3> ) );
  BUFX2 U2454 ( .A(n4805), .Y(\data_out<4> ) );
  BUFX2 U2455 ( .A(n4804), .Y(\data_out<5> ) );
  BUFX2 U2456 ( .A(n4803), .Y(\data_out<6> ) );
  BUFX2 U2457 ( .A(n4802), .Y(\data_out<7> ) );
  OR2X1 U2458 ( .A(N181), .B(n2678), .Y(n273) );
  INVX1 U2459 ( .A(n273), .Y(n274) );
  OR2X1 U2460 ( .A(N181), .B(N180), .Y(n275) );
  INVX1 U2461 ( .A(n275), .Y(n276) );
  INVX1 U2462 ( .A(n3739), .Y(n277) );
  INVX1 U2463 ( .A(n3740), .Y(n278) );
  INVX1 U2464 ( .A(n3741), .Y(n279) );
  INVX1 U2465 ( .A(n3742), .Y(n3200) );
  INVX1 U2466 ( .A(n3800), .Y(n280) );
  INVX1 U2467 ( .A(n3801), .Y(n281) );
  INVX1 U2468 ( .A(n3802), .Y(n282) );
  INVX1 U2469 ( .A(n3844), .Y(n283) );
  INVX1 U2470 ( .A(n3845), .Y(n284) );
  INVX1 U2471 ( .A(n3846), .Y(n285) );
  INVX1 U2472 ( .A(n3888), .Y(n286) );
  INVX1 U2473 ( .A(n3889), .Y(n287) );
  INVX1 U2474 ( .A(n3890), .Y(n288) );
  INVX1 U2475 ( .A(n3932), .Y(n289) );
  INVX1 U2476 ( .A(n3933), .Y(n290) );
  INVX1 U2477 ( .A(n3934), .Y(n291) );
  INVX1 U2478 ( .A(n3976), .Y(n292) );
  INVX1 U2479 ( .A(n3977), .Y(n293) );
  INVX1 U2480 ( .A(n3978), .Y(n294) );
  INVX1 U2481 ( .A(n4020), .Y(n295) );
  INVX1 U2482 ( .A(n4021), .Y(n296) );
  INVX1 U2483 ( .A(n4022), .Y(n297) );
  INVX1 U2484 ( .A(n4064), .Y(n298) );
  INVX1 U2485 ( .A(n4065), .Y(n299) );
  INVX1 U2486 ( .A(n4066), .Y(n300) );
  INVX1 U2487 ( .A(n3749), .Y(n301) );
  INVX1 U2488 ( .A(n3750), .Y(n302) );
  INVX1 U2489 ( .A(n3751), .Y(n303) );
  INVX1 U2490 ( .A(n3782), .Y(n304) );
  INVX1 U2491 ( .A(n3783), .Y(n305) );
  INVX1 U2492 ( .A(n3784), .Y(n306) );
  INVX1 U2493 ( .A(n3805), .Y(n307) );
  INVX1 U2494 ( .A(n3806), .Y(n308) );
  INVX1 U2495 ( .A(n3807), .Y(n309) );
  INVX1 U2496 ( .A(n3826), .Y(n310) );
  INVX1 U2497 ( .A(n3827), .Y(n311) );
  INVX1 U2498 ( .A(n3828), .Y(n312) );
  INVX1 U2499 ( .A(n3849), .Y(n313) );
  INVX1 U2500 ( .A(n3850), .Y(n314) );
  INVX1 U2501 ( .A(n3851), .Y(n315) );
  INVX1 U2502 ( .A(n3870), .Y(n316) );
  INVX1 U2503 ( .A(n3871), .Y(n317) );
  INVX1 U2504 ( .A(n3872), .Y(n318) );
  INVX1 U2505 ( .A(n3893), .Y(n319) );
  INVX1 U2506 ( .A(n3894), .Y(n320) );
  INVX1 U2507 ( .A(n3895), .Y(n321) );
  INVX1 U2508 ( .A(n3914), .Y(n322) );
  INVX1 U2509 ( .A(n3915), .Y(n323) );
  INVX1 U2510 ( .A(n3916), .Y(n324) );
  INVX1 U2511 ( .A(n3937), .Y(n325) );
  INVX1 U2512 ( .A(n3938), .Y(n326) );
  INVX1 U2513 ( .A(n3939), .Y(n327) );
  INVX1 U2514 ( .A(n3958), .Y(n328) );
  INVX1 U2515 ( .A(n3959), .Y(n329) );
  INVX1 U2516 ( .A(n3960), .Y(n330) );
  INVX1 U2517 ( .A(n3981), .Y(n331) );
  INVX1 U2518 ( .A(n3982), .Y(n332) );
  INVX1 U2519 ( .A(n3983), .Y(n333) );
  INVX1 U2520 ( .A(n4002), .Y(n334) );
  INVX1 U2521 ( .A(n4003), .Y(n335) );
  INVX1 U2522 ( .A(n4004), .Y(n336) );
  INVX1 U2523 ( .A(n4025), .Y(n337) );
  INVX1 U2524 ( .A(n4026), .Y(n338) );
  INVX1 U2525 ( .A(n4027), .Y(n339) );
  INVX1 U2526 ( .A(n4046), .Y(n340) );
  INVX1 U2527 ( .A(n4047), .Y(n341) );
  INVX1 U2528 ( .A(n4048), .Y(n342) );
  INVX1 U2529 ( .A(n4070), .Y(n343) );
  INVX1 U2530 ( .A(n4071), .Y(n344) );
  INVX1 U2531 ( .A(n4072), .Y(n345) );
  INVX1 U2532 ( .A(n4091), .Y(n346) );
  INVX1 U2533 ( .A(n4092), .Y(n347) );
  INVX1 U2534 ( .A(n4093), .Y(n348) );
  BUFX2 U2535 ( .A(n4127), .Y(n2611) );
  BUFX2 U2536 ( .A(n4138), .Y(n2612) );
  BUFX2 U2537 ( .A(n4149), .Y(n2613) );
  BUFX2 U2538 ( .A(n4160), .Y(n2614) );
  BUFX2 U2539 ( .A(n4171), .Y(n2615) );
  BUFX2 U2540 ( .A(n4182), .Y(n2616) );
  BUFX2 U2541 ( .A(n4193), .Y(n2617) );
  BUFX2 U2542 ( .A(n4204), .Y(n2618) );
  BUFX2 U2543 ( .A(n4215), .Y(n2619) );
  BUFX2 U2544 ( .A(n4226), .Y(n2620) );
  BUFX2 U2545 ( .A(n4237), .Y(n2621) );
  BUFX2 U2546 ( .A(n4248), .Y(n2622) );
  BUFX2 U2547 ( .A(n4259), .Y(n2623) );
  BUFX2 U2548 ( .A(n4270), .Y(n2624) );
  BUFX2 U2549 ( .A(n4281), .Y(n2625) );
  BUFX2 U2550 ( .A(n4292), .Y(n2626) );
  BUFX2 U2551 ( .A(n4303), .Y(n2627) );
  BUFX2 U2552 ( .A(n4314), .Y(n2628) );
  BUFX2 U2553 ( .A(n4325), .Y(n2629) );
  BUFX2 U2554 ( .A(n4336), .Y(n2630) );
  BUFX2 U2555 ( .A(n4347), .Y(n2631) );
  BUFX2 U2556 ( .A(n4358), .Y(n2632) );
  BUFX2 U2557 ( .A(n4369), .Y(n2633) );
  BUFX2 U2558 ( .A(n4380), .Y(n2634) );
  BUFX2 U2559 ( .A(n4391), .Y(n2635) );
  BUFX2 U2560 ( .A(n4402), .Y(n2636) );
  BUFX2 U2561 ( .A(n4413), .Y(n2637) );
  BUFX2 U2562 ( .A(n4424), .Y(n2638) );
  BUFX2 U2563 ( .A(n4435), .Y(n2639) );
  BUFX2 U2564 ( .A(n4446), .Y(n2640) );
  BUFX2 U2565 ( .A(n4457), .Y(n2641) );
  BUFX2 U2566 ( .A(n4468), .Y(n2642) );
  BUFX2 U2567 ( .A(n4479), .Y(n2643) );
  BUFX2 U2568 ( .A(n4490), .Y(n2644) );
  BUFX2 U2569 ( .A(n4501), .Y(n2645) );
  BUFX2 U2570 ( .A(n4512), .Y(n2646) );
  BUFX2 U2571 ( .A(n4523), .Y(n2647) );
  BUFX2 U2572 ( .A(n4534), .Y(n2648) );
  BUFX2 U2573 ( .A(n4545), .Y(n2649) );
  BUFX2 U2574 ( .A(n4556), .Y(n2650) );
  BUFX2 U2575 ( .A(n4567), .Y(n2651) );
  BUFX2 U2576 ( .A(n4578), .Y(n2652) );
  BUFX2 U2577 ( .A(n4589), .Y(n2653) );
  BUFX2 U2578 ( .A(n4600), .Y(n2654) );
  BUFX2 U2579 ( .A(n4611), .Y(n2655) );
  BUFX2 U2580 ( .A(n4622), .Y(n2656) );
  BUFX2 U2581 ( .A(n4633), .Y(n2657) );
  BUFX2 U2582 ( .A(n4644), .Y(n2658) );
  BUFX2 U2583 ( .A(n4655), .Y(n2659) );
  BUFX2 U2584 ( .A(n4666), .Y(n2660) );
  BUFX2 U2585 ( .A(n4677), .Y(n2661) );
  BUFX2 U2586 ( .A(n4688), .Y(n2662) );
  BUFX2 U2587 ( .A(n4699), .Y(n2663) );
  BUFX2 U2588 ( .A(n4710), .Y(n2664) );
  BUFX2 U2589 ( .A(n4721), .Y(n2665) );
  BUFX2 U2590 ( .A(n4732), .Y(n2666) );
  BUFX2 U2591 ( .A(n4743), .Y(n2667) );
  BUFX2 U2592 ( .A(n4754), .Y(n2668) );
  BUFX2 U2593 ( .A(n4765), .Y(n2669) );
  BUFX2 U2594 ( .A(n4776), .Y(n2670) );
  BUFX2 U2595 ( .A(n4788), .Y(n2671) );
  INVX1 U2596 ( .A(n4777), .Y(n2674) );
  INVX1 U2597 ( .A(rst), .Y(n2679) );
  AND2X1 U2598 ( .A(n3766), .B(n3200), .Y(n349) );
  INVX1 U2599 ( .A(n349), .Y(n350) );
  AND2X1 U2600 ( .A(n210), .B(n3773), .Y(n351) );
  INVX1 U2601 ( .A(n351), .Y(n352) );
  AND2X1 U2602 ( .A(n351), .B(n2674), .Y(n353) );
  INVX1 U2603 ( .A(n353), .Y(n354) );
  INVX1 U2604 ( .A(n356), .Y(n355) );
  AND2X1 U2605 ( .A(n3778), .B(n349), .Y(n356) );
  AND2X1 U2606 ( .A(n3196), .B(n3773), .Y(n357) );
  INVX1 U2607 ( .A(n357), .Y(n358) );
  AND2X1 U2608 ( .A(n3201), .B(n3195), .Y(n359) );
  INVX1 U2609 ( .A(n359), .Y(n360) );
  AND2X1 U2610 ( .A(n3196), .B(n3774), .Y(n361) );
  INVX1 U2611 ( .A(n361), .Y(n362) );
  AND2X1 U2612 ( .A(n3196), .B(n3775), .Y(n363) );
  INVX1 U2613 ( .A(n363), .Y(n364) );
  AND2X1 U2614 ( .A(n3196), .B(n3776), .Y(n365) );
  INVX1 U2615 ( .A(n365), .Y(n366) );
  AND2X1 U2616 ( .A(n3196), .B(n3777), .Y(n367) );
  INVX1 U2617 ( .A(n367), .Y(n368) );
  AND2X1 U2618 ( .A(n3196), .B(n3778), .Y(n369) );
  INVX1 U2619 ( .A(n369), .Y(n370) );
  AND2X1 U2620 ( .A(n3196), .B(n3779), .Y(n371) );
  INVX1 U2621 ( .A(n371), .Y(n372) );
  AND2X1 U2622 ( .A(n3201), .B(n3773), .Y(n373) );
  INVX1 U2623 ( .A(n373), .Y(n374) );
  INVX1 U2624 ( .A(n376), .Y(n375) );
  AND2X1 U2625 ( .A(n207), .B(n3195), .Y(n376) );
  AND2X1 U2626 ( .A(n3201), .B(n3774), .Y(n377) );
  INVX1 U2627 ( .A(n377), .Y(n378) );
  INVX1 U2628 ( .A(n380), .Y(n379) );
  AND2X1 U2629 ( .A(n3201), .B(n3775), .Y(n380) );
  AND2X1 U2630 ( .A(n3201), .B(n3776), .Y(n381) );
  INVX1 U2631 ( .A(n381), .Y(n382) );
  INVX1 U2632 ( .A(n384), .Y(n383) );
  AND2X1 U2633 ( .A(n3201), .B(n3777), .Y(n384) );
  AND2X1 U2634 ( .A(n3201), .B(n3778), .Y(n385) );
  INVX1 U2635 ( .A(n385), .Y(n386) );
  INVX1 U2636 ( .A(n388), .Y(n387) );
  AND2X1 U2637 ( .A(n3201), .B(n3779), .Y(n388) );
  AND2X1 U2638 ( .A(n207), .B(n3773), .Y(n389) );
  INVX1 U2639 ( .A(n389), .Y(n390) );
  AND2X1 U2640 ( .A(n210), .B(n3195), .Y(n391) );
  INVX1 U2641 ( .A(n391), .Y(n392) );
  AND2X1 U2642 ( .A(n207), .B(n3774), .Y(n393) );
  INVX1 U2643 ( .A(n393), .Y(n394) );
  INVX1 U2644 ( .A(n396), .Y(n395) );
  AND2X1 U2645 ( .A(n207), .B(n3775), .Y(n396) );
  AND2X1 U2646 ( .A(n207), .B(n3776), .Y(n397) );
  INVX1 U2647 ( .A(n397), .Y(n398) );
  INVX1 U2648 ( .A(n400), .Y(n399) );
  AND2X1 U2649 ( .A(n207), .B(n3777), .Y(n400) );
  AND2X1 U2650 ( .A(n207), .B(n3778), .Y(n401) );
  INVX1 U2651 ( .A(n401), .Y(n402) );
  INVX1 U2652 ( .A(n404), .Y(n403) );
  AND2X1 U2653 ( .A(n207), .B(n3779), .Y(n404) );
  AND2X1 U2654 ( .A(n210), .B(n3774), .Y(n405) );
  INVX1 U2655 ( .A(n405), .Y(n406) );
  AND2X1 U2656 ( .A(n210), .B(n3776), .Y(n407) );
  INVX1 U2657 ( .A(n407), .Y(n408) );
  AND2X1 U2658 ( .A(n210), .B(n3777), .Y(n409) );
  INVX1 U2659 ( .A(n409), .Y(n410) );
  AND2X1 U2660 ( .A(n210), .B(n3778), .Y(n411) );
  INVX1 U2661 ( .A(n411), .Y(n412) );
  AND2X1 U2662 ( .A(n210), .B(n3779), .Y(n413) );
  INVX1 U2663 ( .A(n413), .Y(n414) );
  AND2X1 U2664 ( .A(n3197), .B(n3773), .Y(n415) );
  INVX1 U2665 ( .A(n415), .Y(n416) );
  AND2X1 U2666 ( .A(n3199), .B(n3195), .Y(n417) );
  INVX1 U2667 ( .A(n417), .Y(n418) );
  AND2X1 U2668 ( .A(n3197), .B(n3774), .Y(n419) );
  INVX1 U2669 ( .A(n419), .Y(n420) );
  AND2X1 U2670 ( .A(n3197), .B(n3775), .Y(n421) );
  INVX1 U2671 ( .A(n421), .Y(n422) );
  AND2X1 U2672 ( .A(n3197), .B(n3776), .Y(n423) );
  INVX1 U2673 ( .A(n423), .Y(n424) );
  AND2X1 U2674 ( .A(n3197), .B(n3777), .Y(n425) );
  INVX1 U2675 ( .A(n425), .Y(n426) );
  AND2X1 U2676 ( .A(n3197), .B(n3778), .Y(n427) );
  INVX1 U2677 ( .A(n427), .Y(n428) );
  AND2X1 U2678 ( .A(n3197), .B(n3779), .Y(n429) );
  INVX1 U2679 ( .A(n429), .Y(n430) );
  AND2X1 U2680 ( .A(n3199), .B(n3773), .Y(n431) );
  INVX1 U2681 ( .A(n431), .Y(n432) );
  AND2X1 U2682 ( .A(n3196), .B(n3195), .Y(n433) );
  INVX1 U2683 ( .A(n433), .Y(n434) );
  AND2X1 U2684 ( .A(n3199), .B(n3774), .Y(n435) );
  INVX1 U2685 ( .A(n435), .Y(n436) );
  AND2X1 U2686 ( .A(n3199), .B(n3775), .Y(n437) );
  INVX1 U2687 ( .A(n437), .Y(n438) );
  AND2X1 U2688 ( .A(n3199), .B(n3776), .Y(n439) );
  INVX1 U2689 ( .A(n439), .Y(n440) );
  INVX1 U2690 ( .A(n442), .Y(n441) );
  AND2X1 U2691 ( .A(n3199), .B(n3777), .Y(n442) );
  AND2X1 U2692 ( .A(n3199), .B(n3778), .Y(n443) );
  INVX1 U2693 ( .A(n443), .Y(n444) );
  INVX1 U2694 ( .A(n446), .Y(n445) );
  AND2X1 U2695 ( .A(n3199), .B(n3779), .Y(n446) );
  INVX1 U2696 ( .A(n448), .Y(n447) );
  AND2X1 U2697 ( .A(n3773), .B(n349), .Y(n448) );
  AND2X1 U2698 ( .A(n3198), .B(n3195), .Y(n449) );
  INVX1 U2699 ( .A(n449), .Y(n450) );
  INVX1 U2700 ( .A(n452), .Y(n451) );
  AND2X1 U2701 ( .A(n3774), .B(n349), .Y(n452) );
  AND2X1 U2702 ( .A(n3775), .B(n349), .Y(n453) );
  INVX1 U2703 ( .A(n453), .Y(n454) );
  INVX1 U2704 ( .A(n456), .Y(n455) );
  AND2X1 U2705 ( .A(n3776), .B(n349), .Y(n456) );
  AND2X1 U2706 ( .A(n3777), .B(n349), .Y(n457) );
  INVX1 U2707 ( .A(n457), .Y(n458) );
  AND2X1 U2708 ( .A(n3779), .B(n349), .Y(n459) );
  INVX1 U2709 ( .A(n459), .Y(n460) );
  AND2X1 U2710 ( .A(n3198), .B(n3773), .Y(n461) );
  INVX1 U2711 ( .A(n461), .Y(n462) );
  AND2X1 U2712 ( .A(n3197), .B(n3195), .Y(n463) );
  INVX1 U2713 ( .A(n463), .Y(n464) );
  AND2X1 U2714 ( .A(n3198), .B(n3774), .Y(n465) );
  INVX1 U2715 ( .A(n465), .Y(n466) );
  AND2X1 U2716 ( .A(n3198), .B(n3775), .Y(n467) );
  INVX1 U2717 ( .A(n467), .Y(n468) );
  AND2X1 U2718 ( .A(n3198), .B(n3776), .Y(n469) );
  INVX1 U2719 ( .A(n469), .Y(n470) );
  AND2X1 U2720 ( .A(n3198), .B(n3777), .Y(n471) );
  INVX1 U2721 ( .A(n471), .Y(n472) );
  AND2X1 U2722 ( .A(n3198), .B(n3778), .Y(n473) );
  INVX1 U2723 ( .A(n473), .Y(n474) );
  AND2X1 U2724 ( .A(n3198), .B(n3779), .Y(n475) );
  INVX1 U2725 ( .A(n475), .Y(n476) );
  AND2X1 U2726 ( .A(n210), .B(n3775), .Y(n477) );
  INVX1 U2727 ( .A(n477), .Y(n478) );
  MUX2X1 U2728 ( .B(n480), .A(n481), .S(n2578), .Y(n479) );
  MUX2X1 U2729 ( .B(n483), .A(n484), .S(n2578), .Y(n482) );
  MUX2X1 U2730 ( .B(n486), .A(n487), .S(n2579), .Y(n485) );
  MUX2X1 U2731 ( .B(n489), .A(n490), .S(n2578), .Y(n488) );
  MUX2X1 U2732 ( .B(n492), .A(n493), .S(n2574), .Y(n491) );
  MUX2X1 U2733 ( .B(n495), .A(n496), .S(n2579), .Y(n494) );
  MUX2X1 U2734 ( .B(n498), .A(n499), .S(n2578), .Y(n497) );
  MUX2X1 U2735 ( .B(n501), .A(n502), .S(n2579), .Y(n500) );
  MUX2X1 U2736 ( .B(n504), .A(n505), .S(n2579), .Y(n503) );
  MUX2X1 U2737 ( .B(n507), .A(n508), .S(n2574), .Y(n506) );
  MUX2X1 U2738 ( .B(n510), .A(n511), .S(n2578), .Y(n509) );
  MUX2X1 U2739 ( .B(n513), .A(n514), .S(n2578), .Y(n512) );
  MUX2X1 U2740 ( .B(n516), .A(n517), .S(n2578), .Y(n515) );
  MUX2X1 U2741 ( .B(n519), .A(n520), .S(n2578), .Y(n518) );
  MUX2X1 U2742 ( .B(n522), .A(n523), .S(n2574), .Y(n521) );
  MUX2X1 U2743 ( .B(n525), .A(n526), .S(n2578), .Y(n524) );
  MUX2X1 U2744 ( .B(n528), .A(n529), .S(n2578), .Y(n527) );
  MUX2X1 U2745 ( .B(n531), .A(n532), .S(n2578), .Y(n530) );
  MUX2X1 U2746 ( .B(n534), .A(n535), .S(n2578), .Y(n533) );
  MUX2X1 U2747 ( .B(n537), .A(n538), .S(n2574), .Y(n536) );
  MUX2X1 U2748 ( .B(n539), .A(n540), .S(N182), .Y(N192) );
  MUX2X1 U2749 ( .B(n542), .A(n543), .S(n2578), .Y(n541) );
  MUX2X1 U2750 ( .B(n545), .A(n546), .S(n2578), .Y(n544) );
  MUX2X1 U2751 ( .B(n548), .A(n549), .S(n2578), .Y(n547) );
  MUX2X1 U2752 ( .B(n551), .A(n552), .S(n2578), .Y(n550) );
  MUX2X1 U2753 ( .B(n554), .A(n555), .S(n2574), .Y(n553) );
  MUX2X1 U2754 ( .B(n557), .A(n558), .S(n2579), .Y(n556) );
  MUX2X1 U2755 ( .B(n560), .A(n561), .S(n2579), .Y(n559) );
  MUX2X1 U2756 ( .B(n563), .A(n564), .S(n2579), .Y(n562) );
  MUX2X1 U2757 ( .B(n566), .A(n567), .S(n2579), .Y(n565) );
  MUX2X1 U2758 ( .B(n569), .A(n570), .S(n2574), .Y(n568) );
  MUX2X1 U2759 ( .B(n572), .A(n573), .S(n2579), .Y(n571) );
  MUX2X1 U2760 ( .B(n575), .A(n576), .S(n2579), .Y(n574) );
  MUX2X1 U2761 ( .B(n578), .A(n579), .S(n2579), .Y(n577) );
  MUX2X1 U2762 ( .B(n581), .A(n582), .S(n2579), .Y(n580) );
  MUX2X1 U2763 ( .B(n584), .A(n585), .S(n2574), .Y(n583) );
  MUX2X1 U2764 ( .B(n587), .A(n588), .S(n2579), .Y(n586) );
  MUX2X1 U2765 ( .B(n590), .A(n591), .S(n2579), .Y(n589) );
  MUX2X1 U2766 ( .B(n593), .A(n594), .S(n2579), .Y(n592) );
  MUX2X1 U2767 ( .B(n596), .A(n597), .S(n2579), .Y(n595) );
  MUX2X1 U2768 ( .B(n611), .A(n624), .S(n2574), .Y(n609) );
  MUX2X1 U2769 ( .B(n637), .A(n649), .S(N182), .Y(N191) );
  MUX2X1 U2770 ( .B(n673), .A(n685), .S(n2583), .Y(n661) );
  MUX2X1 U2771 ( .B(n709), .A(n721), .S(n2579), .Y(n697) );
  MUX2X1 U2772 ( .B(n745), .A(n757), .S(n2581), .Y(n733) );
  MUX2X1 U2773 ( .B(n781), .A(n793), .S(n2584), .Y(n769) );
  MUX2X1 U2774 ( .B(n817), .A(n829), .S(n2574), .Y(n805) );
  MUX2X1 U2775 ( .B(n853), .A(n865), .S(n2578), .Y(n841) );
  MUX2X1 U2776 ( .B(n889), .A(n901), .S(n2580), .Y(n877) );
  MUX2X1 U2777 ( .B(n925), .A(n937), .S(n2580), .Y(n913) );
  MUX2X1 U2778 ( .B(n961), .A(n973), .S(n2582), .Y(n949) );
  MUX2X1 U2779 ( .B(n997), .A(n1009), .S(n2574), .Y(n985) );
  MUX2X1 U2780 ( .B(n1033), .A(n1045), .S(n2580), .Y(n1021) );
  MUX2X1 U2781 ( .B(n1069), .A(n1081), .S(n2582), .Y(n1057) );
  MUX2X1 U2782 ( .B(n1105), .A(n1117), .S(n2582), .Y(n1093) );
  MUX2X1 U2783 ( .B(n1141), .A(n1153), .S(n2578), .Y(n1129) );
  MUX2X1 U2784 ( .B(n1177), .A(n1189), .S(n2574), .Y(n1165) );
  MUX2X1 U2785 ( .B(n1213), .A(n1225), .S(n2580), .Y(n1201) );
  MUX2X1 U2786 ( .B(n1249), .A(n1261), .S(n2580), .Y(n1237) );
  MUX2X1 U2787 ( .B(n1285), .A(n1297), .S(n2580), .Y(n1273) );
  MUX2X1 U2788 ( .B(n1321), .A(n1333), .S(n2580), .Y(n1309) );
  MUX2X1 U2789 ( .B(n1357), .A(n1358), .S(n2574), .Y(n1345) );
  MUX2X1 U2790 ( .B(n1371), .A(n1372), .S(N182), .Y(N190) );
  MUX2X1 U2791 ( .B(n1384), .A(n1396), .S(n2580), .Y(n1383) );
  MUX2X1 U2792 ( .B(n1409), .A(n1410), .S(n2580), .Y(n1397) );
  MUX2X1 U2793 ( .B(n1425), .A(n1436), .S(n2580), .Y(n1424) );
  MUX2X1 U2794 ( .B(n1449), .A(n1450), .S(n2580), .Y(n1437) );
  MUX2X1 U2795 ( .B(n1462), .A(n1476), .S(n2573), .Y(n1461) );
  MUX2X1 U2796 ( .B(n1488), .A(n1489), .S(n2580), .Y(n1477) );
  MUX2X1 U2797 ( .B(n1502), .A(n1513), .S(n2580), .Y(n1501) );
  MUX2X1 U2798 ( .B(n1528), .A(n1529), .S(n2580), .Y(n1514) );
  MUX2X1 U2799 ( .B(n1541), .A(n1553), .S(n2580), .Y(n1540) );
  MUX2X1 U2800 ( .B(n1565), .A(n1566), .S(n2573), .Y(n1554) );
  MUX2X1 U2801 ( .B(n1581), .A(n1592), .S(n2581), .Y(n1580) );
  MUX2X1 U2802 ( .B(n1605), .A(n1606), .S(n2581), .Y(n1593) );
  MUX2X1 U2803 ( .B(n1618), .A(n1632), .S(n2581), .Y(n1617) );
  MUX2X1 U2804 ( .B(n1644), .A(n1645), .S(n2581), .Y(n1633) );
  MUX2X1 U2805 ( .B(n1658), .A(n1669), .S(n2573), .Y(n1657) );
  MUX2X1 U2806 ( .B(n1684), .A(n1685), .S(n2581), .Y(n1670) );
  MUX2X1 U2807 ( .B(n1697), .A(n1709), .S(n2581), .Y(n1696) );
  MUX2X1 U2808 ( .B(n1721), .A(n1722), .S(n2581), .Y(n1710) );
  MUX2X1 U2809 ( .B(n1737), .A(n1758), .S(n2581), .Y(n1736) );
  MUX2X1 U2810 ( .B(n1771), .A(n1773), .S(n2573), .Y(n1759) );
  MUX2X1 U2811 ( .B(n1775), .A(n1776), .S(N182), .Y(N189) );
  MUX2X1 U2812 ( .B(n1793), .A(n1795), .S(n2581), .Y(n1783) );
  MUX2X1 U2813 ( .B(n1802), .A(n2328), .S(n2581), .Y(n1796) );
  MUX2X1 U2814 ( .B(n2330), .A(n2331), .S(n2581), .Y(n2329) );
  MUX2X1 U2815 ( .B(n2333), .A(n2334), .S(n2581), .Y(n2332) );
  MUX2X1 U2816 ( .B(n2336), .A(n2337), .S(n2573), .Y(n2335) );
  MUX2X1 U2817 ( .B(n2339), .A(n2340), .S(n2582), .Y(n2338) );
  MUX2X1 U2818 ( .B(n2342), .A(n2343), .S(n2582), .Y(n2341) );
  MUX2X1 U2819 ( .B(n2345), .A(n2346), .S(n2582), .Y(n2344) );
  MUX2X1 U2820 ( .B(n2348), .A(n2349), .S(n2582), .Y(n2347) );
  MUX2X1 U2821 ( .B(n2351), .A(n2352), .S(n2573), .Y(n2350) );
  MUX2X1 U2822 ( .B(n2354), .A(n2355), .S(n2582), .Y(n2353) );
  MUX2X1 U2823 ( .B(n2357), .A(n2358), .S(n2582), .Y(n2356) );
  MUX2X1 U2824 ( .B(n2360), .A(n2361), .S(n2582), .Y(n2359) );
  MUX2X1 U2825 ( .B(n2363), .A(n2364), .S(n2582), .Y(n2362) );
  MUX2X1 U2826 ( .B(n2366), .A(n2367), .S(n2573), .Y(n2365) );
  MUX2X1 U2827 ( .B(n2369), .A(n2370), .S(n2582), .Y(n2368) );
  MUX2X1 U2828 ( .B(n2372), .A(n2373), .S(n2582), .Y(n2371) );
  MUX2X1 U2829 ( .B(n2375), .A(n2376), .S(n2582), .Y(n2374) );
  MUX2X1 U2830 ( .B(n2378), .A(n2379), .S(n2582), .Y(n2377) );
  MUX2X1 U2831 ( .B(n2381), .A(n2382), .S(n2573), .Y(n2380) );
  MUX2X1 U2832 ( .B(n2383), .A(n2384), .S(N182), .Y(N188) );
  MUX2X1 U2833 ( .B(n2386), .A(n2387), .S(n2583), .Y(n2385) );
  MUX2X1 U2834 ( .B(n2389), .A(n2390), .S(n2583), .Y(n2388) );
  MUX2X1 U2835 ( .B(n2392), .A(n2393), .S(n2583), .Y(n2391) );
  MUX2X1 U2836 ( .B(n2395), .A(n2396), .S(n2583), .Y(n2394) );
  MUX2X1 U2837 ( .B(n2398), .A(n2399), .S(n2573), .Y(n2397) );
  MUX2X1 U2838 ( .B(n2401), .A(n2402), .S(n2583), .Y(n2400) );
  MUX2X1 U2839 ( .B(n2404), .A(n2405), .S(n2583), .Y(n2403) );
  MUX2X1 U2840 ( .B(n2407), .A(n2408), .S(n2583), .Y(n2406) );
  MUX2X1 U2841 ( .B(n2410), .A(n2411), .S(n2583), .Y(n2409) );
  MUX2X1 U2842 ( .B(n2413), .A(n2414), .S(n2573), .Y(n2412) );
  MUX2X1 U2843 ( .B(n2416), .A(n2417), .S(n2583), .Y(n2415) );
  MUX2X1 U2844 ( .B(n2419), .A(n2420), .S(n2583), .Y(n2418) );
  MUX2X1 U2845 ( .B(n2422), .A(n2423), .S(n2583), .Y(n2421) );
  MUX2X1 U2846 ( .B(n2425), .A(n2426), .S(n2583), .Y(n2424) );
  MUX2X1 U2847 ( .B(n2428), .A(n2429), .S(n2573), .Y(n2427) );
  MUX2X1 U2848 ( .B(n2431), .A(n2432), .S(n2584), .Y(n2430) );
  MUX2X1 U2849 ( .B(n2434), .A(n2435), .S(n2584), .Y(n2433) );
  MUX2X1 U2850 ( .B(n2437), .A(n2438), .S(n2584), .Y(n2436) );
  MUX2X1 U2851 ( .B(n2440), .A(n2441), .S(n2584), .Y(n2439) );
  MUX2X1 U2852 ( .B(n2443), .A(n2444), .S(n2573), .Y(n2442) );
  MUX2X1 U2853 ( .B(n2445), .A(n2446), .S(N182), .Y(N187) );
  MUX2X1 U2854 ( .B(n2448), .A(n2449), .S(n2584), .Y(n2447) );
  MUX2X1 U2855 ( .B(n2451), .A(n2452), .S(n2584), .Y(n2450) );
  MUX2X1 U2856 ( .B(n2454), .A(n2455), .S(n2584), .Y(n2453) );
  MUX2X1 U2857 ( .B(n2457), .A(n2458), .S(n2584), .Y(n2456) );
  MUX2X1 U2858 ( .B(n2460), .A(n2461), .S(n2573), .Y(n2459) );
  MUX2X1 U2859 ( .B(n2463), .A(n2464), .S(n2584), .Y(n2462) );
  MUX2X1 U2860 ( .B(n2466), .A(n2467), .S(n2584), .Y(n2465) );
  MUX2X1 U2861 ( .B(n2469), .A(n2470), .S(n2584), .Y(n2468) );
  MUX2X1 U2862 ( .B(n2472), .A(n2473), .S(n2584), .Y(n2471) );
  MUX2X1 U2863 ( .B(n2475), .A(n2476), .S(n2573), .Y(n2474) );
  MUX2X1 U2864 ( .B(n2478), .A(n2479), .S(n2584), .Y(n2477) );
  MUX2X1 U2865 ( .B(n2481), .A(n2482), .S(n2583), .Y(n2480) );
  MUX2X1 U2866 ( .B(n2484), .A(n2485), .S(n2580), .Y(n2483) );
  MUX2X1 U2867 ( .B(n2487), .A(n2488), .S(n2579), .Y(n2486) );
  MUX2X1 U2868 ( .B(n2490), .A(n2491), .S(n2573), .Y(n2489) );
  MUX2X1 U2869 ( .B(n2493), .A(n2494), .S(n2580), .Y(n2492) );
  MUX2X1 U2870 ( .B(n2496), .A(n2497), .S(n2581), .Y(n2495) );
  MUX2X1 U2871 ( .B(n2499), .A(n2500), .S(n2581), .Y(n2498) );
  MUX2X1 U2872 ( .B(n2502), .A(n2503), .S(n2581), .Y(n2501) );
  MUX2X1 U2873 ( .B(n2505), .A(n2506), .S(n2573), .Y(n2504) );
  MUX2X1 U2874 ( .B(n2507), .A(n2508), .S(N182), .Y(N186) );
  MUX2X1 U2875 ( .B(n2510), .A(n2511), .S(n2580), .Y(n2509) );
  MUX2X1 U2876 ( .B(n2513), .A(n2514), .S(n2580), .Y(n2512) );
  MUX2X1 U2877 ( .B(n2516), .A(n2517), .S(n2581), .Y(n2515) );
  MUX2X1 U2878 ( .B(n2519), .A(n2520), .S(n2581), .Y(n2518) );
  MUX2X1 U2879 ( .B(n2522), .A(n2523), .S(n2574), .Y(n2521) );
  MUX2X1 U2880 ( .B(n2525), .A(n2526), .S(n2583), .Y(n2524) );
  MUX2X1 U2881 ( .B(n2528), .A(n2529), .S(n2584), .Y(n2527) );
  MUX2X1 U2882 ( .B(n2531), .A(n2532), .S(n2584), .Y(n2530) );
  MUX2X1 U2883 ( .B(n2534), .A(n2535), .S(n2583), .Y(n2533) );
  MUX2X1 U2884 ( .B(n2537), .A(n2538), .S(n2574), .Y(n2536) );
  MUX2X1 U2885 ( .B(n2540), .A(n2541), .S(n2583), .Y(n2539) );
  MUX2X1 U2886 ( .B(n2543), .A(n2544), .S(n2582), .Y(n2542) );
  MUX2X1 U2887 ( .B(n2546), .A(n2547), .S(n2582), .Y(n2545) );
  MUX2X1 U2888 ( .B(n2549), .A(n2550), .S(n2582), .Y(n2548) );
  MUX2X1 U2889 ( .B(n2552), .A(n2553), .S(n2574), .Y(n2551) );
  MUX2X1 U2890 ( .B(n2555), .A(n2556), .S(n2583), .Y(n2554) );
  MUX2X1 U2891 ( .B(n2558), .A(n2559), .S(n2582), .Y(n2557) );
  MUX2X1 U2892 ( .B(n2561), .A(n2562), .S(n2584), .Y(n2560) );
  MUX2X1 U2893 ( .B(n2564), .A(n2565), .S(n2584), .Y(n2563) );
  MUX2X1 U2894 ( .B(n2567), .A(n2568), .S(n2574), .Y(n2566) );
  MUX2X1 U2895 ( .B(n2569), .A(n2570), .S(N182), .Y(N185) );
  MUX2X1 U2896 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n2591), .Y(n481) );
  MUX2X1 U2897 ( .B(\mem<60><0> ), .A(\mem<61><0> ), .S(n2593), .Y(n480) );
  MUX2X1 U2898 ( .B(\mem<58><0> ), .A(\mem<59><0> ), .S(n2593), .Y(n484) );
  MUX2X1 U2899 ( .B(\mem<56><0> ), .A(\mem<57><0> ), .S(n2593), .Y(n483) );
  MUX2X1 U2900 ( .B(n482), .A(n479), .S(n2577), .Y(n493) );
  MUX2X1 U2901 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n2590), .Y(n487) );
  MUX2X1 U2902 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n2590), .Y(n486) );
  MUX2X1 U2903 ( .B(\mem<50><0> ), .A(\mem<51><0> ), .S(n2590), .Y(n490) );
  MUX2X1 U2904 ( .B(\mem<48><0> ), .A(\mem<49><0> ), .S(n2590), .Y(n489) );
  MUX2X1 U2905 ( .B(n488), .A(n485), .S(n2577), .Y(n492) );
  MUX2X1 U2906 ( .B(\mem<46><0> ), .A(\mem<47><0> ), .S(n2590), .Y(n496) );
  MUX2X1 U2907 ( .B(\mem<44><0> ), .A(\mem<45><0> ), .S(n2590), .Y(n495) );
  MUX2X1 U2908 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n2590), .Y(n499) );
  MUX2X1 U2909 ( .B(\mem<40><0> ), .A(\mem<41><0> ), .S(n2590), .Y(n498) );
  MUX2X1 U2910 ( .B(n497), .A(n494), .S(n2577), .Y(n508) );
  MUX2X1 U2911 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n2590), .Y(n502) );
  MUX2X1 U2912 ( .B(\mem<36><0> ), .A(\mem<37><0> ), .S(n2590), .Y(n501) );
  MUX2X1 U2913 ( .B(\mem<34><0> ), .A(\mem<35><0> ), .S(n2590), .Y(n505) );
  MUX2X1 U2914 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n2590), .Y(n504) );
  MUX2X1 U2915 ( .B(n503), .A(n500), .S(n2577), .Y(n507) );
  MUX2X1 U2916 ( .B(n506), .A(n491), .S(n2572), .Y(n540) );
  MUX2X1 U2917 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n2590), .Y(n511) );
  MUX2X1 U2918 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n2590), .Y(n510) );
  MUX2X1 U2919 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n2590), .Y(n514) );
  MUX2X1 U2920 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n2590), .Y(n513) );
  MUX2X1 U2921 ( .B(n512), .A(n509), .S(n2577), .Y(n523) );
  MUX2X1 U2922 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n2590), .Y(n517) );
  MUX2X1 U2923 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n2590), .Y(n516) );
  MUX2X1 U2924 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n2590), .Y(n520) );
  MUX2X1 U2925 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n2590), .Y(n519) );
  MUX2X1 U2926 ( .B(n518), .A(n515), .S(n2577), .Y(n522) );
  MUX2X1 U2927 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n2590), .Y(n526) );
  MUX2X1 U2928 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n2590), .Y(n525) );
  MUX2X1 U2929 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n2590), .Y(n529) );
  MUX2X1 U2930 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n2590), .Y(n528) );
  MUX2X1 U2931 ( .B(n527), .A(n524), .S(n2577), .Y(n538) );
  MUX2X1 U2932 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n2591), .Y(n532) );
  MUX2X1 U2933 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n2591), .Y(n531) );
  MUX2X1 U2934 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n2591), .Y(n535) );
  MUX2X1 U2935 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n2591), .Y(n534) );
  MUX2X1 U2936 ( .B(n533), .A(n530), .S(n2577), .Y(n537) );
  MUX2X1 U2937 ( .B(n536), .A(n521), .S(n2572), .Y(n539) );
  MUX2X1 U2938 ( .B(\mem<62><1> ), .A(\mem<63><1> ), .S(n2591), .Y(n543) );
  MUX2X1 U2939 ( .B(\mem<60><1> ), .A(\mem<61><1> ), .S(n2591), .Y(n542) );
  MUX2X1 U2940 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n2591), .Y(n546) );
  MUX2X1 U2941 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n2591), .Y(n545) );
  MUX2X1 U2942 ( .B(n544), .A(n541), .S(n2577), .Y(n555) );
  MUX2X1 U2943 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n2591), .Y(n549) );
  MUX2X1 U2944 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n2591), .Y(n548) );
  MUX2X1 U2945 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n2591), .Y(n552) );
  MUX2X1 U2946 ( .B(\mem<48><1> ), .A(\mem<49><1> ), .S(n2591), .Y(n551) );
  MUX2X1 U2947 ( .B(n550), .A(n547), .S(n2577), .Y(n554) );
  MUX2X1 U2948 ( .B(\mem<46><1> ), .A(\mem<47><1> ), .S(n2592), .Y(n558) );
  MUX2X1 U2949 ( .B(\mem<44><1> ), .A(\mem<45><1> ), .S(n2592), .Y(n557) );
  MUX2X1 U2950 ( .B(\mem<42><1> ), .A(\mem<43><1> ), .S(n2592), .Y(n561) );
  MUX2X1 U2951 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n2592), .Y(n560) );
  MUX2X1 U2952 ( .B(n559), .A(n556), .S(n2577), .Y(n570) );
  MUX2X1 U2953 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n2592), .Y(n564) );
  MUX2X1 U2954 ( .B(\mem<36><1> ), .A(\mem<37><1> ), .S(n2592), .Y(n563) );
  MUX2X1 U2955 ( .B(\mem<34><1> ), .A(\mem<35><1> ), .S(n2592), .Y(n567) );
  MUX2X1 U2956 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n2592), .Y(n566) );
  MUX2X1 U2957 ( .B(n565), .A(n562), .S(n2577), .Y(n569) );
  MUX2X1 U2958 ( .B(n568), .A(n553), .S(n2572), .Y(n649) );
  MUX2X1 U2959 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n2592), .Y(n573) );
  MUX2X1 U2960 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n2592), .Y(n572) );
  MUX2X1 U2961 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n2592), .Y(n576) );
  MUX2X1 U2962 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n2592), .Y(n575) );
  MUX2X1 U2963 ( .B(n574), .A(n571), .S(n2576), .Y(n585) );
  MUX2X1 U2964 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n2593), .Y(n579) );
  MUX2X1 U2965 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2593), .Y(n578) );
  MUX2X1 U2966 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n2593), .Y(n582) );
  MUX2X1 U2967 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n2593), .Y(n581) );
  MUX2X1 U2968 ( .B(n580), .A(n577), .S(n2576), .Y(n584) );
  MUX2X1 U2969 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n2593), .Y(n588) );
  MUX2X1 U2970 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n2593), .Y(n587) );
  MUX2X1 U2971 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n2593), .Y(n591) );
  MUX2X1 U2972 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2593), .Y(n590) );
  MUX2X1 U2973 ( .B(n589), .A(n586), .S(n2576), .Y(n624) );
  MUX2X1 U2974 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n2593), .Y(n594) );
  MUX2X1 U2975 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n2593), .Y(n593) );
  MUX2X1 U2976 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n2593), .Y(n597) );
  MUX2X1 U2977 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n2593), .Y(n596) );
  MUX2X1 U2978 ( .B(n595), .A(n592), .S(n2576), .Y(n611) );
  MUX2X1 U2979 ( .B(n609), .A(n583), .S(n2572), .Y(n637) );
  MUX2X1 U2980 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n2594), .Y(n685) );
  MUX2X1 U2981 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n2594), .Y(n673) );
  MUX2X1 U2982 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n2594), .Y(n721) );
  MUX2X1 U2983 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n2594), .Y(n709) );
  MUX2X1 U2984 ( .B(n697), .A(n661), .S(n2576), .Y(n829) );
  MUX2X1 U2985 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n2594), .Y(n757) );
  MUX2X1 U2986 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n2594), .Y(n745) );
  MUX2X1 U2987 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n2594), .Y(n793) );
  MUX2X1 U2988 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n2594), .Y(n781) );
  MUX2X1 U2989 ( .B(n769), .A(n733), .S(n2576), .Y(n817) );
  MUX2X1 U2990 ( .B(\mem<46><2> ), .A(\mem<47><2> ), .S(n2594), .Y(n865) );
  MUX2X1 U2991 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n2594), .Y(n853) );
  MUX2X1 U2992 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n2594), .Y(n901) );
  MUX2X1 U2993 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n2594), .Y(n889) );
  MUX2X1 U2994 ( .B(n877), .A(n841), .S(n2576), .Y(n1009) );
  MUX2X1 U2995 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n2595), .Y(n937) );
  MUX2X1 U2996 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n2595), .Y(n925) );
  MUX2X1 U2997 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n2595), .Y(n973) );
  MUX2X1 U2998 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n2595), .Y(n961) );
  MUX2X1 U2999 ( .B(n949), .A(n913), .S(n2576), .Y(n997) );
  MUX2X1 U3000 ( .B(n985), .A(n805), .S(n2572), .Y(n1372) );
  MUX2X1 U3001 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2595), .Y(n1045) );
  MUX2X1 U3002 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n2595), .Y(n1033) );
  MUX2X1 U3003 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n2595), .Y(n1081) );
  MUX2X1 U3004 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n2595), .Y(n1069) );
  MUX2X1 U3005 ( .B(n1057), .A(n1021), .S(n2576), .Y(n1189) );
  MUX2X1 U3006 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2595), .Y(n1117) );
  MUX2X1 U3007 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n2595), .Y(n1105) );
  MUX2X1 U3008 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n2595), .Y(n1153) );
  MUX2X1 U3009 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n2595), .Y(n1141) );
  MUX2X1 U3010 ( .B(n1129), .A(n1093), .S(n2576), .Y(n1177) );
  MUX2X1 U3011 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2595), .Y(n1225) );
  MUX2X1 U3012 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n2595), .Y(n1213) );
  MUX2X1 U3013 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n2595), .Y(n1261) );
  MUX2X1 U3014 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n2595), .Y(n1249) );
  MUX2X1 U3015 ( .B(n1237), .A(n1201), .S(n2576), .Y(n1358) );
  MUX2X1 U3016 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n2594), .Y(n1297) );
  MUX2X1 U3017 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n2595), .Y(n1285) );
  MUX2X1 U3018 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n2595), .Y(n1333) );
  MUX2X1 U3019 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2594), .Y(n1321) );
  MUX2X1 U3020 ( .B(n1309), .A(n1273), .S(n2576), .Y(n1357) );
  MUX2X1 U3021 ( .B(n1345), .A(n1165), .S(n2572), .Y(n1371) );
  MUX2X1 U3022 ( .B(\mem<62><3> ), .A(\mem<63><3> ), .S(n2594), .Y(n1396) );
  MUX2X1 U3023 ( .B(\mem<60><3> ), .A(\mem<61><3> ), .S(n2594), .Y(n1384) );
  MUX2X1 U3024 ( .B(\mem<58><3> ), .A(\mem<59><3> ), .S(n2595), .Y(n1410) );
  MUX2X1 U3025 ( .B(\mem<56><3> ), .A(\mem<57><3> ), .S(n2594), .Y(n1409) );
  MUX2X1 U3026 ( .B(n1397), .A(n1383), .S(n2577), .Y(n1476) );
  MUX2X1 U3027 ( .B(\mem<54><3> ), .A(\mem<55><3> ), .S(n2596), .Y(n1436) );
  MUX2X1 U3028 ( .B(\mem<52><3> ), .A(\mem<53><3> ), .S(n2596), .Y(n1425) );
  MUX2X1 U3029 ( .B(\mem<50><3> ), .A(\mem<51><3> ), .S(n2596), .Y(n1450) );
  MUX2X1 U3030 ( .B(\mem<48><3> ), .A(\mem<49><3> ), .S(n2596), .Y(n1449) );
  MUX2X1 U3031 ( .B(n1437), .A(n1424), .S(n2577), .Y(n1462) );
  MUX2X1 U3032 ( .B(\mem<46><3> ), .A(\mem<47><3> ), .S(n2596), .Y(n1489) );
  MUX2X1 U3033 ( .B(\mem<44><3> ), .A(\mem<45><3> ), .S(n2596), .Y(n1488) );
  MUX2X1 U3034 ( .B(\mem<42><3> ), .A(\mem<43><3> ), .S(n2596), .Y(n1513) );
  MUX2X1 U3035 ( .B(\mem<40><3> ), .A(\mem<41><3> ), .S(n2596), .Y(n1502) );
  MUX2X1 U3036 ( .B(n1501), .A(n1477), .S(n2577), .Y(n1566) );
  MUX2X1 U3037 ( .B(\mem<38><3> ), .A(\mem<39><3> ), .S(n2596), .Y(n1529) );
  MUX2X1 U3038 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n2596), .Y(n1528) );
  MUX2X1 U3039 ( .B(\mem<34><3> ), .A(\mem<35><3> ), .S(n2596), .Y(n1553) );
  MUX2X1 U3040 ( .B(\mem<32><3> ), .A(\mem<33><3> ), .S(n2596), .Y(n1541) );
  MUX2X1 U3041 ( .B(n1540), .A(n1514), .S(n2577), .Y(n1565) );
  MUX2X1 U3042 ( .B(n1554), .A(n1461), .S(n2572), .Y(n1776) );
  MUX2X1 U3043 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n2597), .Y(n1592) );
  MUX2X1 U3044 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n2597), .Y(n1581) );
  MUX2X1 U3045 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2597), .Y(n1606) );
  MUX2X1 U3046 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n2597), .Y(n1605) );
  MUX2X1 U3047 ( .B(n1593), .A(n1580), .S(n2576), .Y(n1669) );
  MUX2X1 U3048 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n2597), .Y(n1632) );
  MUX2X1 U3049 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n2597), .Y(n1618) );
  MUX2X1 U3050 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n2597), .Y(n1645) );
  MUX2X1 U3051 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n2597), .Y(n1644) );
  MUX2X1 U3052 ( .B(n1633), .A(n1617), .S(n2577), .Y(n1658) );
  MUX2X1 U3053 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n2597), .Y(n1685) );
  MUX2X1 U3054 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n2597), .Y(n1684) );
  MUX2X1 U3055 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n2597), .Y(n1709) );
  MUX2X1 U3056 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n2597), .Y(n1697) );
  MUX2X1 U3057 ( .B(n1696), .A(n1670), .S(n2576), .Y(n1773) );
  MUX2X1 U3058 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n2598), .Y(n1722) );
  MUX2X1 U3059 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n2598), .Y(n1721) );
  MUX2X1 U3060 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n2598), .Y(n1758) );
  MUX2X1 U3061 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2598), .Y(n1737) );
  MUX2X1 U3062 ( .B(n1736), .A(n1710), .S(n2577), .Y(n1771) );
  MUX2X1 U3063 ( .B(n1759), .A(n1657), .S(n2572), .Y(n1775) );
  MUX2X1 U3064 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n2598), .Y(n1795) );
  MUX2X1 U3065 ( .B(\mem<60><4> ), .A(\mem<61><4> ), .S(n2598), .Y(n1793) );
  MUX2X1 U3066 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n2598), .Y(n2328) );
  MUX2X1 U3067 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n2598), .Y(n1802) );
  MUX2X1 U3068 ( .B(n1796), .A(n1783), .S(n2576), .Y(n2337) );
  MUX2X1 U3069 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n2598), .Y(n2331) );
  MUX2X1 U3070 ( .B(\mem<52><4> ), .A(\mem<53><4> ), .S(n2598), .Y(n2330) );
  MUX2X1 U3071 ( .B(\mem<50><4> ), .A(\mem<51><4> ), .S(n2598), .Y(n2334) );
  MUX2X1 U3072 ( .B(\mem<48><4> ), .A(\mem<49><4> ), .S(n2598), .Y(n2333) );
  MUX2X1 U3073 ( .B(n2332), .A(n2329), .S(n2576), .Y(n2336) );
  MUX2X1 U3074 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n2599), .Y(n2340) );
  MUX2X1 U3075 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n2599), .Y(n2339) );
  MUX2X1 U3076 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n2599), .Y(n2343) );
  MUX2X1 U3077 ( .B(\mem<40><4> ), .A(\mem<41><4> ), .S(n2599), .Y(n2342) );
  MUX2X1 U3078 ( .B(n2341), .A(n2338), .S(n2576), .Y(n2352) );
  MUX2X1 U3079 ( .B(\mem<38><4> ), .A(\mem<39><4> ), .S(n2599), .Y(n2346) );
  MUX2X1 U3080 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n2599), .Y(n2345) );
  MUX2X1 U3081 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n2599), .Y(n2349) );
  MUX2X1 U3082 ( .B(\mem<32><4> ), .A(\mem<33><4> ), .S(n2599), .Y(n2348) );
  MUX2X1 U3083 ( .B(n2347), .A(n2344), .S(n2576), .Y(n2351) );
  MUX2X1 U3084 ( .B(n2350), .A(n2335), .S(n2572), .Y(n2384) );
  MUX2X1 U3085 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n2599), .Y(n2355) );
  MUX2X1 U3086 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n2599), .Y(n2354) );
  MUX2X1 U3087 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n2599), .Y(n2358) );
  MUX2X1 U3088 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n2599), .Y(n2357) );
  MUX2X1 U3089 ( .B(n2356), .A(n2353), .S(n2575), .Y(n2367) );
  MUX2X1 U3090 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n2600), .Y(n2361) );
  MUX2X1 U3091 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2600), .Y(n2360) );
  MUX2X1 U3092 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n2600), .Y(n2364) );
  MUX2X1 U3093 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n2600), .Y(n2363) );
  MUX2X1 U3094 ( .B(n2362), .A(n2359), .S(n2575), .Y(n2366) );
  MUX2X1 U3095 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2600), .Y(n2370) );
  MUX2X1 U3096 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n2600), .Y(n2369) );
  MUX2X1 U3097 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n2600), .Y(n2373) );
  MUX2X1 U3098 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n2600), .Y(n2372) );
  MUX2X1 U3099 ( .B(n2371), .A(n2368), .S(n2575), .Y(n2382) );
  MUX2X1 U3100 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n2600), .Y(n2376) );
  MUX2X1 U3101 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2600), .Y(n2375) );
  MUX2X1 U3102 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n2600), .Y(n2379) );
  MUX2X1 U3103 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n2600), .Y(n2378) );
  MUX2X1 U3104 ( .B(n2377), .A(n2374), .S(n2575), .Y(n2381) );
  MUX2X1 U3105 ( .B(n2380), .A(n2365), .S(n2572), .Y(n2383) );
  MUX2X1 U3106 ( .B(\mem<62><5> ), .A(\mem<63><5> ), .S(n2601), .Y(n2387) );
  MUX2X1 U3107 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n2601), .Y(n2386) );
  MUX2X1 U3108 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n2601), .Y(n2390) );
  MUX2X1 U3109 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n2601), .Y(n2389) );
  MUX2X1 U3110 ( .B(n2388), .A(n2385), .S(n2575), .Y(n2399) );
  MUX2X1 U3111 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n2601), .Y(n2393) );
  MUX2X1 U3112 ( .B(\mem<52><5> ), .A(\mem<53><5> ), .S(n2601), .Y(n2392) );
  MUX2X1 U3113 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n2601), .Y(n2396) );
  MUX2X1 U3114 ( .B(\mem<48><5> ), .A(\mem<49><5> ), .S(n2601), .Y(n2395) );
  MUX2X1 U3115 ( .B(n2394), .A(n2391), .S(n2575), .Y(n2398) );
  MUX2X1 U3116 ( .B(\mem<46><5> ), .A(\mem<47><5> ), .S(n2601), .Y(n2402) );
  MUX2X1 U3117 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n2601), .Y(n2401) );
  MUX2X1 U3118 ( .B(\mem<42><5> ), .A(\mem<43><5> ), .S(n2601), .Y(n2405) );
  MUX2X1 U3119 ( .B(\mem<40><5> ), .A(\mem<41><5> ), .S(n2601), .Y(n2404) );
  MUX2X1 U3120 ( .B(n2403), .A(n2400), .S(n2575), .Y(n2414) );
  MUX2X1 U3121 ( .B(\mem<38><5> ), .A(\mem<39><5> ), .S(n2602), .Y(n2408) );
  MUX2X1 U3122 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n2602), .Y(n2407) );
  MUX2X1 U3123 ( .B(\mem<34><5> ), .A(\mem<35><5> ), .S(n2602), .Y(n2411) );
  MUX2X1 U3124 ( .B(\mem<32><5> ), .A(\mem<33><5> ), .S(n2602), .Y(n2410) );
  MUX2X1 U3125 ( .B(n2409), .A(n2406), .S(n2575), .Y(n2413) );
  MUX2X1 U3126 ( .B(n2412), .A(n2397), .S(n2572), .Y(n2446) );
  MUX2X1 U3127 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n2602), .Y(n2417) );
  MUX2X1 U3128 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n2602), .Y(n2416) );
  MUX2X1 U3129 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n2602), .Y(n2420) );
  MUX2X1 U3130 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n2602), .Y(n2419) );
  MUX2X1 U3131 ( .B(n2418), .A(n2415), .S(n2575), .Y(n2429) );
  MUX2X1 U3132 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n2602), .Y(n2423) );
  MUX2X1 U3133 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n2602), .Y(n2422) );
  MUX2X1 U3134 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n2602), .Y(n2426) );
  MUX2X1 U3135 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n2602), .Y(n2425) );
  MUX2X1 U3136 ( .B(n2424), .A(n2421), .S(n2575), .Y(n2428) );
  MUX2X1 U3137 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n2603), .Y(n2432) );
  MUX2X1 U3138 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n2603), .Y(n2431) );
  MUX2X1 U3139 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n2603), .Y(n2435) );
  MUX2X1 U3140 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n2603), .Y(n2434) );
  MUX2X1 U3141 ( .B(n2433), .A(n2430), .S(n2575), .Y(n2444) );
  MUX2X1 U3142 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n2603), .Y(n2438) );
  MUX2X1 U3143 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n2603), .Y(n2437) );
  MUX2X1 U3144 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n2603), .Y(n2441) );
  MUX2X1 U3145 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n2603), .Y(n2440) );
  MUX2X1 U3146 ( .B(n2439), .A(n2436), .S(n2575), .Y(n2443) );
  MUX2X1 U3147 ( .B(n2442), .A(n2427), .S(n2572), .Y(n2445) );
  MUX2X1 U3148 ( .B(\mem<62><6> ), .A(\mem<63><6> ), .S(n2603), .Y(n2449) );
  MUX2X1 U3149 ( .B(\mem<60><6> ), .A(\mem<61><6> ), .S(n2603), .Y(n2448) );
  MUX2X1 U3150 ( .B(\mem<58><6> ), .A(\mem<59><6> ), .S(n2603), .Y(n2452) );
  MUX2X1 U3151 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n2603), .Y(n2451) );
  MUX2X1 U3152 ( .B(n2450), .A(n2447), .S(n2577), .Y(n2461) );
  MUX2X1 U3153 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n2604), .Y(n2455) );
  MUX2X1 U3154 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n2604), .Y(n2454) );
  MUX2X1 U3155 ( .B(\mem<50><6> ), .A(\mem<51><6> ), .S(n2604), .Y(n2458) );
  MUX2X1 U3156 ( .B(\mem<48><6> ), .A(\mem<49><6> ), .S(n2604), .Y(n2457) );
  MUX2X1 U3157 ( .B(n2456), .A(n2453), .S(n2577), .Y(n2460) );
  MUX2X1 U3158 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n2604), .Y(n2464) );
  MUX2X1 U3159 ( .B(\mem<44><6> ), .A(\mem<45><6> ), .S(n2604), .Y(n2463) );
  MUX2X1 U3160 ( .B(\mem<42><6> ), .A(\mem<43><6> ), .S(n2604), .Y(n2467) );
  MUX2X1 U3161 ( .B(\mem<40><6> ), .A(\mem<41><6> ), .S(n2604), .Y(n2466) );
  MUX2X1 U3162 ( .B(n2465), .A(n2462), .S(n2575), .Y(n2476) );
  MUX2X1 U3163 ( .B(\mem<38><6> ), .A(\mem<39><6> ), .S(n2604), .Y(n2470) );
  MUX2X1 U3164 ( .B(\mem<36><6> ), .A(\mem<37><6> ), .S(n2604), .Y(n2469) );
  MUX2X1 U3165 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n2604), .Y(n2473) );
  MUX2X1 U3166 ( .B(\mem<32><6> ), .A(\mem<33><6> ), .S(n2604), .Y(n2472) );
  MUX2X1 U3167 ( .B(n2471), .A(n2468), .S(n2575), .Y(n2475) );
  MUX2X1 U3168 ( .B(n2474), .A(n2459), .S(n2572), .Y(n2508) );
  MUX2X1 U3169 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n2605), .Y(n2479) );
  MUX2X1 U3170 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n2605), .Y(n2478) );
  MUX2X1 U3171 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n2605), .Y(n2482) );
  MUX2X1 U3172 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n2605), .Y(n2481) );
  MUX2X1 U3173 ( .B(n2480), .A(n2477), .S(n2575), .Y(n2491) );
  MUX2X1 U3174 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n2605), .Y(n2485) );
  MUX2X1 U3175 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n2605), .Y(n2484) );
  MUX2X1 U3176 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n2605), .Y(n2488) );
  MUX2X1 U3177 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n2605), .Y(n2487) );
  MUX2X1 U3178 ( .B(n2486), .A(n2483), .S(n2576), .Y(n2490) );
  MUX2X1 U3179 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n2605), .Y(n2494) );
  MUX2X1 U3180 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n2605), .Y(n2493) );
  MUX2X1 U3181 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n2605), .Y(n2497) );
  MUX2X1 U3182 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n2605), .Y(n2496) );
  MUX2X1 U3183 ( .B(n2495), .A(n2492), .S(n2575), .Y(n2506) );
  MUX2X1 U3184 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n2606), .Y(n2500) );
  MUX2X1 U3185 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n2606), .Y(n2499) );
  MUX2X1 U3186 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n2606), .Y(n2503) );
  MUX2X1 U3187 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n2606), .Y(n2502) );
  MUX2X1 U3188 ( .B(n2501), .A(n2498), .S(n2577), .Y(n2505) );
  MUX2X1 U3189 ( .B(n2504), .A(n2489), .S(n2572), .Y(n2507) );
  MUX2X1 U3190 ( .B(\mem<62><7> ), .A(\mem<63><7> ), .S(n2606), .Y(n2511) );
  MUX2X1 U3191 ( .B(\mem<60><7> ), .A(\mem<61><7> ), .S(n2606), .Y(n2510) );
  MUX2X1 U3192 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n2606), .Y(n2514) );
  MUX2X1 U3193 ( .B(\mem<56><7> ), .A(\mem<57><7> ), .S(n2606), .Y(n2513) );
  MUX2X1 U3194 ( .B(n2512), .A(n2509), .S(n2575), .Y(n2523) );
  MUX2X1 U3195 ( .B(\mem<54><7> ), .A(\mem<55><7> ), .S(n2606), .Y(n2517) );
  MUX2X1 U3196 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n2606), .Y(n2516) );
  MUX2X1 U3197 ( .B(\mem<50><7> ), .A(\mem<51><7> ), .S(n2606), .Y(n2520) );
  MUX2X1 U3198 ( .B(\mem<48><7> ), .A(\mem<49><7> ), .S(n2606), .Y(n2519) );
  MUX2X1 U3199 ( .B(n2518), .A(n2515), .S(n2576), .Y(n2522) );
  MUX2X1 U3200 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n2607), .Y(n2526) );
  MUX2X1 U3201 ( .B(\mem<44><7> ), .A(\mem<45><7> ), .S(n2607), .Y(n2525) );
  MUX2X1 U3202 ( .B(\mem<42><7> ), .A(\mem<43><7> ), .S(n2607), .Y(n2529) );
  MUX2X1 U3203 ( .B(\mem<40><7> ), .A(\mem<41><7> ), .S(n2607), .Y(n2528) );
  MUX2X1 U3204 ( .B(n2527), .A(n2524), .S(n2575), .Y(n2538) );
  MUX2X1 U3205 ( .B(\mem<38><7> ), .A(\mem<39><7> ), .S(n2607), .Y(n2532) );
  MUX2X1 U3206 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n2607), .Y(n2531) );
  MUX2X1 U3207 ( .B(\mem<34><7> ), .A(\mem<35><7> ), .S(n2607), .Y(n2535) );
  MUX2X1 U3208 ( .B(\mem<32><7> ), .A(\mem<33><7> ), .S(n2607), .Y(n2534) );
  MUX2X1 U3209 ( .B(n2533), .A(n2530), .S(n2575), .Y(n2537) );
  MUX2X1 U3210 ( .B(n2536), .A(n2521), .S(n2572), .Y(n2570) );
  MUX2X1 U3211 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n2607), .Y(n2541) );
  MUX2X1 U3212 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n2607), .Y(n2540) );
  MUX2X1 U3213 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n2607), .Y(n2544) );
  MUX2X1 U3214 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n2607), .Y(n2543) );
  MUX2X1 U3215 ( .B(n2542), .A(n2539), .S(n2575), .Y(n2553) );
  MUX2X1 U3216 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n2592), .Y(n2547) );
  MUX2X1 U3217 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n2591), .Y(n2546) );
  MUX2X1 U3218 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n2591), .Y(n2550) );
  MUX2X1 U3219 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n2593), .Y(n2549) );
  MUX2X1 U3220 ( .B(n2548), .A(n2545), .S(n2575), .Y(n2552) );
  MUX2X1 U3221 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n2591), .Y(n2556) );
  MUX2X1 U3222 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n2593), .Y(n2555) );
  MUX2X1 U3223 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n2592), .Y(n2559) );
  MUX2X1 U3224 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n2593), .Y(n2558) );
  MUX2X1 U3225 ( .B(n2557), .A(n2554), .S(n2575), .Y(n2568) );
  MUX2X1 U3226 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n2591), .Y(n2562) );
  MUX2X1 U3227 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n2592), .Y(n2561) );
  MUX2X1 U3228 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n2591), .Y(n2565) );
  MUX2X1 U3229 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n2591), .Y(n2564) );
  MUX2X1 U3230 ( .B(n2563), .A(n2560), .S(n2576), .Y(n2567) );
  MUX2X1 U3231 ( .B(n2566), .A(n2551), .S(n2572), .Y(n2569) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module fetch ( .BranchPC({\BranchPC<15> , \BranchPC<14> , \BranchPC<13> , 
        \BranchPC<12> , \BranchPC<11> , \BranchPC<10> , \BranchPC<9> , 
        \BranchPC<8> , \BranchPC<7> , \BranchPC<6> , \BranchPC<5> , 
        \BranchPC<4> , \BranchPC<3> , \BranchPC<2> , \BranchPC<1> , 
        \BranchPC<0> }), BranchJumpTaken, clk, rst, Halt, Rti, Exception, 
        Stall, .Instr({\Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , 
        \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , 
        \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> , 
        \Instr<0> }), .IncPC({\IncPC<15> , \IncPC<14> , \IncPC<13> , 
        \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , 
        \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , 
        \IncPC<1> , \IncPC<0> }) );
  input \BranchPC<15> , \BranchPC<14> , \BranchPC<13> , \BranchPC<12> ,
         \BranchPC<11> , \BranchPC<10> , \BranchPC<9> , \BranchPC<8> ,
         \BranchPC<7> , \BranchPC<6> , \BranchPC<5> , \BranchPC<4> ,
         \BranchPC<3> , \BranchPC<2> , \BranchPC<1> , \BranchPC<0> ,
         BranchJumpTaken, clk, rst, Halt, Rti, Exception, Stall;
  output \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> , \Instr<11> ,
         \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> , \Instr<6> ,
         \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , \Instr<1> ,
         \Instr<0> , \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> ,
         \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> ,
         \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> ,
         \IncPC<1> , \IncPC<0> ;
  wire   \pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , \pc<10> , \pc<9> ,
         \pc<8> , \pc<7> , \pc<6> , \pc<5> , \pc<4> , \pc<3> , \pc<2> ,
         \pc<1> , \pc<0> , \nextEPC<15> , \nextEPC<14> , \nextEPC<13> ,
         \nextEPC<12> , \nextEPC<11> , \nextEPC<10> , \nextEPC<9> ,
         \nextEPC<8> , \nextEPC<7> , \nextEPC<6> , \nextEPC<5> , \nextEPC<4> ,
         \nextEPC<3> , \nextEPC<2> , \nextEPC<1> , \nextEPC<0> , \epc<15> ,
         \epc<14> , \epc<13> , \epc<12> , \epc<11> , \epc<10> , \epc<9> ,
         \epc<8> , \epc<7> , \epc<6> , \epc<5> , \epc<4> , \epc<3> , \epc<2> ,
         \epc<1> , \epc<0> , nextExcptState, curExcptState, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n58, n72, n78, n79, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73, n74,
         n75, n76, n77, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145;

  XOR2X1 U27 ( .A(curExcptState), .B(Exception), .Y(n24) );
  OAI21X1 U28 ( .A(n25), .B(n134), .C(n26), .Y(\nextEPC<9> ) );
  NAND2X1 U29 ( .A(\epc<9> ), .B(n25), .Y(n26) );
  OAI21X1 U30 ( .A(n25), .B(n133), .C(n27), .Y(\nextEPC<8> ) );
  NAND2X1 U31 ( .A(\epc<8> ), .B(n25), .Y(n27) );
  OAI21X1 U32 ( .A(n25), .B(n132), .C(n28), .Y(\nextEPC<7> ) );
  NAND2X1 U33 ( .A(\epc<7> ), .B(n25), .Y(n28) );
  OAI21X1 U34 ( .A(n25), .B(n131), .C(n29), .Y(\nextEPC<6> ) );
  NAND2X1 U35 ( .A(\epc<6> ), .B(n25), .Y(n29) );
  OAI21X1 U36 ( .A(n25), .B(n130), .C(n30), .Y(\nextEPC<5> ) );
  NAND2X1 U37 ( .A(\epc<5> ), .B(n25), .Y(n30) );
  OAI21X1 U38 ( .A(n25), .B(n129), .C(n31), .Y(\nextEPC<4> ) );
  NAND2X1 U39 ( .A(\epc<4> ), .B(n25), .Y(n31) );
  OAI21X1 U40 ( .A(n25), .B(n142), .C(n32), .Y(\nextEPC<3> ) );
  NAND2X1 U41 ( .A(\epc<3> ), .B(n25), .Y(n32) );
  OAI21X1 U42 ( .A(n25), .B(n141), .C(n33), .Y(\nextEPC<2> ) );
  NAND2X1 U43 ( .A(\epc<2> ), .B(n25), .Y(n33) );
  OAI21X1 U44 ( .A(n25), .B(n143), .C(n34), .Y(\nextEPC<1> ) );
  NAND2X1 U45 ( .A(\epc<1> ), .B(n25), .Y(n34) );
  OAI21X1 U46 ( .A(n25), .B(n140), .C(n35), .Y(\nextEPC<15> ) );
  NAND2X1 U47 ( .A(\epc<15> ), .B(n25), .Y(n35) );
  OAI21X1 U48 ( .A(n25), .B(n139), .C(n36), .Y(\nextEPC<14> ) );
  NAND2X1 U49 ( .A(\epc<14> ), .B(n25), .Y(n36) );
  OAI21X1 U50 ( .A(n25), .B(n138), .C(n37), .Y(\nextEPC<13> ) );
  NAND2X1 U51 ( .A(\epc<13> ), .B(n25), .Y(n37) );
  OAI21X1 U52 ( .A(n25), .B(n137), .C(n38), .Y(\nextEPC<12> ) );
  NAND2X1 U53 ( .A(\epc<12> ), .B(n25), .Y(n38) );
  OAI21X1 U54 ( .A(n25), .B(n136), .C(n39), .Y(\nextEPC<11> ) );
  NAND2X1 U55 ( .A(\epc<11> ), .B(n25), .Y(n39) );
  OAI21X1 U56 ( .A(n25), .B(n135), .C(n40), .Y(\nextEPC<10> ) );
  NAND2X1 U57 ( .A(\epc<10> ), .B(n25), .Y(n40) );
  OAI21X1 U58 ( .A(n25), .B(n145), .C(n41), .Y(\nextEPC<0> ) );
  NAND2X1 U59 ( .A(\epc<0> ), .B(n25), .Y(n41) );
  AOI22X1 U86 ( .A(\IncPC<1> ), .B(n97), .C(\BranchPC<1> ), .D(n95), .Y(n58)
         );
  AOI22X1 U107 ( .A(\IncPC<0> ), .B(n97), .C(\BranchPC<0> ), .D(n95), .Y(n72)
         );
  NOR2X1 U110 ( .A(Stall), .B(Halt), .Y(n78) );
  NOR2X1 U112 ( .A(n105), .B(Halt), .Y(n79) );
  dff_388 \pc_reg[0]  ( .q(\pc<0> ), .d(n89), .clk(clk), .rst(n105) );
  dff_389 \pc_reg[1]  ( .q(\pc<1> ), .d(n91), .clk(clk), .rst(n105) );
  dff_390 \pc_reg[2]  ( .q(\pc<2> ), .d(n44), .clk(clk), .rst(n104) );
  dff_391 \pc_reg[3]  ( .q(\pc<3> ), .d(n42), .clk(clk), .rst(n104) );
  dff_392 \pc_reg[4]  ( .q(\pc<4> ), .d(n22), .clk(clk), .rst(n104) );
  dff_393 \pc_reg[5]  ( .q(\pc<5> ), .d(n20), .clk(clk), .rst(n104) );
  dff_394 \pc_reg[6]  ( .q(\pc<6> ), .d(n18), .clk(clk), .rst(n104) );
  dff_395 \pc_reg[7]  ( .q(\pc<7> ), .d(n16), .clk(clk), .rst(n104) );
  dff_396 \pc_reg[8]  ( .q(\pc<8> ), .d(n14), .clk(clk), .rst(n104) );
  dff_397 \pc_reg[9]  ( .q(\pc<9> ), .d(n46), .clk(clk), .rst(n104) );
  dff_398 \pc_reg[10]  ( .q(\pc<10> ), .d(n12), .clk(clk), .rst(n104) );
  dff_399 \pc_reg[11]  ( .q(\pc<11> ), .d(n10), .clk(clk), .rst(n104) );
  dff_400 \pc_reg[12]  ( .q(\pc<12> ), .d(n8), .clk(clk), .rst(n105) );
  dff_401 \pc_reg[13]  ( .q(\pc<13> ), .d(n6), .clk(clk), .rst(n105) );
  dff_402 \pc_reg[14]  ( .q(\pc<14> ), .d(n4), .clk(clk), .rst(n104) );
  dff_403 \pc_reg[15]  ( .q(\pc<15> ), .d(n2), .clk(clk), .rst(n105) );
  dff_372 \epc_reg[0]  ( .q(\epc<0> ), .d(\nextEPC<0> ), .clk(clk), .rst(n105)
         );
  dff_373 \epc_reg[1]  ( .q(\epc<1> ), .d(\nextEPC<1> ), .clk(clk), .rst(n105)
         );
  dff_374 \epc_reg[2]  ( .q(\epc<2> ), .d(\nextEPC<2> ), .clk(clk), .rst(n105)
         );
  dff_375 \epc_reg[3]  ( .q(\epc<3> ), .d(\nextEPC<3> ), .clk(clk), .rst(n105)
         );
  dff_376 \epc_reg[4]  ( .q(\epc<4> ), .d(\nextEPC<4> ), .clk(clk), .rst(n105)
         );
  dff_377 \epc_reg[5]  ( .q(\epc<5> ), .d(\nextEPC<5> ), .clk(clk), .rst(n105)
         );
  dff_378 \epc_reg[6]  ( .q(\epc<6> ), .d(\nextEPC<6> ), .clk(clk), .rst(n105)
         );
  dff_379 \epc_reg[7]  ( .q(\epc<7> ), .d(\nextEPC<7> ), .clk(clk), .rst(n105)
         );
  dff_380 \epc_reg[8]  ( .q(\epc<8> ), .d(\nextEPC<8> ), .clk(clk), .rst(n105)
         );
  dff_381 \epc_reg[9]  ( .q(\epc<9> ), .d(\nextEPC<9> ), .clk(clk), .rst(n105)
         );
  dff_382 \epc_reg[10]  ( .q(\epc<10> ), .d(\nextEPC<10> ), .clk(clk), .rst(
        n105) );
  dff_383 \epc_reg[11]  ( .q(\epc<11> ), .d(\nextEPC<11> ), .clk(clk), .rst(
        n105) );
  dff_384 \epc_reg[12]  ( .q(\epc<12> ), .d(\nextEPC<12> ), .clk(clk), .rst(
        n105) );
  dff_385 \epc_reg[13]  ( .q(\epc<13> ), .d(\nextEPC<13> ), .clk(clk), .rst(
        n105) );
  dff_386 \epc_reg[14]  ( .q(\epc<14> ), .d(\nextEPC<14> ), .clk(clk), .rst(
        n105) );
  dff_387 \epc_reg[15]  ( .q(\epc<15> ), .d(\nextEPC<15> ), .clk(clk), .rst(
        n105) );
  dff_404 excpt_reg ( .q(curExcptState), .d(nextExcptState), .clk(clk), .rst(
        n105) );
  memory2c_1 instr_mem ( .data_out({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , 
        \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , 
        \Instr<1> , \Instr<0> }), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .addr({
        \pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , \pc<10> , \pc<9> , 
        \pc<8> , \pc<7> , \pc<6> , \pc<5> , n102, n100, n98, \pc<1> , \pc<0> }), .enable(1'b1), .wr(1'b0), .createdump(1'b0), .clk(clk), .rst(n104) );
  cla16_2 pc_inc ( .A({\pc<15> , \pc<14> , \pc<13> , \pc<12> , \pc<11> , 
        \pc<10> , \pc<9> , \pc<8> , \pc<7> , \pc<6> , \pc<5> , n102, n100, n98, 
        \pc<1> , \pc<0> }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .Cin(1'b0), .S({
        \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> , 
        \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> , 
        \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> }), .Cout() );
  INVX1 U3 ( .A(\pc<2> ), .Y(n99) );
  INVX1 U4 ( .A(\pc<4> ), .Y(n103) );
  INVX1 U5 ( .A(rst), .Y(n106) );
  INVX1 U6 ( .A(n106), .Y(n104) );
  INVX1 U7 ( .A(\IncPC<3> ), .Y(n142) );
  INVX1 U8 ( .A(\IncPC<5> ), .Y(n130) );
  INVX1 U9 ( .A(\IncPC<6> ), .Y(n131) );
  INVX1 U10 ( .A(\IncPC<7> ), .Y(n132) );
  INVX1 U11 ( .A(\IncPC<8> ), .Y(n133) );
  INVX1 U12 ( .A(\IncPC<9> ), .Y(n134) );
  INVX1 U13 ( .A(\IncPC<10> ), .Y(n135) );
  INVX1 U14 ( .A(\IncPC<12> ), .Y(n137) );
  INVX1 U15 ( .A(\IncPC<13> ), .Y(n138) );
  INVX1 U16 ( .A(\IncPC<14> ), .Y(n139) );
  INVX1 U17 ( .A(Rti), .Y(n144) );
  BUFX2 U18 ( .A(n128), .Y(n95) );
  INVX1 U19 ( .A(\pc<3> ), .Y(n101) );
  INVX1 U20 ( .A(\IncPC<11> ), .Y(n136) );
  INVX1 U21 ( .A(\IncPC<15> ), .Y(n140) );
  INVX1 U22 ( .A(\IncPC<0> ), .Y(n145) );
  INVX1 U23 ( .A(\IncPC<1> ), .Y(n143) );
  INVX1 U24 ( .A(\IncPC<2> ), .Y(n141) );
  INVX1 U25 ( .A(\IncPC<4> ), .Y(n129) );
  AND2X1 U26 ( .A(n24), .B(n144), .Y(nextExcptState) );
  INVX2 U60 ( .A(n99), .Y(n98) );
  AND2X1 U61 ( .A(curExcptState), .B(n144), .Y(n25) );
  BUFX2 U62 ( .A(n126), .Y(n96) );
  AND2X2 U63 ( .A(n111), .B(n60), .Y(n1) );
  INVX1 U64 ( .A(n1), .Y(n2) );
  AND2X2 U65 ( .A(n112), .B(n62), .Y(n3) );
  INVX1 U66 ( .A(n3), .Y(n4) );
  AND2X2 U67 ( .A(n113), .B(n114), .Y(n5) );
  INVX1 U68 ( .A(n5), .Y(n6) );
  AND2X2 U69 ( .A(n115), .B(n64), .Y(n7) );
  INVX1 U70 ( .A(n7), .Y(n8) );
  AND2X2 U71 ( .A(n116), .B(n66), .Y(n9) );
  INVX1 U72 ( .A(n9), .Y(n10) );
  AND2X2 U73 ( .A(n117), .B(n68), .Y(n11) );
  INVX1 U74 ( .A(n11), .Y(n12) );
  AND2X2 U75 ( .A(n119), .B(n73), .Y(n13) );
  INVX1 U76 ( .A(n13), .Y(n14) );
  AND2X2 U77 ( .A(n120), .B(n75), .Y(n15) );
  INVX1 U78 ( .A(n15), .Y(n16) );
  AND2X2 U79 ( .A(n121), .B(n77), .Y(n17) );
  INVX1 U80 ( .A(n17), .Y(n18) );
  AND2X2 U81 ( .A(n122), .B(n81), .Y(n19) );
  INVX1 U82 ( .A(n19), .Y(n20) );
  AND2X2 U83 ( .A(n123), .B(n83), .Y(n21) );
  INVX1 U84 ( .A(n21), .Y(n22) );
  AND2X2 U85 ( .A(n124), .B(n85), .Y(n23) );
  INVX1 U87 ( .A(n23), .Y(n42) );
  AND2X2 U88 ( .A(n125), .B(n87), .Y(n43) );
  INVX1 U89 ( .A(n43), .Y(n44) );
  AND2X2 U90 ( .A(n118), .B(n70), .Y(n45) );
  INVX1 U91 ( .A(n45), .Y(n46) );
  OR2X2 U92 ( .A(n93), .B(n128), .Y(n47) );
  INVX1 U93 ( .A(n47), .Y(n48) );
  AND2X2 U94 ( .A(\pc<0> ), .B(n93), .Y(n49) );
  INVX1 U95 ( .A(n49), .Y(n50) );
  AND2X2 U96 ( .A(\pc<1> ), .B(n93), .Y(n51) );
  INVX1 U97 ( .A(n51), .Y(n52) );
  BUFX2 U98 ( .A(n72), .Y(n53) );
  BUFX2 U99 ( .A(n58), .Y(n54) );
  INVX1 U100 ( .A(n106), .Y(n105) );
  OR2X1 U101 ( .A(Stall), .B(n109), .Y(n55) );
  INVX1 U102 ( .A(n55), .Y(n56) );
  BUFX2 U103 ( .A(n110), .Y(n57) );
  AND2X2 U104 ( .A(\BranchPC<15> ), .B(n95), .Y(n59) );
  INVX1 U105 ( .A(n59), .Y(n60) );
  AND2X2 U106 ( .A(\BranchPC<14> ), .B(n95), .Y(n61) );
  INVX1 U108 ( .A(n61), .Y(n62) );
  AND2X2 U109 ( .A(\BranchPC<12> ), .B(n95), .Y(n63) );
  INVX1 U111 ( .A(n63), .Y(n64) );
  AND2X2 U113 ( .A(\BranchPC<11> ), .B(n95), .Y(n65) );
  INVX1 U114 ( .A(n65), .Y(n66) );
  AND2X2 U115 ( .A(\BranchPC<10> ), .B(n95), .Y(n67) );
  INVX1 U116 ( .A(n67), .Y(n68) );
  AND2X2 U117 ( .A(\BranchPC<9> ), .B(n95), .Y(n69) );
  INVX1 U118 ( .A(n69), .Y(n70) );
  AND2X2 U119 ( .A(\BranchPC<8> ), .B(n95), .Y(n71) );
  INVX1 U120 ( .A(n71), .Y(n73) );
  AND2X2 U121 ( .A(\BranchPC<7> ), .B(n95), .Y(n74) );
  INVX1 U122 ( .A(n74), .Y(n75) );
  AND2X2 U123 ( .A(\BranchPC<6> ), .B(n95), .Y(n76) );
  INVX1 U124 ( .A(n76), .Y(n77) );
  AND2X2 U125 ( .A(\BranchPC<5> ), .B(n95), .Y(n80) );
  INVX1 U126 ( .A(n80), .Y(n81) );
  AND2X2 U127 ( .A(\BranchPC<4> ), .B(n95), .Y(n82) );
  INVX1 U128 ( .A(n82), .Y(n83) );
  AND2X2 U129 ( .A(\BranchPC<3> ), .B(n95), .Y(n84) );
  INVX1 U130 ( .A(n84), .Y(n85) );
  AND2X2 U131 ( .A(\BranchPC<2> ), .B(n95), .Y(n86) );
  INVX1 U132 ( .A(n86), .Y(n87) );
  AND2X2 U133 ( .A(n50), .B(n53), .Y(n88) );
  INVX1 U134 ( .A(n88), .Y(n89) );
  AND2X2 U135 ( .A(n52), .B(n54), .Y(n90) );
  INVX1 U136 ( .A(n90), .Y(n91) );
  INVX2 U137 ( .A(n127), .Y(n92) );
  INVX8 U138 ( .A(n92), .Y(n93) );
  INVX1 U139 ( .A(n108), .Y(n127) );
  INVX1 U140 ( .A(BranchJumpTaken), .Y(n109) );
  AND2X2 U141 ( .A(\BranchPC<13> ), .B(n128), .Y(n94) );
  INVX1 U142 ( .A(n94), .Y(n114) );
  BUFX4 U143 ( .A(n126), .Y(n97) );
  INVX8 U144 ( .A(n101), .Y(n100) );
  INVX8 U145 ( .A(n103), .Y(n102) );
  NOR2X1 U146 ( .A(Halt), .B(n105), .Y(n107) );
  AND2X2 U147 ( .A(n107), .B(n56), .Y(n128) );
  NAND3X1 U148 ( .A(n79), .B(Stall), .C(n109), .Y(n108) );
  NAND3X1 U149 ( .A(n105), .B(n78), .C(n109), .Y(n110) );
  AND2X2 U150 ( .A(n48), .B(n57), .Y(n126) );
  AOI22X1 U151 ( .A(\pc<15> ), .B(n93), .C(\IncPC<15> ), .D(n96), .Y(n111) );
  AOI22X1 U152 ( .A(\pc<14> ), .B(n93), .C(\IncPC<14> ), .D(n96), .Y(n112) );
  AOI22X1 U153 ( .A(\pc<13> ), .B(n93), .C(\IncPC<13> ), .D(n96), .Y(n113) );
  AOI22X1 U154 ( .A(\pc<12> ), .B(n93), .C(\IncPC<12> ), .D(n96), .Y(n115) );
  AOI22X1 U155 ( .A(\pc<11> ), .B(n93), .C(\IncPC<11> ), .D(n96), .Y(n116) );
  AOI22X1 U156 ( .A(\pc<10> ), .B(n93), .C(\IncPC<10> ), .D(n96), .Y(n117) );
  AOI22X1 U157 ( .A(\pc<9> ), .B(n93), .C(\IncPC<9> ), .D(n96), .Y(n118) );
  AOI22X1 U158 ( .A(\pc<8> ), .B(n93), .C(\IncPC<8> ), .D(n96), .Y(n119) );
  AOI22X1 U159 ( .A(\pc<7> ), .B(n93), .C(\IncPC<7> ), .D(n97), .Y(n120) );
  AOI22X1 U160 ( .A(\pc<6> ), .B(n93), .C(\IncPC<6> ), .D(n97), .Y(n121) );
  AOI22X1 U161 ( .A(\pc<5> ), .B(n93), .C(\IncPC<5> ), .D(n97), .Y(n122) );
  AOI22X1 U162 ( .A(n102), .B(n93), .C(\IncPC<4> ), .D(n97), .Y(n123) );
  AOI22X1 U163 ( .A(n100), .B(n93), .C(\IncPC<3> ), .D(n97), .Y(n124) );
  AOI22X1 U164 ( .A(n98), .B(n93), .C(\IncPC<2> ), .D(n97), .Y(n125) );
endmodule


module pipe_fd ( Stall, Flush, rst, clk, .Instr({\Instr<15> , \Instr<14> , 
        \Instr<13> , \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , 
        \Instr<8> , \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , 
        \Instr<2> , \Instr<1> , \Instr<0> }), .IncPC({\IncPC<15> , \IncPC<14> , 
        \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , 
        \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , 
        \IncPC<2> , \IncPC<1> , \IncPC<0> }), .Instr_Out({\Instr_Out<15> , 
        \Instr_Out<14> , \Instr_Out<13> , \Instr_Out<12> , \Instr_Out<11> , 
        \Instr_Out<10> , \Instr_Out<9> , \Instr_Out<8> , \Instr_Out<7> , 
        \Instr_Out<6> , \Instr_Out<5> , \Instr_Out<4> , \Instr_Out<3> , 
        \Instr_Out<2> , \Instr_Out<1> , \Instr_Out<0> }), .IncPC_Out({
        \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> , \IncPC_Out<12> , 
        \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> , \IncPC_Out<8> , 
        \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> , \IncPC_Out<4> , 
        \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> , \IncPC_Out<0> }), 
        CPUActive );
  input Stall, Flush, rst, clk, \Instr<15> , \Instr<14> , \Instr<13> ,
         \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> ,
         \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> ,
         \Instr<2> , \Instr<1> , \Instr<0> , \IncPC<15> , \IncPC<14> ,
         \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> ,
         \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> ,
         \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> ;
  output \Instr_Out<15> , \Instr_Out<14> , \Instr_Out<13> , \Instr_Out<12> ,
         \Instr_Out<11> , \Instr_Out<10> , \Instr_Out<9> , \Instr_Out<8> ,
         \Instr_Out<7> , \Instr_Out<6> , \Instr_Out<5> , \Instr_Out<4> ,
         \Instr_Out<3> , \Instr_Out<2> , \Instr_Out<1> , \Instr_Out<0> ,
         \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> , \IncPC_Out<12> ,
         \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> , \IncPC_Out<8> ,
         \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> , \IncPC_Out<4> ,
         \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> , \IncPC_Out<0> ,
         CPUActive;
  wire   \Instr_Muxed<11> , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n70, n71, n72, n73, n74, n75;

  AOI22X1 U37 ( .A(\Instr_Out<9> ), .B(n4), .C(\Instr<9> ), .D(n5), .Y(n36) );
  AOI22X1 U38 ( .A(\Instr_Out<8> ), .B(n4), .C(\Instr<8> ), .D(n5), .Y(n39) );
  AOI22X1 U39 ( .A(\Instr_Out<7> ), .B(n4), .C(\Instr<7> ), .D(n5), .Y(n40) );
  AOI22X1 U40 ( .A(\Instr_Out<6> ), .B(n4), .C(\Instr<6> ), .D(n5), .Y(n41) );
  AOI22X1 U41 ( .A(\Instr_Out<5> ), .B(n4), .C(\Instr<5> ), .D(n5), .Y(n42) );
  AOI22X1 U42 ( .A(\Instr_Out<4> ), .B(n4), .C(\Instr<4> ), .D(n5), .Y(n43) );
  AOI22X1 U43 ( .A(\Instr_Out<3> ), .B(n4), .C(\Instr<3> ), .D(n5), .Y(n44) );
  AOI22X1 U44 ( .A(\Instr_Out<2> ), .B(n4), .C(\Instr<2> ), .D(n5), .Y(n45) );
  AOI22X1 U45 ( .A(\Instr_Out<1> ), .B(n4), .C(\Instr<1> ), .D(n5), .Y(n46) );
  AOI22X1 U46 ( .A(\Instr_Out<15> ), .B(n4), .C(\Instr<15> ), .D(n5), .Y(n47)
         );
  AOI22X1 U47 ( .A(\Instr_Out<14> ), .B(n4), .C(\Instr<14> ), .D(n5), .Y(n48)
         );
  AOI22X1 U48 ( .A(\Instr_Out<13> ), .B(n4), .C(\Instr<13> ), .D(n5), .Y(n49)
         );
  AOI22X1 U49 ( .A(\Instr_Out<12> ), .B(n4), .C(\Instr<12> ), .D(n5), .Y(n50)
         );
  NAND3X1 U50 ( .A(n9), .B(n8), .C(n51), .Y(\Instr_Muxed<11> ) );
  AOI22X1 U51 ( .A(\Instr_Out<11> ), .B(n4), .C(\Instr<11> ), .D(n5), .Y(n51)
         );
  AOI22X1 U52 ( .A(\Instr_Out<10> ), .B(n4), .C(\Instr<10> ), .D(n5), .Y(n52)
         );
  AOI22X1 U53 ( .A(\Instr_Out<0> ), .B(n4), .C(\Instr<0> ), .D(n5), .Y(n53) );
  NOR3X1 U54 ( .A(n2), .B(n6), .C(Flush), .Y(n38) );
  NOR3X1 U55 ( .A(Flush), .B(n6), .C(n75), .Y(n37) );
  AOI22X1 U56 ( .A(\IncPC<9> ), .B(n75), .C(\IncPC_Out<9> ), .D(n2), .Y(n54)
         );
  AOI22X1 U57 ( .A(\IncPC<8> ), .B(n75), .C(\IncPC_Out<8> ), .D(n3), .Y(n55)
         );
  AOI22X1 U58 ( .A(\IncPC<7> ), .B(n75), .C(\IncPC_Out<7> ), .D(n2), .Y(n56)
         );
  AOI22X1 U59 ( .A(\IncPC<6> ), .B(n75), .C(\IncPC_Out<6> ), .D(n2), .Y(n57)
         );
  AOI22X1 U60 ( .A(\IncPC<5> ), .B(n75), .C(\IncPC_Out<5> ), .D(n3), .Y(n58)
         );
  AOI22X1 U61 ( .A(\IncPC<4> ), .B(n75), .C(\IncPC_Out<4> ), .D(n2), .Y(n59)
         );
  AOI22X1 U62 ( .A(\IncPC<3> ), .B(n75), .C(\IncPC_Out<3> ), .D(n2), .Y(n60)
         );
  AOI22X1 U63 ( .A(\IncPC<2> ), .B(n75), .C(\IncPC_Out<2> ), .D(n3), .Y(n61)
         );
  AOI22X1 U64 ( .A(\IncPC<1> ), .B(n75), .C(\IncPC_Out<1> ), .D(n2), .Y(n62)
         );
  AOI22X1 U65 ( .A(\IncPC<15> ), .B(n75), .C(\IncPC_Out<15> ), .D(n2), .Y(n63)
         );
  AOI22X1 U66 ( .A(\IncPC<14> ), .B(n75), .C(\IncPC_Out<14> ), .D(n3), .Y(n64)
         );
  AOI22X1 U67 ( .A(\IncPC<13> ), .B(n75), .C(\IncPC_Out<13> ), .D(n2), .Y(n65)
         );
  AOI22X1 U68 ( .A(\IncPC<12> ), .B(n75), .C(\IncPC_Out<12> ), .D(n2), .Y(n66)
         );
  AOI22X1 U69 ( .A(\IncPC<11> ), .B(n75), .C(\IncPC_Out<11> ), .D(n3), .Y(n67)
         );
  AOI22X1 U70 ( .A(\IncPC<10> ), .B(n75), .C(\IncPC_Out<10> ), .D(n2), .Y(n68)
         );
  AOI22X1 U71 ( .A(\IncPC<0> ), .B(n75), .C(\IncPC_Out<0> ), .D(n2), .Y(n69)
         );
  dff_355 \instr_reg[0]  ( .q(\Instr_Out<0> ), .d(n32), .clk(clk), .rst(1'b0)
         );
  dff_356 \instr_reg[1]  ( .q(\Instr_Out<1> ), .d(n33), .clk(clk), .rst(1'b0)
         );
  dff_357 \instr_reg[2]  ( .q(\Instr_Out<2> ), .d(n34), .clk(clk), .rst(1'b0)
         );
  dff_358 \instr_reg[3]  ( .q(\Instr_Out<3> ), .d(n35), .clk(clk), .rst(1'b0)
         );
  dff_359 \instr_reg[4]  ( .q(\Instr_Out<4> ), .d(n70), .clk(clk), .rst(1'b0)
         );
  dff_360 \instr_reg[5]  ( .q(\Instr_Out<5> ), .d(n71), .clk(clk), .rst(1'b0)
         );
  dff_361 \instr_reg[6]  ( .q(\Instr_Out<6> ), .d(n72), .clk(clk), .rst(1'b0)
         );
  dff_362 \instr_reg[7]  ( .q(\Instr_Out<7> ), .d(n73), .clk(clk), .rst(1'b0)
         );
  dff_363 \instr_reg[8]  ( .q(\Instr_Out<8> ), .d(n31), .clk(clk), .rst(1'b0)
         );
  dff_364 \instr_reg[9]  ( .q(\Instr_Out<9> ), .d(n30), .clk(clk), .rst(1'b0)
         );
  dff_365 \instr_reg[10]  ( .q(\Instr_Out<10> ), .d(n29), .clk(clk), .rst(1'b0) );
  dff_366 \instr_reg[11]  ( .q(\Instr_Out<11> ), .d(\Instr_Muxed<11> ), .clk(
        clk), .rst(1'b0) );
  dff_367 \instr_reg[12]  ( .q(\Instr_Out<12> ), .d(n28), .clk(clk), .rst(1'b0) );
  dff_368 \instr_reg[13]  ( .q(\Instr_Out<13> ), .d(n27), .clk(clk), .rst(1'b0) );
  dff_369 \instr_reg[14]  ( .q(\Instr_Out<14> ), .d(n26), .clk(clk), .rst(1'b0) );
  dff_370 \instr_reg[15]  ( .q(\Instr_Out<15> ), .d(n25), .clk(clk), .rst(1'b0) );
  dff_339 \incpc_reg[0]  ( .q(\IncPC_Out<0> ), .d(n74), .clk(clk), .rst(n7) );
  dff_340 \incpc_reg[1]  ( .q(\IncPC_Out<1> ), .d(n24), .clk(clk), .rst(n7) );
  dff_341 \incpc_reg[2]  ( .q(\IncPC_Out<2> ), .d(n22), .clk(clk), .rst(n7) );
  dff_342 \incpc_reg[3]  ( .q(\IncPC_Out<3> ), .d(n23), .clk(clk), .rst(n6) );
  dff_343 \incpc_reg[4]  ( .q(\IncPC_Out<4> ), .d(n10), .clk(clk), .rst(n6) );
  dff_344 \incpc_reg[5]  ( .q(\IncPC_Out<5> ), .d(n11), .clk(clk), .rst(n6) );
  dff_345 \incpc_reg[6]  ( .q(\IncPC_Out<6> ), .d(n12), .clk(clk), .rst(n6) );
  dff_346 \incpc_reg[7]  ( .q(\IncPC_Out<7> ), .d(n13), .clk(clk), .rst(n6) );
  dff_347 \incpc_reg[8]  ( .q(\IncPC_Out<8> ), .d(n14), .clk(clk), .rst(n6) );
  dff_348 \incpc_reg[9]  ( .q(\IncPC_Out<9> ), .d(n15), .clk(clk), .rst(n6) );
  dff_349 \incpc_reg[10]  ( .q(\IncPC_Out<10> ), .d(n16), .clk(clk), .rst(n6)
         );
  dff_350 \incpc_reg[11]  ( .q(\IncPC_Out<11> ), .d(n17), .clk(clk), .rst(n6)
         );
  dff_351 \incpc_reg[12]  ( .q(\IncPC_Out<12> ), .d(n18), .clk(clk), .rst(n6)
         );
  dff_352 \incpc_reg[13]  ( .q(\IncPC_Out<13> ), .d(n19), .clk(clk), .rst(n6)
         );
  dff_353 \incpc_reg[14]  ( .q(\IncPC_Out<14> ), .d(n20), .clk(clk), .rst(n6)
         );
  dff_354 \incpc_reg[15]  ( .q(\IncPC_Out<15> ), .d(n21), .clk(clk), .rst(n6)
         );
  dff_371 rst_ff ( .q(CPUActive), .d(n8), .clk(clk), .rst(n6) );
  INVX1 U3 ( .A(n8), .Y(n7) );
  INVX1 U4 ( .A(n8), .Y(n6) );
  INVX1 U5 ( .A(Flush), .Y(n9) );
  INVX2 U6 ( .A(Stall), .Y(n1) );
  INVX1 U7 ( .A(rst), .Y(n8) );
  INVX2 U8 ( .A(n1), .Y(n3) );
  INVX1 U9 ( .A(n69), .Y(n74) );
  INVX1 U10 ( .A(n68), .Y(n16) );
  INVX1 U11 ( .A(n67), .Y(n17) );
  INVX1 U12 ( .A(n66), .Y(n18) );
  INVX1 U13 ( .A(n65), .Y(n19) );
  INVX1 U14 ( .A(n64), .Y(n20) );
  INVX1 U15 ( .A(n63), .Y(n21) );
  INVX1 U16 ( .A(n62), .Y(n24) );
  INVX1 U17 ( .A(n61), .Y(n22) );
  INVX1 U18 ( .A(n60), .Y(n23) );
  INVX1 U19 ( .A(n59), .Y(n10) );
  INVX1 U20 ( .A(n58), .Y(n11) );
  INVX1 U21 ( .A(n57), .Y(n12) );
  INVX1 U22 ( .A(n56), .Y(n13) );
  INVX1 U23 ( .A(n55), .Y(n14) );
  INVX1 U24 ( .A(n54), .Y(n15) );
  INVX1 U25 ( .A(n53), .Y(n32) );
  INVX1 U26 ( .A(n52), .Y(n29) );
  INVX1 U27 ( .A(n50), .Y(n28) );
  INVX1 U28 ( .A(n49), .Y(n27) );
  INVX1 U29 ( .A(n48), .Y(n26) );
  INVX1 U30 ( .A(n47), .Y(n25) );
  INVX1 U31 ( .A(n46), .Y(n33) );
  INVX1 U32 ( .A(n45), .Y(n34) );
  INVX1 U33 ( .A(n44), .Y(n35) );
  INVX1 U34 ( .A(n43), .Y(n70) );
  INVX1 U35 ( .A(n42), .Y(n71) );
  INVX1 U36 ( .A(n41), .Y(n72) );
  INVX1 U72 ( .A(n40), .Y(n73) );
  INVX1 U73 ( .A(n39), .Y(n31) );
  INVX1 U74 ( .A(n36), .Y(n30) );
  BUFX2 U75 ( .A(n37), .Y(n4) );
  BUFX2 U76 ( .A(n38), .Y(n5) );
  INVX8 U77 ( .A(n3), .Y(n75) );
  INVX8 U78 ( .A(n1), .Y(n2) );
endmodule


module decode ( clk, rst, Stall, .Instr({\Instr<15> , \Instr<14> , \Instr<13> , 
        \Instr<12> , \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , 
        \Instr<7> , \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> , 
        \Instr<1> , \Instr<0> }), .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .IncPC({\IncPC<15> , \IncPC<14> , 
        \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , 
        \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , 
        \IncPC<2> , \IncPC<1> , \IncPC<0> }), .ALUOp1({\ALUOp1<15> , 
        \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , 
        \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , 
        \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), 
    .ALUOp2({\ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , 
        \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , 
        \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , 
        \ALUOp2<1> , \ALUOp2<0> }), ALUSrc, .Immediate({\Immediate<15> , 
        \Immediate<14> , \Immediate<13> , \Immediate<12> , \Immediate<11> , 
        \Immediate<10> , \Immediate<9> , \Immediate<8> , \Immediate<7> , 
        \Immediate<6> , \Immediate<5> , \Immediate<4> , \Immediate<3> , 
        \Immediate<2> , \Immediate<1> , \Immediate<0> }), Branch, Jump, 
        JumpReg, Set, Btr, InvA, InvB, Cin, .ALUOpcode({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .Func({\Func<1> , \Func<0> }), 
        MemWrite, MemRead, MemToReg, Halt, Exception, Err, Rti, .Rs({\Rs<2> , 
        \Rs<1> , \Rs<0> }), .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({\Rd<2> , 
        \Rd<1> , \Rd<0> }), RegFileWrEn, RegFileWrEn_Out, .WriteReg({
        \WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), .WriteReg_Out({
        \WriteReg_Out<2> , \WriteReg_Out<1> , \WriteReg_Out<0> }), RtValid, 
        RsValid, RdValid, Link, Store );
  input clk, rst, Stall, \Instr<15> , \Instr<14> , \Instr<13> , \Instr<12> ,
         \Instr<11> , \Instr<10> , \Instr<9> , \Instr<8> , \Instr<7> ,
         \Instr<6> , \Instr<5> , \Instr<4> , \Instr<3> , \Instr<2> ,
         \Instr<1> , \Instr<0> , \WriteData<15> , \WriteData<14> ,
         \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> ,
         \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> ,
         \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> ,
         \WriteData<1> , \WriteData<0> , \IncPC<15> , \IncPC<14> , \IncPC<13> ,
         \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> ,
         \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> ,
         \IncPC<2> , \IncPC<1> , \IncPC<0> , RegFileWrEn, \WriteReg<2> ,
         \WriteReg<1> , \WriteReg<0> ;
  output \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> ,
         \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> ,
         \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> ,
         \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , ALUSrc, \Immediate<15> , \Immediate<14> ,
         \Immediate<13> , \Immediate<12> , \Immediate<11> , \Immediate<10> ,
         \Immediate<9> , \Immediate<8> , \Immediate<7> , \Immediate<6> ,
         \Immediate<5> , \Immediate<4> , \Immediate<3> , \Immediate<2> ,
         \Immediate<1> , \Immediate<0> , Branch, Jump, JumpReg, Set, Btr, InvA,
         InvB, Cin, \ALUOpcode<2> , \ALUOpcode<1> , \ALUOpcode<0> , \Func<1> ,
         \Func<0> , MemWrite, MemRead, MemToReg, Halt, Exception, Err, Rti,
         \Rs<2> , \Rs<1> , \Rs<0> , \Rt<2> , \Rt<1> , \Rt<0> , \Rd<2> ,
         \Rd<1> , \Rd<0> , RegFileWrEn_Out, \WriteReg_Out<2> ,
         \WriteReg_Out<1> , \WriteReg_Out<0> , RtValid, RsValid, RdValid, Link,
         Store;
  wire   Instr_15, Instr_14, Instr_13, n114, Rf, If1, If2, \rs_out<15> ,
         \rs_out<14> , \rs_out<13> , \rs_out<12> , \rs_out<11> , \rs_out<10> ,
         \rs_out<9> , \rs_out<8> , \rs_out<7> , \rs_out<6> , \rs_out<5> ,
         \rs_out<4> , \rs_out<3> , \rs_out<2> , \rs_out<1> , \rs_out<0> ,
         RfError, stu, slbi, lbi, ZeroExt, N73, N74, N75, N76, N77, N83, N84,
         n29, n30, n31, n32, n38, n42, n47, n48, n49, n55, n57, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n33, n34, n35, n36, n37, n39,
         n40, n41, n43, n44, n45, n46, n50, n51, n52, n53, n54, n56, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n81, n83, n85, n87, n92, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113;
  assign Instr_15 = \Instr<15> ;
  assign Instr_14 = \Instr<14> ;
  assign Instr_13 = \Instr<13> ;
  assign Err = 1'b0;

  LATCH \write_reg_reg<2>  ( .CLK(n26), .D(n23), .Q(\WriteReg_Out<2> ) );
  LATCH \write_reg_reg<1>  ( .CLK(n26), .D(n20), .Q(\WriteReg_Out<1> ) );
  LATCH \write_reg_reg<0>  ( .CLK(n26), .D(n17), .Q(\WriteReg_Out<0> ) );
  LATCH \ImmReg_reg<15>  ( .CLK(N83), .D(N84), .Q(\Immediate<15> ) );
  LATCH \ImmReg_reg<14>  ( .CLK(N83), .D(N84), .Q(\Immediate<14> ) );
  LATCH \ImmReg_reg<13>  ( .CLK(N83), .D(N84), .Q(\Immediate<13> ) );
  LATCH \ImmReg_reg<12>  ( .CLK(N83), .D(N84), .Q(\Immediate<12> ) );
  LATCH \ImmReg_reg<11>  ( .CLK(N83), .D(N84), .Q(\Immediate<11> ) );
  LATCH \ImmReg_reg<10>  ( .CLK(N83), .D(N84), .Q(\Immediate<10> ) );
  LATCH \ImmReg_reg<9>  ( .CLK(N83), .D(N77), .Q(\Immediate<9> ) );
  LATCH \ImmReg_reg<8>  ( .CLK(N83), .D(N76), .Q(\Immediate<8> ) );
  LATCH \ImmReg_reg<7>  ( .CLK(N83), .D(N75), .Q(\Immediate<7> ) );
  LATCH \ImmReg_reg<6>  ( .CLK(N83), .D(N74), .Q(\Immediate<6> ) );
  LATCH \ImmReg_reg<5>  ( .CLK(N83), .D(N73), .Q(\Immediate<5> ) );
  LATCH \ImmReg_reg<4>  ( .CLK(N83), .D(\Instr<4> ), .Q(\Immediate<4> ) );
  LATCH \ImmReg_reg<3>  ( .CLK(N83), .D(\Instr<3> ), .Q(\Immediate<3> ) );
  LATCH \ImmReg_reg<2>  ( .CLK(N83), .D(\Instr<2> ), .Q(\Immediate<2> ) );
  LATCH \ImmReg_reg<1>  ( .CLK(N83), .D(\Instr<1> ), .Q(\Immediate<1> ) );
  LATCH \ImmReg_reg<0>  ( .CLK(N83), .D(\Instr<0> ), .Q(\Immediate<0> ) );
  OR2X2 U3 ( .A(Instr_13), .B(Instr_14), .Y(n29) );
  OR2X2 U4 ( .A(RdValid), .B(n14), .Y(RsValid) );
  OR2X2 U5 ( .A(If1), .B(RtValid), .Y(RdValid) );
  AND2X2 U6 ( .A(Rf), .B(n31), .Y(RtValid) );
  NOR3X1 U42 ( .A(n29), .B(n113), .C(n30), .Y(Store) );
  XOR2X1 U43 ( .A(\Instr<12> ), .B(\Instr<11> ), .Y(n30) );
  NAND3X1 U44 ( .A(n110), .B(n112), .C(n32), .Y(n31) );
  NOR2X1 U45 ( .A(Instr_15), .B(Instr_14), .Y(n32) );
  OAI21X1 U46 ( .A(Rf), .B(n92), .C(n6), .Y(\Rd<2> ) );
  OAI21X1 U48 ( .A(Rf), .B(n81), .C(n12), .Y(\Rd<1> ) );
  OAI21X1 U50 ( .A(Rf), .B(n79), .C(n10), .Y(\Rd<0> ) );
  OAI21X1 U52 ( .A(Jump), .B(n68), .C(n105), .Y(N83) );
  OAI21X1 U53 ( .A(n28), .B(n94), .C(n95), .Y(N84) );
  OAI21X1 U54 ( .A(n28), .B(n85), .C(n95), .Y(N77) );
  OAI21X1 U55 ( .A(n28), .B(n83), .C(n95), .Y(N76) );
  OAI21X1 U56 ( .A(n92), .B(n76), .C(n4), .Y(n38) );
  OAI21X1 U57 ( .A(n105), .B(n92), .C(n4), .Y(N75) );
  OAI21X1 U58 ( .A(n105), .B(n81), .C(n4), .Y(N74) );
  OAI21X1 U59 ( .A(n105), .B(n79), .C(n4), .Y(N73) );
  NAND3X1 U62 ( .A(n76), .B(n28), .C(n61), .Y(n42) );
  AOI22X1 U68 ( .A(\Rs<2> ), .B(n48), .C(n49), .D(\Instr<4> ), .Y(n47) );
  AOI22X1 U73 ( .A(\Instr<9> ), .B(n48), .C(n49), .D(\Instr<3> ), .Y(n55) );
  AOI22X1 U76 ( .A(\Instr<8> ), .B(n48), .C(n49), .D(\Instr<2> ), .Y(n57) );
  NOR3X1 U77 ( .A(If1), .B(n16), .C(n109), .Y(n49) );
  OAI21X1 U78 ( .A(n73), .B(n107), .C(n66), .Y(n48) );
  OAI21X1 U85 ( .A(n78), .B(n97), .C(n58), .Y(\ALUOp1<9> ) );
  OAI21X1 U87 ( .A(n78), .B(n96), .C(n54), .Y(\ALUOp1<8> ) );
  OAI21X1 U89 ( .A(n78), .B(n103), .C(n52), .Y(\ALUOp1<15> ) );
  OAI21X1 U91 ( .A(n78), .B(n102), .C(n50), .Y(\ALUOp1<14> ) );
  OAI21X1 U93 ( .A(n78), .B(n101), .C(n45), .Y(\ALUOp1<13> ) );
  OAI21X1 U95 ( .A(n78), .B(n100), .C(n43), .Y(\ALUOp1<12> ) );
  OAI21X1 U97 ( .A(n78), .B(n99), .C(n40), .Y(\ALUOp1<11> ) );
  OAI21X1 U99 ( .A(n78), .B(n98), .C(n37), .Y(\ALUOp1<10> ) );
  rf_bypass regfile ( .read1data({\rs_out<15> , \rs_out<14> , \rs_out<13> , 
        \rs_out<12> , \rs_out<11> , \rs_out<10> , \rs_out<9> , \rs_out<8> , 
        \rs_out<7> , \rs_out<6> , \rs_out<5> , \rs_out<4> , \rs_out<3> , 
        \rs_out<2> , \rs_out<1> , \rs_out<0> }), .read2data({\ALUOp2<15> , 
        \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , 
        \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , 
        \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), 
        .err(RfError), .clk(clk), .rst(rst), .read1regsel({\Rs<2> , \Instr<9> , 
        \Instr<8> }), .read2regsel({\Rt<2> , \Instr<6> , \Instr<5> }), 
        .writeregsel({\WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), 
        .writedata({\WriteData<15> , \WriteData<14> , \WriteData<13> , 
        \WriteData<12> , \WriteData<11> , \WriteData<10> , \WriteData<9> , 
        \WriteData<8> , \WriteData<7> , \WriteData<6> , \WriteData<5> , 
        \WriteData<4> , \WriteData<3> , \WriteData<2> , \WriteData<1> , 
        \WriteData<0> }), .write(RegFileWrEn) );
  control_unit cu ( .opcode({Instr_15, Instr_14, Instr_13, \Instr<12> , 
        \Instr<11> }), .func({\Instr<1> , \Instr<0> }), .aluop({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .alusrc(ALUSrc), .branch(n114), 
        .jump(Jump), .i1(If1), .i2(If2), .r(Rf), .jumpreg(JumpReg), .set(Set), 
        .btr(Btr), .regwrite(RegFileWrEn_Out), .memwrite(MemWrite), .memread(
        MemRead), .memtoreg(MemToReg), .invA(InvA), .invB(InvB), .cin(Cin), 
        .excp(Exception), .zeroext(ZeroExt), .halt(Halt), .slbi(slbi), .link(
        Link), .lbi(lbi), .stu(stu), .rti(Rti) );
  INVX1 U7 ( .A(lbi), .Y(n104) );
  INVX1 U8 ( .A(Instr_13), .Y(n112) );
  AND2X1 U9 ( .A(\rs_out<2> ), .B(n64), .Y(\ALUOp1<2> ) );
  AND2X1 U10 ( .A(\rs_out<3> ), .B(n64), .Y(\ALUOp1<3> ) );
  AND2X1 U11 ( .A(\rs_out<4> ), .B(n64), .Y(\ALUOp1<4> ) );
  AND2X1 U12 ( .A(\rs_out<5> ), .B(n64), .Y(\ALUOp1<5> ) );
  AND2X1 U13 ( .A(\rs_out<6> ), .B(n64), .Y(\ALUOp1<6> ) );
  AND2X1 U14 ( .A(\rs_out<7> ), .B(n64), .Y(\ALUOp1<7> ) );
  INVX1 U15 ( .A(\rs_out<0> ), .Y(n96) );
  INVX1 U16 ( .A(\rs_out<1> ), .Y(n97) );
  INVX1 U17 ( .A(\rs_out<3> ), .Y(n99) );
  INVX1 U18 ( .A(\rs_out<4> ), .Y(n100) );
  INVX1 U19 ( .A(\rs_out<5> ), .Y(n101) );
  INVX1 U20 ( .A(\rs_out<6> ), .Y(n102) );
  INVX1 U21 ( .A(\rs_out<7> ), .Y(n103) );
  INVX1 U22 ( .A(\Instr<7> ), .Y(n92) );
  INVX1 U23 ( .A(\Instr<10> ), .Y(n94) );
  INVX1 U24 ( .A(Instr_15), .Y(n113) );
  INVX1 U25 ( .A(ZeroExt), .Y(n108) );
  INVX1 U26 ( .A(stu), .Y(n107) );
  AND2X1 U27 ( .A(\rs_out<0> ), .B(n64), .Y(\ALUOp1<0> ) );
  AND2X1 U28 ( .A(n64), .B(\rs_out<1> ), .Y(\ALUOp1<1> ) );
  INVX1 U29 ( .A(\rs_out<2> ), .Y(n98) );
  INVX1 U30 ( .A(n38), .Y(n95) );
  AND2X1 U31 ( .A(n72), .B(\Rt<2> ), .Y(n8) );
  AND2X1 U32 ( .A(n70), .B(n108), .Y(n75) );
  AND2X1 U33 ( .A(n72), .B(\Instr<6> ), .Y(n1) );
  AND2X1 U34 ( .A(n72), .B(\Instr<5> ), .Y(n2) );
  INVX1 U35 ( .A(\Instr<12> ), .Y(n110) );
  OR2X1 U36 ( .A(n62), .B(n7), .Y(n3) );
  INVX1 U37 ( .A(Jump), .Y(n111) );
  OR2X1 U38 ( .A(n68), .B(n3), .Y(n4) );
  AND2X2 U39 ( .A(\Instr<4> ), .B(Rf), .Y(n5) );
  INVX1 U40 ( .A(n5), .Y(n6) );
  INVX1 U41 ( .A(\Instr<4> ), .Y(n7) );
  AND2X2 U47 ( .A(\Instr<2> ), .B(Rf), .Y(n9) );
  INVX1 U49 ( .A(n9), .Y(n10) );
  AND2X2 U51 ( .A(\Instr<3> ), .B(Rf), .Y(n11) );
  INVX1 U60 ( .A(n11), .Y(n12) );
  INVX1 U61 ( .A(If2), .Y(n13) );
  INVX1 U63 ( .A(n13), .Y(n14) );
  BUFX2 U64 ( .A(n114), .Y(Branch) );
  BUFX2 U65 ( .A(n14), .Y(n16) );
  OR2X1 U66 ( .A(n2), .B(n18), .Y(n17) );
  OR2X1 U67 ( .A(n19), .B(Link), .Y(n18) );
  INVX1 U69 ( .A(n57), .Y(n19) );
  OR2X1 U70 ( .A(n1), .B(n21), .Y(n20) );
  OR2X1 U71 ( .A(n22), .B(Link), .Y(n21) );
  INVX1 U72 ( .A(n55), .Y(n22) );
  OR2X1 U74 ( .A(n8), .B(n24), .Y(n23) );
  OR2X1 U75 ( .A(n25), .B(Link), .Y(n24) );
  INVX1 U79 ( .A(n47), .Y(n25) );
  OR2X1 U80 ( .A(n74), .B(n27), .Y(n26) );
  OR2X1 U81 ( .A(n34), .B(n65), .Y(n27) );
  OR2X1 U82 ( .A(n75), .B(n33), .Y(n28) );
  OR2X1 U83 ( .A(n35), .B(n111), .Y(n33) );
  OR2X1 U84 ( .A(n49), .B(Link), .Y(n34) );
  OR2X1 U86 ( .A(ZeroExt), .B(If1), .Y(n35) );
  AND2X1 U88 ( .A(\rs_out<10> ), .B(n64), .Y(n36) );
  INVX1 U90 ( .A(n36), .Y(n37) );
  AND2X1 U92 ( .A(\rs_out<11> ), .B(n64), .Y(n39) );
  INVX1 U94 ( .A(n39), .Y(n40) );
  AND2X1 U96 ( .A(\rs_out<12> ), .B(n64), .Y(n41) );
  INVX1 U98 ( .A(n41), .Y(n43) );
  AND2X1 U100 ( .A(\rs_out<13> ), .B(n64), .Y(n44) );
  INVX1 U101 ( .A(n44), .Y(n45) );
  AND2X1 U102 ( .A(\rs_out<14> ), .B(n64), .Y(n46) );
  INVX1 U103 ( .A(n46), .Y(n50) );
  AND2X1 U104 ( .A(\rs_out<15> ), .B(n64), .Y(n51) );
  INVX1 U105 ( .A(n51), .Y(n52) );
  AND2X1 U106 ( .A(\rs_out<8> ), .B(n64), .Y(n53) );
  INVX1 U107 ( .A(n53), .Y(n54) );
  AND2X1 U108 ( .A(\rs_out<9> ), .B(n64), .Y(n56) );
  INVX1 U109 ( .A(n56), .Y(n58) );
  INVX1 U110 ( .A(n94), .Y(\Rs<2> ) );
  INVX1 U111 ( .A(n92), .Y(\Rt<2> ) );
  BUFX2 U112 ( .A(n42), .Y(n59) );
  INVX1 U113 ( .A(n59), .Y(n105) );
  AND2X1 U114 ( .A(n70), .B(n111), .Y(n60) );
  INVX1 U115 ( .A(n60), .Y(n61) );
  OR2X1 U116 ( .A(ZeroExt), .B(Jump), .Y(n62) );
  OR2X1 U117 ( .A(lbi), .B(slbi), .Y(n63) );
  INVX1 U118 ( .A(n63), .Y(n64) );
  AND2X1 U119 ( .A(n70), .B(n109), .Y(n65) );
  INVX1 U120 ( .A(n65), .Y(n66) );
  AND2X1 U121 ( .A(If1), .B(n106), .Y(n67) );
  INVX1 U122 ( .A(n67), .Y(n68) );
  OR2X1 U123 ( .A(n106), .B(If1), .Y(n69) );
  INVX1 U124 ( .A(n69), .Y(n70) );
  OR2X1 U125 ( .A(n73), .B(stu), .Y(n71) );
  INVX1 U126 ( .A(n71), .Y(n72) );
  INVX1 U127 ( .A(n74), .Y(n73) );
  AND2X1 U128 ( .A(n67), .B(n109), .Y(n74) );
  INVX1 U129 ( .A(n75), .Y(n76) );
  INVX1 U130 ( .A(n16), .Y(n106) );
  INVX1 U131 ( .A(Rf), .Y(n109) );
  AND2X1 U132 ( .A(slbi), .B(n104), .Y(n77) );
  INVX1 U133 ( .A(n77), .Y(n78) );
  INVX1 U134 ( .A(n110), .Y(\Func<1> ) );
  INVX1 U135 ( .A(n87), .Y(\Func<0> ) );
  INVX1 U136 ( .A(\Instr<11> ), .Y(n87) );
  INVX1 U137 ( .A(n85), .Y(\Rs<1> ) );
  INVX1 U138 ( .A(\Instr<9> ), .Y(n85) );
  INVX1 U139 ( .A(n83), .Y(\Rs<0> ) );
  INVX1 U140 ( .A(\Instr<8> ), .Y(n83) );
  INVX1 U141 ( .A(n81), .Y(\Rt<1> ) );
  INVX1 U142 ( .A(\Instr<6> ), .Y(n81) );
  INVX1 U143 ( .A(n79), .Y(\Rt<0> ) );
  INVX1 U144 ( .A(\Instr<5> ), .Y(n79) );
endmodule


module pipe_de ( clk, rst, Stall, Flush, .ALUOp1({\ALUOp1<15> , \ALUOp1<14> , 
        \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , 
        \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , 
        \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), .ALUOp2({
        \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , 
        \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , 
        \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , 
        \ALUOp2<0> }), .Immediate({\Immediate<15> , \Immediate<14> , 
        \Immediate<13> , \Immediate<12> , \Immediate<11> , \Immediate<10> , 
        \Immediate<9> , \Immediate<8> , \Immediate<7> , \Immediate<6> , 
        \Immediate<5> , \Immediate<4> , \Immediate<3> , \Immediate<2> , 
        \Immediate<1> , \Immediate<0> }), .ALUOpcode({\ALUOpcode<2> , 
        \ALUOpcode<1> , \ALUOpcode<0> }), .Func({\Func<1> , \Func<0> }), 
        ALUSrc, Branch, Jump, JumpReg, Set, Btr, MemWrite, MemRead, MemToReg, 
        Halt, InvA, InvB, Cin, .IncPC({\IncPC<15> , \IncPC<14> , \IncPC<13> , 
        \IncPC<12> , \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , 
        \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , 
        \IncPC<1> , \IncPC<0> }), CPUActive, .ALUOp1_Out({\ALUOp1_Out<15> , 
        \ALUOp1_Out<14> , \ALUOp1_Out<13> , \ALUOp1_Out<12> , \ALUOp1_Out<11> , 
        \ALUOp1_Out<10> , \ALUOp1_Out<9> , \ALUOp1_Out<8> , \ALUOp1_Out<7> , 
        \ALUOp1_Out<6> , \ALUOp1_Out<5> , \ALUOp1_Out<4> , \ALUOp1_Out<3> , 
        \ALUOp1_Out<2> , \ALUOp1_Out<1> , \ALUOp1_Out<0> }), .ALUOp2_Out({
        \ALUOp2_Out<15> , \ALUOp2_Out<14> , \ALUOp2_Out<13> , \ALUOp2_Out<12> , 
        \ALUOp2_Out<11> , \ALUOp2_Out<10> , \ALUOp2_Out<9> , \ALUOp2_Out<8> , 
        \ALUOp2_Out<7> , \ALUOp2_Out<6> , \ALUOp2_Out<5> , \ALUOp2_Out<4> , 
        \ALUOp2_Out<3> , \ALUOp2_Out<2> , \ALUOp2_Out<1> , \ALUOp2_Out<0> }), 
    .Immediate_Out({\Immediate_Out<15> , \Immediate_Out<14> , 
        \Immediate_Out<13> , \Immediate_Out<12> , \Immediate_Out<11> , 
        \Immediate_Out<10> , \Immediate_Out<9> , \Immediate_Out<8> , 
        \Immediate_Out<7> , \Immediate_Out<6> , \Immediate_Out<5> , 
        \Immediate_Out<4> , \Immediate_Out<3> , \Immediate_Out<2> , 
        \Immediate_Out<1> , \Immediate_Out<0> }), .ALUOpcode_Out({
        \ALUOpcode_Out<2> , \ALUOpcode_Out<1> , \ALUOpcode_Out<0> }), 
    .Func_Out({\Func_Out<1> , \Func_Out<0> }), ALUSrc_Out, Branch_Out, 
        Jump_Out, JumpReg_Out, Set_Out, Btr_Out, MemWrite_Out, MemRead_Out, 
        MemToReg_Out, Halt_Out, InvA_Out, InvB_Out, Cin_Out, .Rs({\Rs<2> , 
        \Rs<1> , \Rs<0> }), .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({\Rd<2> , 
        \Rd<1> , \Rd<0> }), .Rs_Out({\Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> }), 
    .Rt_Out({\Rt_Out<2> , \Rt_Out<1> , \Rt_Out<0> }), .Rd_Out({\Rd_Out<2> , 
        \Rd_Out<1> , \Rd_Out<0> }), RegFileWrEn, RegFileWrEn_Out, .IncPC_Out({
        \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> , \IncPC_Out<12> , 
        \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> , \IncPC_Out<8> , 
        \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> , \IncPC_Out<4> , 
        \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> , \IncPC_Out<0> }), 
    .WriteReg({\WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), .WriteReg_Out({
        \WriteReg_Out<2> , \WriteReg_Out<1> , \WriteReg_Out<0> }), RtValid, 
        RtValid_Out, CPUActive_Out, RsValid, RdValid, RsValid_Out, RdValid_Out, 
    .DecodeIncPC({\DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> , 
        \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> , 
        \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> , \DecodeIncPC<6> , 
        \DecodeIncPC<5> , \DecodeIncPC<4> , \DecodeIncPC<3> , \DecodeIncPC<2> , 
        \DecodeIncPC<1> , \DecodeIncPC<0> }), .DecodeIncPC_Out({
        \DecodeIncPC_Out<15> , \DecodeIncPC_Out<14> , \DecodeIncPC_Out<13> , 
        \DecodeIncPC_Out<12> , \DecodeIncPC_Out<11> , \DecodeIncPC_Out<10> , 
        \DecodeIncPC_Out<9> , \DecodeIncPC_Out<8> , \DecodeIncPC_Out<7> , 
        \DecodeIncPC_Out<6> , \DecodeIncPC_Out<5> , \DecodeIncPC_Out<4> , 
        \DecodeIncPC_Out<3> , \DecodeIncPC_Out<2> , \DecodeIncPC_Out<1> , 
        \DecodeIncPC_Out<0> }), Link, Link_Out );
  input clk, rst, Stall, Flush, \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> ,
         \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> ,
         \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> ,
         \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> ,
         \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> ,
         \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> ,
         \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> , \Immediate<15> ,
         \Immediate<14> , \Immediate<13> , \Immediate<12> , \Immediate<11> ,
         \Immediate<10> , \Immediate<9> , \Immediate<8> , \Immediate<7> ,
         \Immediate<6> , \Immediate<5> , \Immediate<4> , \Immediate<3> ,
         \Immediate<2> , \Immediate<1> , \Immediate<0> , \ALUOpcode<2> ,
         \ALUOpcode<1> , \ALUOpcode<0> , \Func<1> , \Func<0> , ALUSrc, Branch,
         Jump, JumpReg, Set, Btr, MemWrite, MemRead, MemToReg, Halt, InvA,
         InvB, Cin, \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> ,
         \IncPC<11> , \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> ,
         \IncPC<6> , \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> ,
         \IncPC<1> , \IncPC<0> , CPUActive, \Rs<2> , \Rs<1> , \Rs<0> , \Rt<2> ,
         \Rt<1> , \Rt<0> , \Rd<2> , \Rd<1> , \Rd<0> , RegFileWrEn,
         \WriteReg<2> , \WriteReg<1> , \WriteReg<0> , RtValid, RsValid,
         RdValid, \DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> ,
         \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> ,
         \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> ,
         \DecodeIncPC<6> , \DecodeIncPC<5> , \DecodeIncPC<4> ,
         \DecodeIncPC<3> , \DecodeIncPC<2> , \DecodeIncPC<1> ,
         \DecodeIncPC<0> , Link;
  output \ALUOp1_Out<15> , \ALUOp1_Out<14> , \ALUOp1_Out<13> ,
         \ALUOp1_Out<12> , \ALUOp1_Out<11> , \ALUOp1_Out<10> , \ALUOp1_Out<9> ,
         \ALUOp1_Out<8> , \ALUOp1_Out<7> , \ALUOp1_Out<6> , \ALUOp1_Out<5> ,
         \ALUOp1_Out<4> , \ALUOp1_Out<3> , \ALUOp1_Out<2> , \ALUOp1_Out<1> ,
         \ALUOp1_Out<0> , \ALUOp2_Out<15> , \ALUOp2_Out<14> , \ALUOp2_Out<13> ,
         \ALUOp2_Out<12> , \ALUOp2_Out<11> , \ALUOp2_Out<10> , \ALUOp2_Out<9> ,
         \ALUOp2_Out<8> , \ALUOp2_Out<7> , \ALUOp2_Out<6> , \ALUOp2_Out<5> ,
         \ALUOp2_Out<4> , \ALUOp2_Out<3> , \ALUOp2_Out<2> , \ALUOp2_Out<1> ,
         \ALUOp2_Out<0> , \Immediate_Out<15> , \Immediate_Out<14> ,
         \Immediate_Out<13> , \Immediate_Out<12> , \Immediate_Out<11> ,
         \Immediate_Out<10> , \Immediate_Out<9> , \Immediate_Out<8> ,
         \Immediate_Out<7> , \Immediate_Out<6> , \Immediate_Out<5> ,
         \Immediate_Out<4> , \Immediate_Out<3> , \Immediate_Out<2> ,
         \Immediate_Out<1> , \Immediate_Out<0> , \ALUOpcode_Out<2> ,
         \ALUOpcode_Out<1> , \ALUOpcode_Out<0> , \Func_Out<1> , \Func_Out<0> ,
         ALUSrc_Out, Branch_Out, Jump_Out, JumpReg_Out, Set_Out, Btr_Out,
         MemWrite_Out, MemRead_Out, MemToReg_Out, Halt_Out, InvA_Out, InvB_Out,
         Cin_Out, \Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> , \Rt_Out<2> ,
         \Rt_Out<1> , \Rt_Out<0> , \Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> ,
         RegFileWrEn_Out, \IncPC_Out<15> , \IncPC_Out<14> , \IncPC_Out<13> ,
         \IncPC_Out<12> , \IncPC_Out<11> , \IncPC_Out<10> , \IncPC_Out<9> ,
         \IncPC_Out<8> , \IncPC_Out<7> , \IncPC_Out<6> , \IncPC_Out<5> ,
         \IncPC_Out<4> , \IncPC_Out<3> , \IncPC_Out<2> , \IncPC_Out<1> ,
         \IncPC_Out<0> , \WriteReg_Out<2> , \WriteReg_Out<1> ,
         \WriteReg_Out<0> , RtValid_Out, CPUActive_Out, RsValid_Out,
         RdValid_Out, \DecodeIncPC_Out<15> , \DecodeIncPC_Out<14> ,
         \DecodeIncPC_Out<13> , \DecodeIncPC_Out<12> , \DecodeIncPC_Out<11> ,
         \DecodeIncPC_Out<10> , \DecodeIncPC_Out<9> , \DecodeIncPC_Out<8> ,
         \DecodeIncPC_Out<7> , \DecodeIncPC_Out<6> , \DecodeIncPC_Out<5> ,
         \DecodeIncPC_Out<4> , \DecodeIncPC_Out<3> , \DecodeIncPC_Out<2> ,
         \DecodeIncPC_Out<1> , \DecodeIncPC_Out<0> , Link_Out;
  wire   n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246;

  AOI22X1 U117 ( .A(\WriteReg<2> ), .B(n246), .C(\WriteReg_Out<2> ), .D(Stall), 
        .Y(n118) );
  AOI22X1 U118 ( .A(\WriteReg<1> ), .B(n246), .C(\WriteReg_Out<1> ), .D(Stall), 
        .Y(n119) );
  AOI22X1 U119 ( .A(\WriteReg<0> ), .B(n246), .C(\WriteReg_Out<0> ), .D(Stall), 
        .Y(n120) );
  AOI22X1 U120 ( .A(Set), .B(n246), .C(Set_Out), .D(Stall), .Y(n121) );
  AOI22X1 U121 ( .A(\Rt<2> ), .B(n246), .C(\Rt_Out<2> ), .D(Stall), .Y(n122)
         );
  AOI22X1 U122 ( .A(\Rt<1> ), .B(n246), .C(\Rt_Out<1> ), .D(Stall), .Y(n123)
         );
  AOI22X1 U123 ( .A(\Rt<0> ), .B(n246), .C(\Rt_Out<0> ), .D(Stall), .Y(n124)
         );
  AOI22X1 U124 ( .A(RtValid), .B(n246), .C(RtValid_Out), .D(Stall), .Y(n125)
         );
  AOI22X1 U125 ( .A(\Rs<2> ), .B(n246), .C(\Rs_Out<2> ), .D(Stall), .Y(n126)
         );
  AOI22X1 U126 ( .A(\Rs<1> ), .B(n246), .C(\Rs_Out<1> ), .D(Stall), .Y(n127)
         );
  AOI22X1 U127 ( .A(\Rs<0> ), .B(n246), .C(\Rs_Out<0> ), .D(Stall), .Y(n128)
         );
  AOI22X1 U128 ( .A(RsValid), .B(n246), .C(RsValid_Out), .D(Stall), .Y(n129)
         );
  AOI22X1 U129 ( .A(RegFileWrEn), .B(n246), .C(RegFileWrEn_Out), .D(Stall), 
        .Y(n130) );
  AOI22X1 U130 ( .A(\Rd<2> ), .B(n246), .C(\Rd_Out<2> ), .D(Stall), .Y(n131)
         );
  AOI22X1 U131 ( .A(\Rd<1> ), .B(n246), .C(\Rd_Out<1> ), .D(Stall), .Y(n132)
         );
  AOI22X1 U132 ( .A(\Rd<0> ), .B(n246), .C(\Rd_Out<0> ), .D(Stall), .Y(n133)
         );
  AOI22X1 U133 ( .A(RdValid), .B(n246), .C(RdValid_Out), .D(Stall), .Y(n134)
         );
  AOI22X1 U134 ( .A(MemWrite), .B(n246), .C(MemWrite_Out), .D(Stall), .Y(n135)
         );
  AOI22X1 U135 ( .A(MemToReg), .B(n246), .C(MemToReg_Out), .D(Stall), .Y(n136)
         );
  AOI22X1 U136 ( .A(MemRead), .B(n246), .C(MemRead_Out), .D(Stall), .Y(n137)
         );
  AOI22X1 U137 ( .A(Link), .B(n246), .C(n5), .D(Stall), .Y(n138) );
  AOI22X1 U138 ( .A(Jump), .B(n246), .C(Jump_Out), .D(Stall), .Y(n139) );
  AOI22X1 U139 ( .A(JumpReg), .B(n246), .C(n4), .D(Stall), .Y(n140) );
  AOI22X1 U140 ( .A(InvB), .B(n246), .C(InvB_Out), .D(Stall), .Y(n141) );
  AOI22X1 U141 ( .A(InvA), .B(n246), .C(InvA_Out), .D(Stall), .Y(n142) );
  AOI22X1 U142 ( .A(\IncPC<9> ), .B(n246), .C(\IncPC_Out<9> ), .D(Stall), .Y(
        n143) );
  AOI22X1 U143 ( .A(\IncPC<8> ), .B(n246), .C(\IncPC_Out<8> ), .D(Stall), .Y(
        n144) );
  AOI22X1 U144 ( .A(\IncPC<7> ), .B(n246), .C(\IncPC_Out<7> ), .D(Stall), .Y(
        n145) );
  AOI22X1 U145 ( .A(\IncPC<6> ), .B(n246), .C(\IncPC_Out<6> ), .D(Stall), .Y(
        n146) );
  AOI22X1 U146 ( .A(\IncPC<5> ), .B(n246), .C(\IncPC_Out<5> ), .D(Stall), .Y(
        n147) );
  AOI22X1 U147 ( .A(\IncPC<4> ), .B(n246), .C(\IncPC_Out<4> ), .D(Stall), .Y(
        n148) );
  AOI22X1 U148 ( .A(\IncPC<3> ), .B(n246), .C(\IncPC_Out<3> ), .D(Stall), .Y(
        n149) );
  AOI22X1 U149 ( .A(\IncPC<2> ), .B(n246), .C(\IncPC_Out<2> ), .D(Stall), .Y(
        n150) );
  AOI22X1 U150 ( .A(\IncPC<1> ), .B(n246), .C(\IncPC_Out<1> ), .D(Stall), .Y(
        n151) );
  AOI22X1 U151 ( .A(\IncPC<15> ), .B(n246), .C(\IncPC_Out<15> ), .D(Stall), 
        .Y(n152) );
  AOI22X1 U152 ( .A(\IncPC<14> ), .B(n246), .C(\IncPC_Out<14> ), .D(Stall), 
        .Y(n153) );
  AOI22X1 U153 ( .A(\IncPC<13> ), .B(n246), .C(\IncPC_Out<13> ), .D(Stall), 
        .Y(n154) );
  AOI22X1 U154 ( .A(\IncPC<12> ), .B(n246), .C(\IncPC_Out<12> ), .D(Stall), 
        .Y(n155) );
  AOI22X1 U155 ( .A(\IncPC<11> ), .B(n246), .C(\IncPC_Out<11> ), .D(Stall), 
        .Y(n156) );
  AOI22X1 U156 ( .A(\IncPC<10> ), .B(n246), .C(\IncPC_Out<10> ), .D(Stall), 
        .Y(n157) );
  AOI22X1 U157 ( .A(\IncPC<0> ), .B(n246), .C(\IncPC_Out<0> ), .D(Stall), .Y(
        n158) );
  AOI22X1 U158 ( .A(\Immediate<9> ), .B(n246), .C(n1), .D(Stall), .Y(n159) );
  AOI22X1 U159 ( .A(\Immediate<8> ), .B(n246), .C(\Immediate_Out<8> ), .D(
        Stall), .Y(n160) );
  AOI22X1 U160 ( .A(\Immediate<7> ), .B(n246), .C(\Immediate_Out<7> ), .D(
        Stall), .Y(n161) );
  AOI22X1 U161 ( .A(\Immediate<6> ), .B(n246), .C(\Immediate_Out<6> ), .D(
        Stall), .Y(n162) );
  AOI22X1 U162 ( .A(\Immediate<5> ), .B(n246), .C(\Immediate_Out<5> ), .D(
        Stall), .Y(n163) );
  AOI22X1 U163 ( .A(\Immediate<4> ), .B(n246), .C(\Immediate_Out<4> ), .D(
        Stall), .Y(n164) );
  AOI22X1 U164 ( .A(\Immediate<3> ), .B(n246), .C(\Immediate_Out<3> ), .D(
        Stall), .Y(n165) );
  AOI22X1 U165 ( .A(\Immediate<2> ), .B(n246), .C(\Immediate_Out<2> ), .D(
        Stall), .Y(n166) );
  AOI22X1 U166 ( .A(\Immediate<1> ), .B(n246), .C(\Immediate_Out<1> ), .D(
        Stall), .Y(n167) );
  AOI22X1 U167 ( .A(\Immediate<15> ), .B(n246), .C(\Immediate_Out<15> ), .D(
        Stall), .Y(n168) );
  AOI22X1 U168 ( .A(\Immediate<14> ), .B(n246), .C(\Immediate_Out<14> ), .D(
        Stall), .Y(n169) );
  AOI22X1 U169 ( .A(\Immediate<13> ), .B(n246), .C(\Immediate_Out<13> ), .D(
        Stall), .Y(n170) );
  AOI22X1 U170 ( .A(\Immediate<12> ), .B(n246), .C(\Immediate_Out<12> ), .D(
        Stall), .Y(n171) );
  AOI22X1 U171 ( .A(\Immediate<11> ), .B(n246), .C(\Immediate_Out<11> ), .D(
        Stall), .Y(n172) );
  AOI22X1 U172 ( .A(\Immediate<10> ), .B(n246), .C(\Immediate_Out<10> ), .D(
        Stall), .Y(n173) );
  AOI22X1 U173 ( .A(\Immediate<0> ), .B(n246), .C(\Immediate_Out<0> ), .D(
        Stall), .Y(n174) );
  AOI22X1 U174 ( .A(Halt), .B(n246), .C(Halt_Out), .D(Stall), .Y(n175) );
  AOI22X1 U175 ( .A(\Func<1> ), .B(n246), .C(\Func_Out<1> ), .D(Stall), .Y(
        n176) );
  AOI22X1 U176 ( .A(\Func<0> ), .B(n246), .C(\Func_Out<0> ), .D(Stall), .Y(
        n177) );
  AOI22X1 U177 ( .A(\DecodeIncPC<9> ), .B(n246), .C(\DecodeIncPC_Out<9> ), .D(
        Stall), .Y(n178) );
  AOI22X1 U178 ( .A(\DecodeIncPC<8> ), .B(n246), .C(\DecodeIncPC_Out<8> ), .D(
        Stall), .Y(n179) );
  AOI22X1 U179 ( .A(\DecodeIncPC<7> ), .B(n246), .C(\DecodeIncPC_Out<7> ), .D(
        Stall), .Y(n180) );
  AOI22X1 U180 ( .A(\DecodeIncPC<6> ), .B(n246), .C(\DecodeIncPC_Out<6> ), .D(
        Stall), .Y(n181) );
  AOI22X1 U181 ( .A(\DecodeIncPC<5> ), .B(n246), .C(\DecodeIncPC_Out<5> ), .D(
        Stall), .Y(n182) );
  AOI22X1 U182 ( .A(\DecodeIncPC<4> ), .B(n246), .C(\DecodeIncPC_Out<4> ), .D(
        Stall), .Y(n183) );
  AOI22X1 U183 ( .A(\DecodeIncPC<3> ), .B(n246), .C(\DecodeIncPC_Out<3> ), .D(
        Stall), .Y(n184) );
  AOI22X1 U184 ( .A(\DecodeIncPC<2> ), .B(n246), .C(\DecodeIncPC_Out<2> ), .D(
        Stall), .Y(n185) );
  AOI22X1 U185 ( .A(\DecodeIncPC<1> ), .B(n246), .C(\DecodeIncPC_Out<1> ), .D(
        Stall), .Y(n186) );
  AOI22X1 U186 ( .A(\DecodeIncPC<15> ), .B(n246), .C(\DecodeIncPC_Out<15> ), 
        .D(Stall), .Y(n187) );
  AOI22X1 U187 ( .A(\DecodeIncPC<14> ), .B(n246), .C(\DecodeIncPC_Out<14> ), 
        .D(Stall), .Y(n188) );
  AOI22X1 U188 ( .A(\DecodeIncPC<13> ), .B(n246), .C(\DecodeIncPC_Out<13> ), 
        .D(Stall), .Y(n189) );
  AOI22X1 U189 ( .A(\DecodeIncPC<12> ), .B(n246), .C(\DecodeIncPC_Out<12> ), 
        .D(Stall), .Y(n190) );
  AOI22X1 U190 ( .A(\DecodeIncPC<11> ), .B(n246), .C(\DecodeIncPC_Out<11> ), 
        .D(Stall), .Y(n191) );
  AOI22X1 U191 ( .A(\DecodeIncPC<10> ), .B(n246), .C(n2), .D(Stall), .Y(n192)
         );
  AOI22X1 U192 ( .A(\DecodeIncPC<0> ), .B(n246), .C(\DecodeIncPC_Out<0> ), .D(
        Stall), .Y(n193) );
  AOI22X1 U193 ( .A(Cin), .B(n246), .C(Cin_Out), .D(Stall), .Y(n194) );
  AOI22X1 U194 ( .A(Btr), .B(n246), .C(Btr_Out), .D(Stall), .Y(n195) );
  AOI22X1 U195 ( .A(Branch), .B(n246), .C(Branch_Out), .D(Stall), .Y(n196) );
  AOI22X1 U196 ( .A(ALUSrc), .B(n246), .C(ALUSrc_Out), .D(Stall), .Y(n197) );
  AOI22X1 U197 ( .A(\ALUOpcode<2> ), .B(n246), .C(\ALUOpcode_Out<2> ), .D(
        Stall), .Y(n198) );
  AOI22X1 U198 ( .A(\ALUOpcode<1> ), .B(n246), .C(n3), .D(Stall), .Y(n199) );
  AOI22X1 U199 ( .A(\ALUOpcode<0> ), .B(n246), .C(\ALUOpcode_Out<0> ), .D(
        Stall), .Y(n200) );
  AOI22X1 U200 ( .A(\ALUOp2<9> ), .B(n246), .C(\ALUOp2_Out<9> ), .D(Stall), 
        .Y(n201) );
  AOI22X1 U201 ( .A(\ALUOp2<8> ), .B(n246), .C(\ALUOp2_Out<8> ), .D(Stall), 
        .Y(n202) );
  AOI22X1 U202 ( .A(\ALUOp2<7> ), .B(n246), .C(\ALUOp2_Out<7> ), .D(Stall), 
        .Y(n203) );
  AOI22X1 U203 ( .A(\ALUOp2<6> ), .B(n246), .C(\ALUOp2_Out<6> ), .D(Stall), 
        .Y(n204) );
  AOI22X1 U204 ( .A(\ALUOp2<5> ), .B(n246), .C(\ALUOp2_Out<5> ), .D(Stall), 
        .Y(n205) );
  AOI22X1 U205 ( .A(\ALUOp2<4> ), .B(n246), .C(\ALUOp2_Out<4> ), .D(Stall), 
        .Y(n206) );
  AOI22X1 U206 ( .A(\ALUOp2<3> ), .B(n246), .C(\ALUOp2_Out<3> ), .D(Stall), 
        .Y(n207) );
  AOI22X1 U207 ( .A(\ALUOp2<2> ), .B(n246), .C(\ALUOp2_Out<2> ), .D(Stall), 
        .Y(n208) );
  AOI22X1 U208 ( .A(\ALUOp2<1> ), .B(n246), .C(\ALUOp2_Out<1> ), .D(Stall), 
        .Y(n209) );
  AOI22X1 U209 ( .A(\ALUOp2<15> ), .B(n246), .C(\ALUOp2_Out<15> ), .D(Stall), 
        .Y(n210) );
  AOI22X1 U210 ( .A(\ALUOp2<14> ), .B(n246), .C(\ALUOp2_Out<14> ), .D(Stall), 
        .Y(n211) );
  AOI22X1 U211 ( .A(\ALUOp2<13> ), .B(n246), .C(\ALUOp2_Out<13> ), .D(Stall), 
        .Y(n212) );
  AOI22X1 U212 ( .A(\ALUOp2<12> ), .B(n246), .C(\ALUOp2_Out<12> ), .D(Stall), 
        .Y(n213) );
  AOI22X1 U213 ( .A(\ALUOp2<11> ), .B(n246), .C(\ALUOp2_Out<11> ), .D(Stall), 
        .Y(n214) );
  AOI22X1 U214 ( .A(\ALUOp2<10> ), .B(n246), .C(\ALUOp2_Out<10> ), .D(Stall), 
        .Y(n215) );
  AOI22X1 U215 ( .A(\ALUOp2<0> ), .B(n246), .C(\ALUOp2_Out<0> ), .D(Stall), 
        .Y(n216) );
  AOI22X1 U216 ( .A(\ALUOp1<9> ), .B(n246), .C(\ALUOp1_Out<9> ), .D(Stall), 
        .Y(n217) );
  AOI22X1 U217 ( .A(\ALUOp1<8> ), .B(n246), .C(\ALUOp1_Out<8> ), .D(Stall), 
        .Y(n218) );
  AOI22X1 U218 ( .A(\ALUOp1<7> ), .B(n246), .C(\ALUOp1_Out<7> ), .D(Stall), 
        .Y(n219) );
  AOI22X1 U219 ( .A(\ALUOp1<6> ), .B(n246), .C(\ALUOp1_Out<6> ), .D(Stall), 
        .Y(n220) );
  AOI22X1 U220 ( .A(\ALUOp1<5> ), .B(n246), .C(\ALUOp1_Out<5> ), .D(Stall), 
        .Y(n221) );
  AOI22X1 U221 ( .A(\ALUOp1<4> ), .B(n246), .C(\ALUOp1_Out<4> ), .D(Stall), 
        .Y(n222) );
  AOI22X1 U222 ( .A(\ALUOp1<3> ), .B(n246), .C(\ALUOp1_Out<3> ), .D(Stall), 
        .Y(n223) );
  AOI22X1 U223 ( .A(\ALUOp1<2> ), .B(n246), .C(\ALUOp1_Out<2> ), .D(Stall), 
        .Y(n224) );
  AOI22X1 U224 ( .A(\ALUOp1<1> ), .B(n246), .C(\ALUOp1_Out<1> ), .D(Stall), 
        .Y(n225) );
  AOI22X1 U225 ( .A(\ALUOp1<15> ), .B(n246), .C(\ALUOp1_Out<15> ), .D(Stall), 
        .Y(n226) );
  AOI22X1 U226 ( .A(\ALUOp1<14> ), .B(n246), .C(\ALUOp1_Out<14> ), .D(Stall), 
        .Y(n227) );
  AOI22X1 U227 ( .A(\ALUOp1<13> ), .B(n246), .C(\ALUOp1_Out<13> ), .D(Stall), 
        .Y(n228) );
  AOI22X1 U228 ( .A(\ALUOp1<12> ), .B(n246), .C(\ALUOp1_Out<12> ), .D(Stall), 
        .Y(n229) );
  AOI22X1 U229 ( .A(\ALUOp1<11> ), .B(n246), .C(\ALUOp1_Out<11> ), .D(Stall), 
        .Y(n230) );
  AOI22X1 U230 ( .A(\ALUOp1<10> ), .B(n246), .C(\ALUOp1_Out<10> ), .D(Stall), 
        .Y(n231) );
  AOI22X1 U231 ( .A(\ALUOp1<0> ), .B(n246), .C(\ALUOp1_Out<0> ), .D(Stall), 
        .Y(n232) );
  dff_338 LinkReg ( .q(Link_Out), .d(n93), .clk(clk), .rst(n14) );
  dff_304 \DecodeIncPC_Reg[0]  ( .q(\DecodeIncPC_Out<0> ), .d(n95), .clk(clk), 
        .rst(n14) );
  dff_305 \DecodeIncPC_Reg[1]  ( .q(\DecodeIncPC_Out<1> ), .d(n96), .clk(clk), 
        .rst(n14) );
  dff_306 \DecodeIncPC_Reg[2]  ( .q(\DecodeIncPC_Out<2> ), .d(n97), .clk(clk), 
        .rst(n14) );
  dff_307 \DecodeIncPC_Reg[3]  ( .q(\DecodeIncPC_Out<3> ), .d(n98), .clk(clk), 
        .rst(n14) );
  dff_308 \DecodeIncPC_Reg[4]  ( .q(\DecodeIncPC_Out<4> ), .d(n99), .clk(clk), 
        .rst(n14) );
  dff_309 \DecodeIncPC_Reg[5]  ( .q(\DecodeIncPC_Out<5> ), .d(n100), .clk(clk), 
        .rst(n14) );
  dff_310 \DecodeIncPC_Reg[6]  ( .q(\DecodeIncPC_Out<6> ), .d(n101), .clk(clk), 
        .rst(n14) );
  dff_311 \DecodeIncPC_Reg[7]  ( .q(\DecodeIncPC_Out<7> ), .d(n102), .clk(clk), 
        .rst(n14) );
  dff_312 \DecodeIncPC_Reg[8]  ( .q(\DecodeIncPC_Out<8> ), .d(n103), .clk(clk), 
        .rst(n14) );
  dff_313 \DecodeIncPC_Reg[9]  ( .q(\DecodeIncPC_Out<9> ), .d(n104), .clk(clk), 
        .rst(n14) );
  dff_314 \DecodeIncPC_Reg[10]  ( .q(\DecodeIncPC_Out<10> ), .d(n105), .clk(
        clk), .rst(n14) );
  dff_315 \DecodeIncPC_Reg[11]  ( .q(\DecodeIncPC_Out<11> ), .d(n106), .clk(
        clk), .rst(n13) );
  dff_316 \DecodeIncPC_Reg[12]  ( .q(\DecodeIncPC_Out<12> ), .d(n107), .clk(
        clk), .rst(n13) );
  dff_317 \DecodeIncPC_Reg[13]  ( .q(\DecodeIncPC_Out<13> ), .d(n108), .clk(
        clk), .rst(n13) );
  dff_318 \DecodeIncPC_Reg[14]  ( .q(\DecodeIncPC_Out<14> ), .d(n109), .clk(
        clk), .rst(n13) );
  dff_319 \DecodeIncPC_Reg[15]  ( .q(\DecodeIncPC_Out<15> ), .d(n110), .clk(
        clk), .rst(n13) );
  dff_337 RtValid_reg ( .q(RtValid_Out), .d(n43), .clk(clk), .rst(n13) );
  dff_336 RsValid_reg ( .q(RsValid_Out), .d(n90), .clk(clk), .rst(n13) );
  dff_335 RdValid_reg ( .q(RdValid_Out), .d(n91), .clk(clk), .rst(n13) );
  dff_301 \WriteReg_reg[0]  ( .q(\WriteReg_Out<0> ), .d(n111), .clk(clk), 
        .rst(n13) );
  dff_302 \WriteReg_reg[1]  ( .q(\WriteReg_Out<1> ), .d(n112), .clk(clk), 
        .rst(n13) );
  dff_303 \WriteReg_reg[2]  ( .q(\WriteReg_Out<2> ), .d(n113), .clk(clk), 
        .rst(n13) );
  dff_285 \incpc_reg[0]  ( .q(\IncPC_Out<0> ), .d(n114), .clk(clk), .rst(n13)
         );
  dff_286 \incpc_reg[1]  ( .q(\IncPC_Out<1> ), .d(n30), .clk(clk), .rst(n13)
         );
  dff_287 \incpc_reg[2]  ( .q(\IncPC_Out<2> ), .d(n28), .clk(clk), .rst(n12)
         );
  dff_288 \incpc_reg[3]  ( .q(\IncPC_Out<3> ), .d(n29), .clk(clk), .rst(n12)
         );
  dff_289 \incpc_reg[4]  ( .q(\IncPC_Out<4> ), .d(n16), .clk(clk), .rst(n12)
         );
  dff_290 \incpc_reg[5]  ( .q(\IncPC_Out<5> ), .d(n17), .clk(clk), .rst(n12)
         );
  dff_291 \incpc_reg[6]  ( .q(\IncPC_Out<6> ), .d(n18), .clk(clk), .rst(n12)
         );
  dff_292 \incpc_reg[7]  ( .q(\IncPC_Out<7> ), .d(n19), .clk(clk), .rst(n12)
         );
  dff_293 \incpc_reg[8]  ( .q(\IncPC_Out<8> ), .d(n20), .clk(clk), .rst(n12)
         );
  dff_294 \incpc_reg[9]  ( .q(\IncPC_Out<9> ), .d(n21), .clk(clk), .rst(n12)
         );
  dff_295 \incpc_reg[10]  ( .q(\IncPC_Out<10> ), .d(n22), .clk(clk), .rst(n12)
         );
  dff_296 \incpc_reg[11]  ( .q(\IncPC_Out<11> ), .d(n23), .clk(clk), .rst(n12)
         );
  dff_297 \incpc_reg[12]  ( .q(\IncPC_Out<12> ), .d(n24), .clk(clk), .rst(n12)
         );
  dff_298 \incpc_reg[13]  ( .q(\IncPC_Out<13> ), .d(n25), .clk(clk), .rst(n12)
         );
  dff_299 \incpc_reg[14]  ( .q(\IncPC_Out<14> ), .d(n26), .clk(clk), .rst(n12)
         );
  dff_300 \incpc_reg[15]  ( .q(\IncPC_Out<15> ), .d(n27), .clk(clk), .rst(n11)
         );
  dff_334 rf_wr_en_reg ( .q(RegFileWrEn_Out), .d(n44), .clk(clk), .rst(n11) );
  dff_282 \rs_reg[0]  ( .q(\Rs_Out<0> ), .d(n87), .clk(clk), .rst(n11) );
  dff_283 \rs_reg[1]  ( .q(\Rs_Out<1> ), .d(n88), .clk(clk), .rst(n11) );
  dff_284 \rs_reg[2]  ( .q(\Rs_Out<2> ), .d(n89), .clk(clk), .rst(n11) );
  dff_279 \rt_reg[0]  ( .q(\Rt_Out<0> ), .d(n68), .clk(clk), .rst(n11) );
  dff_280 \rt_reg[1]  ( .q(\Rt_Out<1> ), .d(n69), .clk(clk), .rst(n11) );
  dff_281 \rt_reg[2]  ( .q(\Rt_Out<2> ), .d(n70), .clk(clk), .rst(n11) );
  dff_276 \rd_reg[0]  ( .q(\Rd_Out<0> ), .d(n36), .clk(clk), .rst(n11) );
  dff_277 \rd_reg[1]  ( .q(\Rd_Out<1> ), .d(n50), .clk(clk), .rst(n11) );
  dff_278 \rd_reg[2]  ( .q(\Rd_Out<2> ), .d(n51), .clk(clk), .rst(n11) );
  dff_260 \ALUOp1_reg[0]  ( .q(\ALUOp1_Out<0> ), .d(n72), .clk(clk), .rst(n11)
         );
  dff_261 \ALUOp1_reg[1]  ( .q(\ALUOp1_Out<1> ), .d(n80), .clk(clk), .rst(n11)
         );
  dff_262 \ALUOp1_reg[2]  ( .q(\ALUOp1_Out<2> ), .d(n81), .clk(clk), .rst(n10)
         );
  dff_263 \ALUOp1_reg[3]  ( .q(\ALUOp1_Out<3> ), .d(n82), .clk(clk), .rst(n10)
         );
  dff_264 \ALUOp1_reg[4]  ( .q(\ALUOp1_Out<4> ), .d(n83), .clk(clk), .rst(n10)
         );
  dff_265 \ALUOp1_reg[5]  ( .q(\ALUOp1_Out<5> ), .d(n84), .clk(clk), .rst(n10)
         );
  dff_266 \ALUOp1_reg[6]  ( .q(\ALUOp1_Out<6> ), .d(n85), .clk(clk), .rst(n10)
         );
  dff_267 \ALUOp1_reg[7]  ( .q(\ALUOp1_Out<7> ), .d(n86), .clk(clk), .rst(n10)
         );
  dff_268 \ALUOp1_reg[8]  ( .q(\ALUOp1_Out<8> ), .d(n71), .clk(clk), .rst(n10)
         );
  dff_269 \ALUOp1_reg[9]  ( .q(\ALUOp1_Out<9> ), .d(n79), .clk(clk), .rst(n10)
         );
  dff_270 \ALUOp1_reg[10]  ( .q(\ALUOp1_Out<10> ), .d(n73), .clk(clk), .rst(
        n10) );
  dff_271 \ALUOp1_reg[11]  ( .q(\ALUOp1_Out<11> ), .d(n74), .clk(clk), .rst(
        n10) );
  dff_272 \ALUOp1_reg[12]  ( .q(\ALUOp1_Out<12> ), .d(n75), .clk(clk), .rst(
        n10) );
  dff_273 \ALUOp1_reg[13]  ( .q(\ALUOp1_Out<13> ), .d(n76), .clk(clk), .rst(
        n10) );
  dff_274 \ALUOp1_reg[14]  ( .q(\ALUOp1_Out<14> ), .d(n77), .clk(clk), .rst(
        n10) );
  dff_275 \ALUOp1_reg[15]  ( .q(\ALUOp1_Out<15> ), .d(n78), .clk(clk), .rst(n9) );
  dff_244 \ALUOp2_reg[0]  ( .q(\ALUOp2_Out<0> ), .d(n52), .clk(clk), .rst(n9)
         );
  dff_245 \ALUOp2_reg[1]  ( .q(\ALUOp2_Out<1> ), .d(n59), .clk(clk), .rst(n9)
         );
  dff_246 \ALUOp2_reg[2]  ( .q(\ALUOp2_Out<2> ), .d(n60), .clk(clk), .rst(n9)
         );
  dff_247 \ALUOp2_reg[3]  ( .q(\ALUOp2_Out<3> ), .d(n61), .clk(clk), .rst(n9)
         );
  dff_248 \ALUOp2_reg[4]  ( .q(\ALUOp2_Out<4> ), .d(n62), .clk(clk), .rst(n9)
         );
  dff_249 \ALUOp2_reg[5]  ( .q(\ALUOp2_Out<5> ), .d(n63), .clk(clk), .rst(n9)
         );
  dff_250 \ALUOp2_reg[6]  ( .q(\ALUOp2_Out<6> ), .d(n64), .clk(clk), .rst(n9)
         );
  dff_251 \ALUOp2_reg[7]  ( .q(\ALUOp2_Out<7> ), .d(n65), .clk(clk), .rst(n9)
         );
  dff_252 \ALUOp2_reg[8]  ( .q(\ALUOp2_Out<8> ), .d(n66), .clk(clk), .rst(n9)
         );
  dff_253 \ALUOp2_reg[9]  ( .q(\ALUOp2_Out<9> ), .d(n67), .clk(clk), .rst(n9)
         );
  dff_254 \ALUOp2_reg[10]  ( .q(\ALUOp2_Out<10> ), .d(n53), .clk(clk), .rst(n9) );
  dff_255 \ALUOp2_reg[11]  ( .q(\ALUOp2_Out<11> ), .d(n54), .clk(clk), .rst(n9) );
  dff_256 \ALUOp2_reg[12]  ( .q(\ALUOp2_Out<12> ), .d(n55), .clk(clk), .rst(n8) );
  dff_257 \ALUOp2_reg[13]  ( .q(\ALUOp2_Out<13> ), .d(n56), .clk(clk), .rst(n8) );
  dff_258 \ALUOp2_reg[14]  ( .q(\ALUOp2_Out<14> ), .d(n57), .clk(clk), .rst(n8) );
  dff_259 \ALUOp2_reg[15]  ( .q(\ALUOp2_Out<15> ), .d(n58), .clk(clk), .rst(n8) );
  dff_228 \Immediate_reg[0]  ( .q(\Immediate_Out<0> ), .d(n115), .clk(clk), 
        .rst(n8) );
  dff_229 \Immediate_reg[1]  ( .q(\Immediate_Out<1> ), .d(n116), .clk(clk), 
        .rst(n8) );
  dff_230 \Immediate_reg[2]  ( .q(\Immediate_Out<2> ), .d(n117), .clk(clk), 
        .rst(n8) );
  dff_231 \Immediate_reg[3]  ( .q(\Immediate_Out<3> ), .d(n233), .clk(clk), 
        .rst(n8) );
  dff_232 \Immediate_reg[4]  ( .q(\Immediate_Out<4> ), .d(n234), .clk(clk), 
        .rst(n8) );
  dff_233 \Immediate_reg[5]  ( .q(\Immediate_Out<5> ), .d(n235), .clk(clk), 
        .rst(n8) );
  dff_234 \Immediate_reg[6]  ( .q(\Immediate_Out<6> ), .d(n236), .clk(clk), 
        .rst(n8) );
  dff_235 \Immediate_reg[7]  ( .q(\Immediate_Out<7> ), .d(n237), .clk(clk), 
        .rst(n8) );
  dff_236 \Immediate_reg[8]  ( .q(\Immediate_Out<8> ), .d(n238), .clk(clk), 
        .rst(n8) );
  dff_237 \Immediate_reg[9]  ( .q(\Immediate_Out<9> ), .d(n239), .clk(clk), 
        .rst(n7) );
  dff_238 \Immediate_reg[10]  ( .q(\Immediate_Out<10> ), .d(n240), .clk(clk), 
        .rst(n7) );
  dff_239 \Immediate_reg[11]  ( .q(\Immediate_Out<11> ), .d(n241), .clk(clk), 
        .rst(n7) );
  dff_240 \Immediate_reg[12]  ( .q(\Immediate_Out<12> ), .d(n242), .clk(clk), 
        .rst(n7) );
  dff_241 \Immediate_reg[13]  ( .q(\Immediate_Out<13> ), .d(n243), .clk(clk), 
        .rst(n7) );
  dff_242 \Immediate_reg[14]  ( .q(\Immediate_Out<14> ), .d(n244), .clk(clk), 
        .rst(n7) );
  dff_243 \Immediate_reg[15]  ( .q(\Immediate_Out<15> ), .d(n245), .clk(clk), 
        .rst(n7) );
  dff_225 \ALUOpcode_reg[0]  ( .q(\ALUOpcode_Out<0> ), .d(n31), .clk(clk), 
        .rst(n7) );
  dff_226 \ALUOpcode_reg[1]  ( .q(\ALUOpcode_Out<1> ), .d(n35), .clk(clk), 
        .rst(n7) );
  dff_227 \ALUOpcode_reg[2]  ( .q(\ALUOpcode_Out<2> ), .d(n92), .clk(clk), 
        .rst(n7) );
  dff_223 \Func_reg[0]  ( .q(\Func_Out<0> ), .d(n45), .clk(clk), .rst(n7) );
  dff_224 \Func_reg[1]  ( .q(\Func_Out<1> ), .d(n94), .clk(clk), .rst(n7) );
  dff_333 ALUSrc_reg ( .q(ALUSrc_Out), .d(n46), .clk(clk), .rst(n7) );
  dff_332 Branch_reg ( .q(Branch_Out), .d(n47), .clk(clk), .rst(n6) );
  dff_331 Jump_reg ( .q(Jump_Out), .d(n48), .clk(clk), .rst(n6) );
  dff_330 JumpReg_reg ( .q(JumpReg_Out), .d(n49), .clk(clk), .rst(n6) );
  dff_329 Set_reg ( .q(Set_Out), .d(n38), .clk(clk), .rst(n6) );
  dff_328 Btr_reg ( .q(Btr_Out), .d(n39), .clk(clk), .rst(n6) );
  dff_327 MemWrite_reg ( .q(MemWrite_Out), .d(n40), .clk(clk), .rst(n6) );
  dff_326 MemRead_reg ( .q(MemRead_Out), .d(n41), .clk(clk), .rst(n6) );
  dff_325 MemToReg_reg ( .q(MemToReg_Out), .d(n42), .clk(clk), .rst(n6) );
  dff_324 Halt_reg ( .q(Halt_Out), .d(n37), .clk(clk), .rst(n6) );
  dff_323 InvA_reg ( .q(InvA_Out), .d(n33), .clk(clk), .rst(n6) );
  dff_322 InvB_reg ( .q(InvB_Out), .d(n32), .clk(clk), .rst(n6) );
  dff_321 Cin_reg ( .q(Cin_Out), .d(n34), .clk(clk), .rst(n6) );
  dff_320 CPUActive_reg ( .q(CPUActive_Out), .d(CPUActive), .clk(clk), .rst(n6) );
  INVX1 U1 ( .A(n232), .Y(n72) );
  INVX1 U2 ( .A(n225), .Y(n80) );
  INVX1 U3 ( .A(n137), .Y(n41) );
  INVX1 U4 ( .A(n136), .Y(n42) );
  INVX1 U5 ( .A(n125), .Y(n43) );
  INVX1 U6 ( .A(n224), .Y(n81) );
  INVX1 U7 ( .A(n223), .Y(n82) );
  INVX1 U8 ( .A(n222), .Y(n83) );
  INVX1 U9 ( .A(n221), .Y(n84) );
  INVX1 U10 ( .A(n220), .Y(n85) );
  INVX1 U11 ( .A(n219), .Y(n86) );
  INVX1 U12 ( .A(n177), .Y(n45) );
  INVX1 U13 ( .A(n139), .Y(n48) );
  INVX1 U14 ( .A(n140), .Y(n49) );
  INVX1 U15 ( .A(n121), .Y(n38) );
  INVX1 U16 ( .A(n195), .Y(n39) );
  INVX1 U17 ( .A(n142), .Y(n33) );
  INVX1 U18 ( .A(n141), .Y(n32) );
  INVX1 U19 ( .A(n194), .Y(n34) );
  INVX1 U20 ( .A(rst), .Y(n15) );
  BUFX2 U21 ( .A(\Immediate_Out<9> ), .Y(n1) );
  BUFX2 U22 ( .A(\DecodeIncPC_Out<10> ), .Y(n2) );
  INVX1 U23 ( .A(n138), .Y(n93) );
  INVX1 U24 ( .A(n134), .Y(n91) );
  INVX1 U25 ( .A(n15), .Y(n6) );
  INVX1 U26 ( .A(n15), .Y(n7) );
  INVX1 U27 ( .A(n15), .Y(n8) );
  INVX1 U28 ( .A(n15), .Y(n9) );
  INVX1 U29 ( .A(n15), .Y(n10) );
  INVX1 U30 ( .A(n15), .Y(n11) );
  INVX1 U31 ( .A(n15), .Y(n12) );
  INVX1 U32 ( .A(n15), .Y(n13) );
  INVX1 U33 ( .A(n15), .Y(n14) );
  INVX1 U34 ( .A(n231), .Y(n73) );
  INVX1 U35 ( .A(n230), .Y(n74) );
  INVX1 U36 ( .A(n229), .Y(n75) );
  INVX1 U37 ( .A(n228), .Y(n76) );
  INVX1 U38 ( .A(n227), .Y(n77) );
  INVX1 U39 ( .A(n226), .Y(n78) );
  INVX1 U40 ( .A(n218), .Y(n71) );
  INVX1 U41 ( .A(n217), .Y(n79) );
  INVX1 U42 ( .A(n216), .Y(n52) );
  INVX1 U43 ( .A(n215), .Y(n53) );
  INVX1 U44 ( .A(n214), .Y(n54) );
  INVX1 U45 ( .A(n213), .Y(n55) );
  INVX1 U46 ( .A(n212), .Y(n56) );
  INVX1 U47 ( .A(n211), .Y(n57) );
  INVX1 U48 ( .A(n210), .Y(n58) );
  INVX1 U49 ( .A(n209), .Y(n59) );
  INVX1 U50 ( .A(n208), .Y(n60) );
  INVX1 U51 ( .A(n207), .Y(n61) );
  INVX1 U52 ( .A(n206), .Y(n62) );
  INVX1 U53 ( .A(n205), .Y(n63) );
  INVX1 U54 ( .A(n204), .Y(n64) );
  INVX1 U55 ( .A(n203), .Y(n65) );
  INVX1 U56 ( .A(n202), .Y(n66) );
  INVX1 U57 ( .A(n201), .Y(n67) );
  INVX1 U58 ( .A(n200), .Y(n31) );
  INVX1 U59 ( .A(n199), .Y(n35) );
  INVX1 U60 ( .A(n198), .Y(n92) );
  INVX1 U61 ( .A(n197), .Y(n46) );
  INVX1 U62 ( .A(n196), .Y(n47) );
  INVX1 U63 ( .A(n193), .Y(n95) );
  INVX1 U64 ( .A(n192), .Y(n105) );
  INVX1 U65 ( .A(n191), .Y(n106) );
  INVX1 U66 ( .A(n190), .Y(n107) );
  INVX1 U67 ( .A(n189), .Y(n108) );
  INVX1 U68 ( .A(n188), .Y(n109) );
  INVX1 U69 ( .A(n187), .Y(n110) );
  INVX1 U70 ( .A(n186), .Y(n96) );
  INVX1 U71 ( .A(n185), .Y(n97) );
  INVX1 U72 ( .A(n184), .Y(n98) );
  INVX1 U73 ( .A(n183), .Y(n99) );
  INVX1 U74 ( .A(n182), .Y(n100) );
  INVX1 U75 ( .A(n181), .Y(n101) );
  INVX1 U76 ( .A(n180), .Y(n102) );
  INVX1 U77 ( .A(n179), .Y(n103) );
  INVX1 U78 ( .A(n178), .Y(n104) );
  INVX1 U79 ( .A(n176), .Y(n94) );
  INVX1 U80 ( .A(n175), .Y(n37) );
  INVX1 U81 ( .A(n174), .Y(n115) );
  INVX1 U82 ( .A(n173), .Y(n240) );
  INVX1 U83 ( .A(n172), .Y(n241) );
  INVX1 U84 ( .A(n171), .Y(n242) );
  INVX1 U85 ( .A(n170), .Y(n243) );
  INVX1 U86 ( .A(n169), .Y(n244) );
  INVX1 U87 ( .A(n168), .Y(n245) );
  INVX1 U88 ( .A(n167), .Y(n116) );
  INVX1 U89 ( .A(n166), .Y(n117) );
  INVX1 U90 ( .A(n165), .Y(n233) );
  INVX1 U91 ( .A(n164), .Y(n234) );
  INVX1 U92 ( .A(n163), .Y(n235) );
  INVX1 U93 ( .A(n162), .Y(n236) );
  INVX1 U94 ( .A(n161), .Y(n237) );
  INVX1 U95 ( .A(n160), .Y(n238) );
  INVX1 U96 ( .A(n159), .Y(n239) );
  INVX1 U97 ( .A(n158), .Y(n114) );
  INVX1 U98 ( .A(n157), .Y(n22) );
  INVX1 U99 ( .A(n156), .Y(n23) );
  INVX1 U100 ( .A(n155), .Y(n24) );
  INVX1 U101 ( .A(n154), .Y(n25) );
  INVX1 U102 ( .A(n153), .Y(n26) );
  INVX1 U103 ( .A(n152), .Y(n27) );
  INVX1 U104 ( .A(n151), .Y(n30) );
  INVX1 U105 ( .A(n150), .Y(n28) );
  INVX1 U106 ( .A(n149), .Y(n29) );
  INVX1 U107 ( .A(n148), .Y(n16) );
  INVX1 U108 ( .A(n147), .Y(n17) );
  INVX1 U109 ( .A(n146), .Y(n18) );
  INVX1 U110 ( .A(n145), .Y(n19) );
  INVX1 U111 ( .A(n144), .Y(n20) );
  INVX1 U112 ( .A(n143), .Y(n21) );
  INVX1 U113 ( .A(n135), .Y(n40) );
  INVX1 U114 ( .A(n133), .Y(n36) );
  INVX1 U115 ( .A(n132), .Y(n50) );
  INVX1 U116 ( .A(n131), .Y(n51) );
  INVX1 U232 ( .A(n130), .Y(n44) );
  INVX1 U233 ( .A(n129), .Y(n90) );
  INVX1 U234 ( .A(n128), .Y(n87) );
  INVX1 U235 ( .A(n127), .Y(n88) );
  INVX1 U236 ( .A(n126), .Y(n89) );
  INVX1 U237 ( .A(n124), .Y(n68) );
  INVX1 U238 ( .A(n123), .Y(n69) );
  INVX1 U239 ( .A(n122), .Y(n70) );
  INVX1 U240 ( .A(n120), .Y(n111) );
  INVX1 U241 ( .A(n119), .Y(n112) );
  INVX1 U242 ( .A(n118), .Y(n113) );
  BUFX2 U243 ( .A(\ALUOpcode_Out<1> ), .Y(n3) );
  BUFX2 U244 ( .A(JumpReg_Out), .Y(n4) );
  BUFX2 U245 ( .A(Link_Out), .Y(n5) );
  INVX2 U246 ( .A(Stall), .Y(n246) );
endmodule


module execute ( .ALUOp1({\ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , 
        \ALUOp1<12> , \ALUOp1<11> , \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , 
        \ALUOp1<7> , \ALUOp1<6> , \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , 
        \ALUOp1<2> , \ALUOp1<1> , \ALUOp1<0> }), .ALUOp2({\ALUOp2<15> , 
        \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , 
        \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , 
        \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), 
    .Opcode({\Opcode<2> , \Opcode<1> , \Opcode<0> }), .IncPC({\IncPC<15> , 
        \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> , \IncPC<10> , 
        \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> , \IncPC<5> , \IncPC<4> , 
        \IncPC<3> , \IncPC<2> , \IncPC<1> , \IncPC<0> }), Jump, Branch, 
        JumpReg, Set, InvA, InvB, Cin, Btr, .Func({\Func<1> , \Func<0> }), 
    .Imm({\Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> , \Imm<11> , \Imm<10> , 
        \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> , \Imm<5> , \Imm<4> , \Imm<3> , 
        \Imm<2> , \Imm<1> , \Imm<0> }), ALUSrc, .Result({\Result<15> , 
        \Result<14> , \Result<13> , \Result<12> , \Result<11> , \Result<10> , 
        \Result<9> , \Result<8> , \Result<7> , \Result<6> , \Result<5> , 
        \Result<4> , \Result<3> , \Result<2> , \Result<1> , \Result<0> }), 
    .NextPC({\NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> , 
        \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> , 
        \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> , 
        \NextPC<1> , \NextPC<0> }), Err, BranchJumpTaken, rst, .DecodeIncPC({
        \DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> , 
        \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> , 
        \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> , \DecodeIncPC<6> , 
        \DecodeIncPC<5> , \DecodeIncPC<4> , \DecodeIncPC<3> , \DecodeIncPC<2> , 
        \DecodeIncPC<1> , \DecodeIncPC<0> }), Link, .ForwardALUOp1({
        \ForwardALUOp1<1> , \ForwardALUOp1<0> }), .ForwardALUOp2({
        \ForwardALUOp2<1> , \ForwardALUOp2<0> }), .PipeMW_Result({
        \PipeMW_Result<15> , \PipeMW_Result<14> , \PipeMW_Result<13> , 
        \PipeMW_Result<12> , \PipeMW_Result<11> , \PipeMW_Result<10> , 
        \PipeMW_Result<9> , \PipeMW_Result<8> , \PipeMW_Result<7> , 
        \PipeMW_Result<6> , \PipeMW_Result<5> , \PipeMW_Result<4> , 
        \PipeMW_Result<3> , \PipeMW_Result<2> , \PipeMW_Result<1> , 
        \PipeMW_Result<0> }), .PipeEM_Result({\PipeEM_Result<15> , 
        \PipeEM_Result<14> , \PipeEM_Result<13> , \PipeEM_Result<12> , 
        \PipeEM_Result<11> , \PipeEM_Result<10> , \PipeEM_Result<9> , 
        \PipeEM_Result<8> , \PipeEM_Result<7> , \PipeEM_Result<6> , 
        \PipeEM_Result<5> , \PipeEM_Result<4> , \PipeEM_Result<3> , 
        \PipeEM_Result<2> , \PipeEM_Result<1> , \PipeEM_Result<0> }) );
  input \ALUOp1<15> , \ALUOp1<14> , \ALUOp1<13> , \ALUOp1<12> , \ALUOp1<11> ,
         \ALUOp1<10> , \ALUOp1<9> , \ALUOp1<8> , \ALUOp1<7> , \ALUOp1<6> ,
         \ALUOp1<5> , \ALUOp1<4> , \ALUOp1<3> , \ALUOp1<2> , \ALUOp1<1> ,
         \ALUOp1<0> , \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , \Opcode<2> , \Opcode<1> , \Opcode<0> ,
         \IncPC<15> , \IncPC<14> , \IncPC<13> , \IncPC<12> , \IncPC<11> ,
         \IncPC<10> , \IncPC<9> , \IncPC<8> , \IncPC<7> , \IncPC<6> ,
         \IncPC<5> , \IncPC<4> , \IncPC<3> , \IncPC<2> , \IncPC<1> ,
         \IncPC<0> , Jump, Branch, JumpReg, Set, InvA, InvB, Cin, Btr,
         \Func<1> , \Func<0> , \Imm<15> , \Imm<14> , \Imm<13> , \Imm<12> ,
         \Imm<11> , \Imm<10> , \Imm<9> , \Imm<8> , \Imm<7> , \Imm<6> ,
         \Imm<5> , \Imm<4> , \Imm<3> , \Imm<2> , \Imm<1> , \Imm<0> , ALUSrc,
         rst, \DecodeIncPC<15> , \DecodeIncPC<14> , \DecodeIncPC<13> ,
         \DecodeIncPC<12> , \DecodeIncPC<11> , \DecodeIncPC<10> ,
         \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> ,
         \DecodeIncPC<6> , \DecodeIncPC<5> , \DecodeIncPC<4> ,
         \DecodeIncPC<3> , \DecodeIncPC<2> , \DecodeIncPC<1> ,
         \DecodeIncPC<0> , Link, \ForwardALUOp1<1> , \ForwardALUOp1<0> ,
         \ForwardALUOp2<1> , \ForwardALUOp2<0> , \PipeMW_Result<15> ,
         \PipeMW_Result<14> , \PipeMW_Result<13> , \PipeMW_Result<12> ,
         \PipeMW_Result<11> , \PipeMW_Result<10> , \PipeMW_Result<9> ,
         \PipeMW_Result<8> , \PipeMW_Result<7> , \PipeMW_Result<6> ,
         \PipeMW_Result<5> , \PipeMW_Result<4> , \PipeMW_Result<3> ,
         \PipeMW_Result<2> , \PipeMW_Result<1> , \PipeMW_Result<0> ,
         \PipeEM_Result<15> , \PipeEM_Result<14> , \PipeEM_Result<13> ,
         \PipeEM_Result<12> , \PipeEM_Result<11> , \PipeEM_Result<10> ,
         \PipeEM_Result<9> , \PipeEM_Result<8> , \PipeEM_Result<7> ,
         \PipeEM_Result<6> , \PipeEM_Result<5> , \PipeEM_Result<4> ,
         \PipeEM_Result<3> , \PipeEM_Result<2> , \PipeEM_Result<1> ,
         \PipeEM_Result<0> ;
  output \Result<15> , \Result<14> , \Result<13> , \Result<12> , \Result<11> ,
         \Result<10> , \Result<9> , \Result<8> , \Result<7> , \Result<6> ,
         \Result<5> , \Result<4> , \Result<3> , \Result<2> , \Result<1> ,
         \Result<0> , \NextPC<15> , \NextPC<14> , \NextPC<13> , \NextPC<12> ,
         \NextPC<11> , \NextPC<10> , \NextPC<9> , \NextPC<8> , \NextPC<7> ,
         \NextPC<6> , \NextPC<5> , \NextPC<4> , \NextPC<3> , \NextPC<2> ,
         \NextPC<1> , \NextPC<0> , Err, BranchJumpTaken;
  wire   n504, n505, n506, n507, \alu_operand_b<15> , \alu_operand_b<14> ,
         \alu_operand_b<13> , \alu_operand_b<12> , \alu_operand_b<11> ,
         \alu_operand_b<8> , \aluResult<15> , \aluResult<14> , \aluResult<13> ,
         \aluResult<12> , \aluResult<11> , \aluResult<10> , \aluResult<9> ,
         \aluResult<8> , \aluResult<7> , \aluResult<6> , \aluResult<5> ,
         \aluResult<4> , \aluResult<3> , \aluResult<2> , \aluResult<1> ,
         \aluResult<0> , Zero, cout, \OpAReg<15> , \OpAReg<14> , \OpAReg<13> ,
         \OpAReg<12> , \OpAReg<11> , \OpAReg<10> , \OpAReg<9> , \OpAReg<8> ,
         \OpAReg<7> , \OpAReg<6> , \OpAReg<5> , \OpAReg<4> , \OpAReg<3> ,
         \OpAReg<2> , \OpAReg<1> , \OpAReg<0> , \OpBReg<15> , \OpBReg<14> ,
         \OpBReg<13> , \OpBReg<12> , \OpBReg<11> , \OpBReg<10> , \OpBReg<9> ,
         \OpBReg<8> , \OpBReg<7> , \OpBReg<6> , \OpBReg<5> , \OpBReg<4> ,
         \OpBReg<3> , \OpBReg<2> , \OpBReg<1> , \OpBReg<0> , N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N54,
         \_2_net_<0> , \setResult<15> , \setResult<14> , \setResult<13> ,
         \setResult<12> , \setResult<11> , \setResult<10> , \setResult<9> ,
         \setResult<8> , \setResult<7> , \setResult<6> , \setResult<5> ,
         \setResult<4> , \setResult<3> , \setResult<2> , \setResult<1> ,
         \setResult<0> , \offsetAddr<15> , \offsetAddr<14> , \offsetAddr<13> ,
         \offsetAddr<12> , \offsetAddr<11> , \offsetAddr<10> , \offsetAddr<9> ,
         \offsetAddr<8> , \offsetAddr<7> , \offsetAddr<6> , \offsetAddr<5> ,
         \offsetAddr<4> , \offsetAddr<3> , \offsetAddr<2> , \offsetAddr<1> ,
         \offsetAddr<0> , branch_en, _7_net_, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n113, n114, n146, n147, n148, n149, n150, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n185, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n80, n82, n93, n95, n97, n99, n101, n103,
         n105, n107, n109, n111, n115, n117, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n144, n145, n151,
         n152, n153, n184, n186, n187, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503;
  assign Err = 1'b0;

  LATCH \OpAReg_reg<15>  ( .CLK(n292), .D(N54), .Q(\OpAReg<15> ) );
  LATCH \OpAReg_reg<14>  ( .CLK(n292), .D(N52), .Q(\OpAReg<14> ) );
  LATCH \OpAReg_reg<13>  ( .CLK(n292), .D(N51), .Q(\OpAReg<13> ) );
  LATCH \OpAReg_reg<12>  ( .CLK(n292), .D(N50), .Q(\OpAReg<12> ) );
  LATCH \OpAReg_reg<11>  ( .CLK(n292), .D(N49), .Q(\OpAReg<11> ) );
  LATCH \OpAReg_reg<10>  ( .CLK(n292), .D(N48), .Q(\OpAReg<10> ) );
  LATCH \OpAReg_reg<9>  ( .CLK(n292), .D(N47), .Q(\OpAReg<9> ) );
  LATCH \OpAReg_reg<8>  ( .CLK(n292), .D(N46), .Q(\OpAReg<8> ) );
  LATCH \OpAReg_reg<7>  ( .CLK(n292), .D(N45), .Q(\OpAReg<7> ) );
  LATCH \OpAReg_reg<6>  ( .CLK(n292), .D(N44), .Q(\OpAReg<6> ) );
  LATCH \OpAReg_reg<5>  ( .CLK(n292), .D(N43), .Q(\OpAReg<5> ) );
  LATCH \OpAReg_reg<4>  ( .CLK(n292), .D(N42), .Q(\OpAReg<4> ) );
  LATCH \OpAReg_reg<3>  ( .CLK(n292), .D(N41), .Q(\OpAReg<3> ) );
  LATCH \OpAReg_reg<2>  ( .CLK(n292), .D(N40), .Q(\OpAReg<2> ) );
  LATCH \OpAReg_reg<1>  ( .CLK(n292), .D(N39), .Q(\OpAReg<1> ) );
  LATCH \OpAReg_reg<0>  ( .CLK(n292), .D(N38), .Q(\OpAReg<0> ) );
  LATCH \OpBReg_reg<15>  ( .CLK(n294), .D(n291), .Q(\OpBReg<15> ) );
  LATCH \OpBReg_reg<14>  ( .CLK(n294), .D(n289), .Q(\OpBReg<14> ) );
  LATCH \OpBReg_reg<13>  ( .CLK(n294), .D(n287), .Q(\OpBReg<13> ) );
  LATCH \OpBReg_reg<12>  ( .CLK(n294), .D(n285), .Q(\OpBReg<12> ) );
  LATCH \OpBReg_reg<11>  ( .CLK(n294), .D(n283), .Q(\OpBReg<11> ) );
  LATCH \OpBReg_reg<10>  ( .CLK(n294), .D(n281), .Q(\OpBReg<10> ) );
  LATCH \OpBReg_reg<9>  ( .CLK(n294), .D(n279), .Q(\OpBReg<9> ) );
  LATCH \OpBReg_reg<8>  ( .CLK(n294), .D(n277), .Q(\OpBReg<8> ) );
  LATCH \OpBReg_reg<7>  ( .CLK(n294), .D(n275), .Q(\OpBReg<7> ) );
  LATCH \OpBReg_reg<6>  ( .CLK(n294), .D(n273), .Q(\OpBReg<6> ) );
  LATCH \OpBReg_reg<5>  ( .CLK(n294), .D(n271), .Q(\OpBReg<5> ) );
  LATCH \OpBReg_reg<4>  ( .CLK(n294), .D(n269), .Q(\OpBReg<4> ) );
  LATCH \OpBReg_reg<3>  ( .CLK(n294), .D(n267), .Q(\OpBReg<3> ) );
  LATCH \OpBReg_reg<2>  ( .CLK(n294), .D(n265), .Q(\OpBReg<2> ) );
  LATCH \OpBReg_reg<1>  ( .CLK(n294), .D(n263), .Q(\OpBReg<1> ) );
  LATCH \OpBReg_reg<0>  ( .CLK(n294), .D(n261), .Q(\OpBReg<0> ) );
  AND2X2 U20 ( .A(n493), .B(n492), .Y(n89) );
  NAND3X1 U120 ( .A(n83), .B(n84), .C(n85), .Y(_7_net_) );
  NOR3X1 U121 ( .A(n86), .B(n87), .C(n88), .Y(n85) );
  NAND2X1 U122 ( .A(n486), .B(n487), .Y(n88) );
  NAND2X1 U123 ( .A(n488), .B(n489), .Y(n87) );
  NAND3X1 U124 ( .A(n490), .B(n491), .C(n89), .Y(n86) );
  NOR3X1 U125 ( .A(n90), .B(\ALUOp1<1> ), .C(\ALUOp1<15> ), .Y(n84) );
  NAND2X1 U126 ( .A(n497), .B(n498), .Y(n90) );
  NOR3X1 U127 ( .A(n91), .B(\ALUOp1<10> ), .C(\ALUOp1<0> ), .Y(n83) );
  NAND2X1 U128 ( .A(n495), .B(n496), .Y(n91) );
  AOI22X1 U158 ( .A(\setResult<1> ), .B(n480), .C(\ALUOp1<14> ), .D(Btr), .Y(
        n113) );
  AOI22X1 U216 ( .A(n379), .B(\ALUOp2<15> ), .C(n150), .D(\Imm<15> ), .Y(n148)
         );
  AOI22X1 U217 ( .A(\PipeEM_Result<15> ), .B(n354), .C(\PipeMW_Result<15> ), 
        .D(n355), .Y(n147) );
  AOI22X1 U220 ( .A(\ALUOp2<14> ), .B(n379), .C(n150), .D(\Imm<14> ), .Y(n155)
         );
  AOI22X1 U221 ( .A(\PipeEM_Result<14> ), .B(n354), .C(\PipeMW_Result<14> ), 
        .D(n355), .Y(n154) );
  AOI22X1 U223 ( .A(\ALUOp2<13> ), .B(n379), .C(n150), .D(\Imm<13> ), .Y(n157)
         );
  AOI22X1 U224 ( .A(\PipeEM_Result<13> ), .B(n354), .C(\PipeMW_Result<13> ), 
        .D(n355), .Y(n156) );
  AOI22X1 U226 ( .A(\ALUOp2<12> ), .B(n379), .C(n150), .D(\Imm<12> ), .Y(n159)
         );
  AOI22X1 U227 ( .A(\PipeEM_Result<12> ), .B(n354), .C(\PipeMW_Result<12> ), 
        .D(n355), .Y(n158) );
  AOI22X1 U229 ( .A(\ALUOp2<11> ), .B(n379), .C(n150), .D(\Imm<11> ), .Y(n161)
         );
  AOI22X1 U230 ( .A(\PipeEM_Result<11> ), .B(n354), .C(\PipeMW_Result<11> ), 
        .D(n355), .Y(n160) );
  AOI22X1 U232 ( .A(\ALUOp2<10> ), .B(n379), .C(n150), .D(\Imm<10> ), .Y(n163)
         );
  AOI22X1 U233 ( .A(\PipeEM_Result<10> ), .B(n354), .C(\PipeMW_Result<10> ), 
        .D(n355), .Y(n162) );
  AOI22X1 U235 ( .A(\ALUOp2<9> ), .B(n379), .C(n150), .D(\Imm<9> ), .Y(n165)
         );
  AOI22X1 U236 ( .A(\PipeEM_Result<9> ), .B(n354), .C(\PipeMW_Result<9> ), .D(
        n355), .Y(n164) );
  AOI22X1 U238 ( .A(\ALUOp2<8> ), .B(n379), .C(n150), .D(\Imm<8> ), .Y(n167)
         );
  AOI22X1 U239 ( .A(\PipeEM_Result<8> ), .B(n354), .C(\PipeMW_Result<8> ), .D(
        n355), .Y(n166) );
  AOI22X1 U241 ( .A(\ALUOp2<7> ), .B(n379), .C(n150), .D(\Imm<7> ), .Y(n169)
         );
  AOI22X1 U242 ( .A(\PipeEM_Result<7> ), .B(n354), .C(\PipeMW_Result<7> ), .D(
        n355), .Y(n168) );
  AOI22X1 U244 ( .A(\ALUOp2<6> ), .B(n379), .C(n150), .D(\Imm<6> ), .Y(n171)
         );
  AOI22X1 U245 ( .A(\PipeEM_Result<6> ), .B(n354), .C(\PipeMW_Result<6> ), .D(
        n355), .Y(n170) );
  AOI22X1 U247 ( .A(\ALUOp2<5> ), .B(n379), .C(n150), .D(\Imm<5> ), .Y(n173)
         );
  AOI22X1 U248 ( .A(\PipeEM_Result<5> ), .B(n354), .C(\PipeMW_Result<5> ), .D(
        n355), .Y(n172) );
  AOI22X1 U250 ( .A(\ALUOp2<4> ), .B(n379), .C(n150), .D(\Imm<4> ), .Y(n175)
         );
  AOI22X1 U251 ( .A(\PipeEM_Result<4> ), .B(n354), .C(\PipeMW_Result<4> ), .D(
        n355), .Y(n174) );
  AOI22X1 U253 ( .A(\ALUOp2<3> ), .B(n379), .C(n150), .D(\Imm<3> ), .Y(n177)
         );
  AOI22X1 U254 ( .A(\PipeEM_Result<3> ), .B(n354), .C(\PipeMW_Result<3> ), .D(
        n355), .Y(n176) );
  AOI22X1 U256 ( .A(\ALUOp2<2> ), .B(n379), .C(n150), .D(\Imm<2> ), .Y(n179)
         );
  AOI22X1 U257 ( .A(\PipeEM_Result<2> ), .B(n354), .C(\PipeMW_Result<2> ), .D(
        n355), .Y(n178) );
  AOI22X1 U259 ( .A(\ALUOp2<1> ), .B(n379), .C(n150), .D(\Imm<1> ), .Y(n181)
         );
  AOI22X1 U260 ( .A(\PipeEM_Result<1> ), .B(n354), .C(\PipeMW_Result<1> ), .D(
        n355), .Y(n180) );
  AOI22X1 U262 ( .A(\ALUOp2<0> ), .B(n379), .C(n150), .D(\Imm<0> ), .Y(n183)
         );
  NOR2X1 U263 ( .A(n357), .B(ALUSrc), .Y(n149) );
  AOI22X1 U265 ( .A(\PipeEM_Result<0> ), .B(n354), .C(\PipeMW_Result<0> ), .D(
        n355), .Y(n182) );
  OAI21X1 U268 ( .A(n499), .B(n378), .C(n185), .Y(N54) );
  AOI22X1 U269 ( .A(n352), .B(\PipeEM_Result<15> ), .C(n353), .D(
        \PipeMW_Result<15> ), .Y(n185) );
  OAI21X1 U271 ( .A(n498), .B(n378), .C(n188), .Y(N52) );
  AOI22X1 U272 ( .A(n352), .B(\PipeEM_Result<14> ), .C(n353), .D(
        \PipeMW_Result<14> ), .Y(n188) );
  OAI21X1 U273 ( .A(n497), .B(n378), .C(n189), .Y(N51) );
  AOI22X1 U274 ( .A(n352), .B(\PipeEM_Result<13> ), .C(n353), .D(
        \PipeMW_Result<13> ), .Y(n189) );
  OAI21X1 U275 ( .A(n496), .B(n378), .C(n190), .Y(N50) );
  AOI22X1 U276 ( .A(n352), .B(\PipeEM_Result<12> ), .C(n353), .D(
        \PipeMW_Result<12> ), .Y(n190) );
  OAI21X1 U277 ( .A(n495), .B(n378), .C(n191), .Y(N49) );
  AOI22X1 U278 ( .A(n352), .B(\PipeEM_Result<11> ), .C(n353), .D(
        \PipeMW_Result<11> ), .Y(n191) );
  OAI21X1 U279 ( .A(n494), .B(n378), .C(n192), .Y(N48) );
  AOI22X1 U280 ( .A(n352), .B(\PipeEM_Result<10> ), .C(n353), .D(
        \PipeMW_Result<10> ), .Y(n192) );
  OAI21X1 U281 ( .A(n493), .B(n378), .C(n193), .Y(N47) );
  AOI22X1 U282 ( .A(n352), .B(\PipeEM_Result<9> ), .C(n353), .D(
        \PipeMW_Result<9> ), .Y(n193) );
  OAI21X1 U283 ( .A(n492), .B(n377), .C(n194), .Y(N46) );
  AOI22X1 U284 ( .A(n352), .B(\PipeEM_Result<8> ), .C(n353), .D(
        \PipeMW_Result<8> ), .Y(n194) );
  OAI21X1 U285 ( .A(n491), .B(n377), .C(n195), .Y(N45) );
  AOI22X1 U286 ( .A(n352), .B(\PipeEM_Result<7> ), .C(n353), .D(
        \PipeMW_Result<7> ), .Y(n195) );
  OAI21X1 U287 ( .A(n490), .B(n377), .C(n196), .Y(N44) );
  AOI22X1 U288 ( .A(n352), .B(\PipeEM_Result<6> ), .C(n353), .D(
        \PipeMW_Result<6> ), .Y(n196) );
  OAI21X1 U289 ( .A(n489), .B(n377), .C(n197), .Y(N43) );
  AOI22X1 U290 ( .A(n352), .B(\PipeEM_Result<5> ), .C(n353), .D(
        \PipeMW_Result<5> ), .Y(n197) );
  OAI21X1 U291 ( .A(n488), .B(n377), .C(n198), .Y(N42) );
  AOI22X1 U292 ( .A(n352), .B(\PipeEM_Result<4> ), .C(n353), .D(
        \PipeMW_Result<4> ), .Y(n198) );
  OAI21X1 U293 ( .A(n487), .B(n377), .C(n199), .Y(N41) );
  AOI22X1 U294 ( .A(n352), .B(\PipeEM_Result<3> ), .C(n353), .D(
        \PipeMW_Result<3> ), .Y(n199) );
  OAI21X1 U295 ( .A(n486), .B(n377), .C(n200), .Y(N40) );
  AOI22X1 U296 ( .A(n352), .B(\PipeEM_Result<2> ), .C(n353), .D(
        \PipeMW_Result<2> ), .Y(n200) );
  OAI21X1 U297 ( .A(n485), .B(n377), .C(n201), .Y(N39) );
  AOI22X1 U298 ( .A(n352), .B(\PipeEM_Result<1> ), .C(n353), .D(
        \PipeMW_Result<1> ), .Y(n201) );
  OAI21X1 U299 ( .A(n484), .B(n377), .C(n202), .Y(N38) );
  AOI22X1 U300 ( .A(n352), .B(\PipeEM_Result<0> ), .C(n353), .D(
        \PipeMW_Result<0> ), .Y(n202) );
  AOI21X1 U305 ( .A(branch_en), .B(Branch), .C(Jump), .Y(n146) );
  alu primary_alu ( .A({n337, n347, n345, n343, n335, n333, n77, n332, n330, 
        n341, n339, n297, n73, n151, n259, n184}), .B({\alu_operand_b<15> , 
        \alu_operand_b<14> , \alu_operand_b<13> , \alu_operand_b<12> , 
        \alu_operand_b<11> , n137, n132, \alu_operand_b<8> , n65, n127, n123, 
        n119, n61, n57, n53, n50}), .Cin(Cin), .Op({\Opcode<2> , \Opcode<1> , 
        \Opcode<0> }), .invA(InvA), .invB(InvB), .sign(1'b1), .Out({
        \aluResult<15> , \aluResult<14> , \aluResult<13> , \aluResult<12> , 
        \aluResult<11> , \aluResult<10> , \aluResult<9> , \aluResult<8> , 
        \aluResult<7> , \aluResult<6> , \aluResult<5> , \aluResult<4> , 
        \aluResult<3> , \aluResult<2> , \aluResult<1> , \aluResult<0> }), 
        .Ofl(), .Z(Zero), .Cout(cout) );
  mux4to1_16_5 set_mux ( .InA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n38}), .InB({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \_2_net_<0> }), .InC({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n75}), .InD({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, cout}), .S({\Func<1> , \Func<0> }), .Out({\setResult<15> , 
        \setResult<14> , \setResult<13> , \setResult<12> , \setResult<11> , 
        \setResult<10> , \setResult<9> , \setResult<8> , \setResult<7> , 
        \setResult<6> , \setResult<5> , \setResult<4> , \setResult<3> , 
        \setResult<2> , \setResult<1> , \setResult<0> }) );
  cla16_1 addr_adder ( .A({\DecodeIncPC<15> , \DecodeIncPC<14> , 
        \DecodeIncPC<13> , \DecodeIncPC<12> , \DecodeIncPC<11> , n19, 
        \DecodeIncPC<9> , \DecodeIncPC<8> , \DecodeIncPC<7> , \DecodeIncPC<6> , 
        \DecodeIncPC<5> , \DecodeIncPC<4> , \DecodeIncPC<3> , \DecodeIncPC<2> , 
        \DecodeIncPC<1> , \DecodeIncPC<0> }), .B({\Imm<15> , \Imm<14> , 
        \Imm<13> , \Imm<12> , \Imm<11> , \Imm<10> , \Imm<9> , \Imm<8> , 
        \Imm<7> , \Imm<6> , \Imm<5> , \Imm<4> , \Imm<3> , \Imm<2> , \Imm<1> , 
        \Imm<0> }), .Cin(1'b0), .S({\offsetAddr<15> , \offsetAddr<14> , 
        \offsetAddr<13> , \offsetAddr<12> , \offsetAddr<11> , \offsetAddr<10> , 
        \offsetAddr<9> , \offsetAddr<8> , \offsetAddr<7> , \offsetAddr<6> , 
        \offsetAddr<5> , \offsetAddr<4> , \offsetAddr<3> , \offsetAddr<2> , 
        \offsetAddr<1> , \offsetAddr<0> }), .Cout() );
  mux4to1 branchMux ( .InA(n350), .InB(n351), .InC(\ALUOp1<15> ), .InD(n499), 
        .S({\Func<1> , \Func<0> }), .Out(branch_en) );
  INVX1 U3 ( .A(n374), .Y(n1) );
  INVX1 U4 ( .A(n369), .Y(n2) );
  INVX1 U5 ( .A(n369), .Y(n385) );
  OR2X2 U6 ( .A(n43), .B(n430), .Y(n331) );
  INVX1 U7 ( .A(n34), .Y(n3) );
  INVX1 U8 ( .A(n34), .Y(n4) );
  INVX1 U9 ( .A(n34), .Y(n35) );
  INVX2 U10 ( .A(n383), .Y(n5) );
  INVX2 U11 ( .A(n385), .Y(n23) );
  INVX1 U12 ( .A(Link), .Y(n6) );
  INVX1 U13 ( .A(n387), .Y(n34) );
  INVX2 U14 ( .A(n387), .Y(n359) );
  INVX1 U15 ( .A(\OpAReg<12> ), .Y(n434) );
  AND2X1 U16 ( .A(\DecodeIncPC<15> ), .B(n479), .Y(n36) );
  INVX1 U17 ( .A(\Imm<2> ), .Y(n32) );
  INVX1 U18 ( .A(\Imm<0> ), .Y(n28) );
  INVX1 U19 ( .A(\OpAReg<13> ), .Y(n435) );
  INVX1 U21 ( .A(\OpAReg<4> ), .Y(n426) );
  INVX1 U22 ( .A(\OpAReg<0> ), .Y(n422) );
  INVX1 U23 ( .A(\OpAReg<10> ), .Y(n432) );
  INVX1 U24 ( .A(\OpBReg<15> ), .Y(n421) );
  INVX1 U25 ( .A(\DecodeIncPC<0> ), .Y(n458) );
  INVX1 U26 ( .A(\OpBReg<12> ), .Y(n415) );
  INVX1 U27 ( .A(\OpBReg<13> ), .Y(n417) );
  INVX1 U28 ( .A(\OpBReg<14> ), .Y(n419) );
  INVX1 U29 ( .A(\ALUOp1<8> ), .Y(n492) );
  INVX1 U30 ( .A(\ALUOp1<9> ), .Y(n493) );
  INVX1 U31 ( .A(\OpBReg<2> ), .Y(n26) );
  INVX1 U32 ( .A(\OpAReg<9> ), .Y(n431) );
  INVX1 U33 ( .A(\OpAReg<5> ), .Y(n427) );
  INVX1 U34 ( .A(\OpAReg<8> ), .Y(n430) );
  INVX1 U35 ( .A(\OpAReg<6> ), .Y(n428) );
  INVX1 U36 ( .A(\OpAReg<7> ), .Y(n429) );
  INVX1 U37 ( .A(\OpAReg<11> ), .Y(n433) );
  INVX1 U38 ( .A(\OpAReg<14> ), .Y(n436) );
  INVX1 U39 ( .A(n18), .Y(n19) );
  INVX1 U40 ( .A(\OpAReg<15> ), .Y(n437) );
  INVX1 U41 ( .A(\aluResult<1> ), .Y(n483) );
  AND2X1 U42 ( .A(n19), .B(n479), .Y(n246) );
  INVX1 U43 ( .A(n438), .Y(n454) );
  OR2X1 U44 ( .A(n25), .B(n37), .Y(n438) );
  INVX1 U45 ( .A(\aluResult<0> ), .Y(n482) );
  INVX1 U46 ( .A(\ForwardALUOp2<1> ), .Y(n501) );
  INVX1 U47 ( .A(\ForwardALUOp2<0> ), .Y(n500) );
  INVX1 U48 ( .A(\ForwardALUOp1<1> ), .Y(n503) );
  INVX1 U49 ( .A(\ForwardALUOp1<0> ), .Y(n502) );
  INVX1 U50 ( .A(\ALUOp1<6> ), .Y(n490) );
  INVX1 U51 ( .A(\ALUOp1<7> ), .Y(n491) );
  BUFX2 U52 ( .A(n349), .Y(n377) );
  INVX1 U53 ( .A(\ALUOp1<15> ), .Y(n499) );
  INVX1 U54 ( .A(\ALUOp1<0> ), .Y(n484) );
  INVX1 U55 ( .A(\ALUOp1<1> ), .Y(n485) );
  INVX1 U56 ( .A(\ALUOp1<10> ), .Y(n494) );
  OR2X1 U57 ( .A(Btr), .B(n360), .Y(n7) );
  AND2X1 U58 ( .A(n257), .B(n205), .Y(n144) );
  AND2X2 U59 ( .A(n363), .B(\OpBReg<5> ), .Y(n8) );
  AND2X2 U60 ( .A(n368), .B(\OpBReg<0> ), .Y(n9) );
  AND2X2 U61 ( .A(n362), .B(\OpBReg<1> ), .Y(n10) );
  AND2X2 U62 ( .A(n363), .B(\OpBReg<7> ), .Y(n11) );
  AND2X2 U63 ( .A(n363), .B(\OpBReg<4> ), .Y(n12) );
  AND2X2 U64 ( .A(n362), .B(\OpBReg<10> ), .Y(n13) );
  INVX1 U65 ( .A(\OpAReg<2> ), .Y(n371) );
  AND2X1 U66 ( .A(\aluResult<5> ), .B(n25), .Y(n212) );
  AND2X1 U67 ( .A(\aluResult<15> ), .B(n478), .Y(n328) );
  INVX1 U68 ( .A(n365), .Y(n366) );
  INVX1 U69 ( .A(n384), .Y(n14) );
  INVX1 U70 ( .A(n383), .Y(n15) );
  INVX1 U71 ( .A(n385), .Y(n16) );
  AND2X2 U72 ( .A(\aluResult<7> ), .B(n478), .Y(n256) );
  AND2X2 U73 ( .A(\aluResult<13> ), .B(n478), .Y(n324) );
  OR2X2 U74 ( .A(n16), .B(n371), .Y(n424) );
  INVX1 U75 ( .A(n382), .Y(n17) );
  INVX1 U76 ( .A(n382), .Y(n381) );
  INVX2 U77 ( .A(n374), .Y(n33) );
  INVX1 U78 ( .A(\DecodeIncPC<10> ), .Y(n18) );
  INVX1 U79 ( .A(n49), .Y(n20) );
  INVX1 U80 ( .A(n20), .Y(n21) );
  INVX1 U81 ( .A(n17), .Y(n22) );
  INVX1 U82 ( .A(\Imm<3> ), .Y(n30) );
  AND2X2 U83 ( .A(\aluResult<12> ), .B(n25), .Y(n226) );
  BUFX2 U84 ( .A(\aluResult<12> ), .Y(n24) );
  AND2X2 U85 ( .A(n24), .B(n478), .Y(n322) );
  BUFX2 U86 ( .A(n2), .Y(n25) );
  INVX1 U87 ( .A(n6), .Y(n380) );
  OR2X2 U88 ( .A(n1), .B(n26), .Y(n394) );
  NOR3X1 U89 ( .A(n358), .B(n4), .C(n28), .Y(n27) );
  NOR3X1 U90 ( .A(n30), .B(n4), .C(n22), .Y(n29) );
  INVX1 U91 ( .A(n386), .Y(n384) );
  NOR3X1 U92 ( .A(n35), .B(n32), .C(n365), .Y(n31) );
  INVX1 U93 ( .A(JumpReg), .Y(n387) );
  BUFX2 U94 ( .A(n146), .Y(n37) );
  BUFX2 U95 ( .A(Zero), .Y(n38) );
  INVX1 U96 ( .A(Link), .Y(n382) );
  NAND2X1 U97 ( .A(\DecodeIncPC<10> ), .B(n3), .Y(n39) );
  AND2X2 U98 ( .A(n5), .B(n40), .Y(n139) );
  INVX1 U99 ( .A(n39), .Y(n40) );
  OR2X2 U100 ( .A(n381), .B(n371), .Y(n376) );
  INVX1 U101 ( .A(n383), .Y(n367) );
  INVX1 U102 ( .A(n21), .Y(n41) );
  INVX1 U103 ( .A(n49), .Y(n42) );
  INVX1 U104 ( .A(n20), .Y(n43) );
  INVX1 U105 ( .A(n42), .Y(n44) );
  INVX1 U106 ( .A(n41), .Y(n45) );
  INVX1 U107 ( .A(n41), .Y(n46) );
  INVX1 U108 ( .A(n42), .Y(n47) );
  INVX1 U109 ( .A(n42), .Y(n48) );
  OR2X2 U110 ( .A(n48), .B(n435), .Y(n344) );
  OR2X2 U111 ( .A(n46), .B(n436), .Y(n346) );
  OR2X2 U112 ( .A(n48), .B(n426), .Y(n296) );
  AND2X2 U113 ( .A(n372), .B(n386), .Y(n49) );
  OR2X2 U114 ( .A(n9), .B(n51), .Y(n50) );
  OR2X2 U115 ( .A(n52), .B(n27), .Y(n51) );
  INVX1 U116 ( .A(n390), .Y(n52) );
  OR2X2 U117 ( .A(n10), .B(n54), .Y(n53) );
  OR2X2 U118 ( .A(n55), .B(n56), .Y(n54) );
  INVX1 U119 ( .A(n391), .Y(n55) );
  INVX1 U129 ( .A(n392), .Y(n56) );
  OR2X2 U130 ( .A(n58), .B(n60), .Y(n57) );
  OR2X2 U131 ( .A(n31), .B(n59), .Y(n58) );
  INVX1 U132 ( .A(n394), .Y(n59) );
  INVX1 U133 ( .A(n393), .Y(n60) );
  OR2X2 U134 ( .A(n64), .B(n62), .Y(n61) );
  OR2X2 U135 ( .A(n29), .B(n63), .Y(n62) );
  INVX1 U136 ( .A(n396), .Y(n63) );
  INVX1 U137 ( .A(n395), .Y(n64) );
  OR2X2 U138 ( .A(n11), .B(n66), .Y(n65) );
  OR2X2 U139 ( .A(n67), .B(n68), .Y(n66) );
  INVX1 U140 ( .A(n404), .Y(n67) );
  INVX1 U141 ( .A(n405), .Y(n68) );
  OR2X2 U142 ( .A(n36), .B(n70), .Y(\Result<15> ) );
  OR2X2 U143 ( .A(n328), .B(n71), .Y(n70) );
  INVX1 U144 ( .A(n477), .Y(n71) );
  OR2X2 U145 ( .A(n43), .B(n425), .Y(n72) );
  INVX1 U146 ( .A(n72), .Y(n73) );
  AND2X2 U147 ( .A(n388), .B(n389), .Y(n74) );
  INVX1 U148 ( .A(n74), .Y(n75) );
  OR2X2 U149 ( .A(n21), .B(n431), .Y(n76) );
  INVX1 U150 ( .A(n76), .Y(n77) );
  AND2X2 U151 ( .A(n441), .B(n207), .Y(n78) );
  INVX1 U152 ( .A(n78), .Y(\NextPC<2> ) );
  AND2X2 U153 ( .A(n442), .B(n209), .Y(n80) );
  INVX1 U154 ( .A(n80), .Y(\NextPC<3> ) );
  AND2X2 U155 ( .A(n443), .B(n211), .Y(n82) );
  INVX1 U156 ( .A(n82), .Y(\NextPC<4> ) );
  AND2X2 U157 ( .A(n444), .B(n213), .Y(n93) );
  INVX1 U159 ( .A(n93), .Y(\NextPC<5> ) );
  AND2X2 U160 ( .A(n445), .B(n215), .Y(n95) );
  INVX1 U161 ( .A(n95), .Y(\NextPC<6> ) );
  AND2X2 U162 ( .A(n446), .B(n217), .Y(n97) );
  INVX1 U163 ( .A(n97), .Y(\NextPC<7> ) );
  AND2X2 U164 ( .A(n447), .B(n219), .Y(n99) );
  INVX1 U165 ( .A(n99), .Y(\NextPC<8> ) );
  AND2X2 U166 ( .A(n448), .B(n221), .Y(n101) );
  INVX1 U167 ( .A(n101), .Y(\NextPC<9> ) );
  AND2X2 U168 ( .A(n449), .B(n223), .Y(n103) );
  INVX1 U169 ( .A(n103), .Y(\NextPC<10> ) );
  AND2X2 U170 ( .A(n450), .B(n225), .Y(n105) );
  INVX1 U171 ( .A(n105), .Y(\NextPC<11> ) );
  AND2X2 U172 ( .A(n451), .B(n227), .Y(n107) );
  INVX1 U173 ( .A(n107), .Y(\NextPC<12> ) );
  AND2X2 U174 ( .A(n452), .B(n229), .Y(n109) );
  INVX1 U175 ( .A(n109), .Y(\NextPC<13> ) );
  AND2X2 U176 ( .A(n453), .B(n231), .Y(n111) );
  INVX1 U177 ( .A(n111), .Y(\NextPC<14> ) );
  AND2X2 U178 ( .A(n456), .B(n457), .Y(n115) );
  INVX1 U179 ( .A(n115), .Y(\NextPC<15> ) );
  AND2X2 U180 ( .A(n113), .B(n114), .Y(n117) );
  INVX1 U181 ( .A(n117), .Y(\Result<1> ) );
  OR2X2 U182 ( .A(n12), .B(n120), .Y(n119) );
  OR2X2 U183 ( .A(n121), .B(n122), .Y(n120) );
  INVX1 U184 ( .A(n397), .Y(n121) );
  INVX1 U185 ( .A(n398), .Y(n122) );
  OR2X2 U186 ( .A(n126), .B(n124), .Y(n123) );
  OR2X2 U187 ( .A(n125), .B(n8), .Y(n124) );
  INVX1 U188 ( .A(n399), .Y(n125) );
  INVX1 U189 ( .A(n400), .Y(n126) );
  OR2X2 U190 ( .A(n131), .B(n128), .Y(n127) );
  OR2X2 U191 ( .A(n129), .B(n130), .Y(n128) );
  INVX1 U192 ( .A(n401), .Y(n129) );
  INVX1 U193 ( .A(n402), .Y(n130) );
  INVX1 U194 ( .A(n403), .Y(n131) );
  OR2X2 U195 ( .A(n136), .B(n133), .Y(n132) );
  OR2X2 U196 ( .A(n135), .B(n134), .Y(n133) );
  INVX1 U197 ( .A(n408), .Y(n134) );
  INVX1 U198 ( .A(n409), .Y(n135) );
  INVX1 U199 ( .A(n410), .Y(n136) );
  OR2X2 U200 ( .A(n140), .B(n138), .Y(n137) );
  OR2X2 U201 ( .A(n13), .B(n139), .Y(n138) );
  INVX1 U202 ( .A(n411), .Y(n140) );
  OR2X1 U203 ( .A(Set), .B(n7), .Y(n141) );
  AND2X2 U204 ( .A(n469), .B(n144), .Y(n142) );
  INVX1 U205 ( .A(n142), .Y(\Result<7> ) );
  AND2X2 U206 ( .A(n424), .B(n376), .Y(n145) );
  INVX1 U207 ( .A(n145), .Y(n151) );
  OR2X2 U208 ( .A(n14), .B(n22), .Y(n152) );
  OR2X1 U209 ( .A(n44), .B(n422), .Y(n153) );
  INVX1 U210 ( .A(n153), .Y(n184) );
  OR2X2 U211 ( .A(n49), .B(n432), .Y(n186) );
  AND2X2 U212 ( .A(n363), .B(\OpBReg<11> ), .Y(n187) );
  INVX1 U213 ( .A(n187), .Y(n203) );
  AND2X2 U214 ( .A(\DecodeIncPC<7> ), .B(n479), .Y(n204) );
  INVX1 U215 ( .A(n204), .Y(n205) );
  AND2X2 U218 ( .A(\aluResult<2> ), .B(n25), .Y(n206) );
  INVX1 U219 ( .A(n206), .Y(n207) );
  AND2X2 U222 ( .A(\aluResult<3> ), .B(n25), .Y(n208) );
  INVX1 U225 ( .A(n208), .Y(n209) );
  AND2X2 U228 ( .A(\aluResult<4> ), .B(n25), .Y(n210) );
  INVX1 U231 ( .A(n210), .Y(n211) );
  INVX1 U234 ( .A(n212), .Y(n213) );
  AND2X2 U237 ( .A(\aluResult<6> ), .B(n25), .Y(n214) );
  INVX1 U240 ( .A(n214), .Y(n215) );
  AND2X2 U243 ( .A(\aluResult<7> ), .B(n25), .Y(n216) );
  INVX1 U246 ( .A(n216), .Y(n217) );
  AND2X2 U249 ( .A(\aluResult<8> ), .B(n25), .Y(n218) );
  INVX1 U252 ( .A(n218), .Y(n219) );
  AND2X2 U255 ( .A(\aluResult<9> ), .B(n25), .Y(n220) );
  INVX1 U258 ( .A(n220), .Y(n221) );
  AND2X2 U261 ( .A(\aluResult<10> ), .B(n25), .Y(n222) );
  INVX1 U264 ( .A(n222), .Y(n223) );
  AND2X2 U266 ( .A(\aluResult<11> ), .B(n25), .Y(n224) );
  INVX1 U267 ( .A(n224), .Y(n225) );
  INVX1 U270 ( .A(n226), .Y(n227) );
  AND2X2 U301 ( .A(\aluResult<13> ), .B(n25), .Y(n228) );
  INVX1 U302 ( .A(n228), .Y(n229) );
  AND2X2 U303 ( .A(\aluResult<14> ), .B(n25), .Y(n230) );
  INVX1 U304 ( .A(n230), .Y(n231) );
  INVX1 U307 ( .A(n372), .Y(n363) );
  AND2X2 U308 ( .A(\DecodeIncPC<2> ), .B(n479), .Y(n232) );
  INVX1 U309 ( .A(n232), .Y(n233) );
  AND2X2 U310 ( .A(\DecodeIncPC<3> ), .B(n479), .Y(n234) );
  INVX1 U311 ( .A(n234), .Y(n235) );
  AND2X2 U312 ( .A(\DecodeIncPC<4> ), .B(n479), .Y(n236) );
  INVX1 U313 ( .A(n236), .Y(n237) );
  AND2X2 U314 ( .A(\DecodeIncPC<5> ), .B(n479), .Y(n238) );
  INVX1 U315 ( .A(n238), .Y(n239) );
  AND2X2 U316 ( .A(\DecodeIncPC<6> ), .B(n479), .Y(n240) );
  INVX1 U317 ( .A(n240), .Y(n241) );
  AND2X2 U318 ( .A(\DecodeIncPC<8> ), .B(n479), .Y(n242) );
  INVX1 U319 ( .A(n242), .Y(n243) );
  AND2X2 U320 ( .A(\DecodeIncPC<9> ), .B(n479), .Y(n244) );
  INVX1 U321 ( .A(n244), .Y(n245) );
  INVX1 U322 ( .A(n246), .Y(n247) );
  AND2X2 U323 ( .A(\DecodeIncPC<11> ), .B(n479), .Y(n248) );
  INVX1 U324 ( .A(n248), .Y(n249) );
  AND2X2 U325 ( .A(\DecodeIncPC<12> ), .B(n479), .Y(n250) );
  INVX1 U326 ( .A(n250), .Y(n251) );
  AND2X2 U327 ( .A(\DecodeIncPC<13> ), .B(n479), .Y(n252) );
  INVX1 U328 ( .A(n252), .Y(n253) );
  AND2X2 U329 ( .A(\DecodeIncPC<14> ), .B(n479), .Y(n254) );
  INVX1 U330 ( .A(n254), .Y(n255) );
  INVX1 U331 ( .A(Btr), .Y(n460) );
  INVX1 U332 ( .A(n256), .Y(n257) );
  AND2X2 U333 ( .A(n373), .B(n423), .Y(n258) );
  INVX1 U334 ( .A(n258), .Y(n259) );
  AND2X2 U335 ( .A(n182), .B(n183), .Y(n260) );
  INVX1 U336 ( .A(n260), .Y(n261) );
  AND2X2 U337 ( .A(n180), .B(n181), .Y(n262) );
  INVX1 U338 ( .A(n262), .Y(n263) );
  AND2X2 U339 ( .A(n178), .B(n179), .Y(n264) );
  INVX1 U340 ( .A(n264), .Y(n265) );
  AND2X2 U341 ( .A(n176), .B(n177), .Y(n266) );
  INVX1 U342 ( .A(n266), .Y(n267) );
  AND2X2 U343 ( .A(n174), .B(n175), .Y(n268) );
  INVX1 U344 ( .A(n268), .Y(n269) );
  AND2X2 U345 ( .A(n172), .B(n173), .Y(n270) );
  INVX1 U346 ( .A(n270), .Y(n271) );
  AND2X2 U347 ( .A(n170), .B(n171), .Y(n272) );
  INVX1 U348 ( .A(n272), .Y(n273) );
  AND2X2 U349 ( .A(n168), .B(n169), .Y(n274) );
  INVX1 U350 ( .A(n274), .Y(n275) );
  AND2X2 U351 ( .A(n166), .B(n167), .Y(n276) );
  INVX1 U352 ( .A(n276), .Y(n277) );
  AND2X2 U353 ( .A(n164), .B(n165), .Y(n278) );
  INVX1 U354 ( .A(n278), .Y(n279) );
  AND2X2 U355 ( .A(n162), .B(n163), .Y(n280) );
  INVX1 U356 ( .A(n280), .Y(n281) );
  AND2X2 U357 ( .A(n160), .B(n161), .Y(n282) );
  INVX1 U358 ( .A(n282), .Y(n283) );
  AND2X2 U359 ( .A(n158), .B(n159), .Y(n284) );
  INVX1 U360 ( .A(n284), .Y(n285) );
  AND2X2 U361 ( .A(n156), .B(n157), .Y(n286) );
  INVX1 U362 ( .A(n286), .Y(n287) );
  AND2X2 U363 ( .A(n154), .B(n155), .Y(n288) );
  INVX1 U364 ( .A(n288), .Y(n289) );
  AND2X2 U365 ( .A(n147), .B(n148), .Y(n290) );
  INVX1 U366 ( .A(n290), .Y(n291) );
  OR2X1 U367 ( .A(n353), .B(n293), .Y(n292) );
  OR2X1 U368 ( .A(n352), .B(n348), .Y(n293) );
  OR2X1 U369 ( .A(n355), .B(n295), .Y(n294) );
  OR2X1 U370 ( .A(n354), .B(n356), .Y(n295) );
  INVX1 U371 ( .A(n296), .Y(n297) );
  AND2X1 U372 ( .A(\aluResult<0> ), .B(n478), .Y(n298) );
  INVX1 U373 ( .A(n298), .Y(n299) );
  BUFX2 U374 ( .A(n149), .Y(n379) );
  AND2X1 U375 ( .A(ALUSrc), .B(n356), .Y(n150) );
  BUFX2 U376 ( .A(n507), .Y(\Result<2> ) );
  BUFX2 U377 ( .A(n506), .Y(\Result<4> ) );
  BUFX2 U378 ( .A(n505), .Y(\Result<5> ) );
  BUFX2 U379 ( .A(n504), .Y(\Result<9> ) );
  AND2X1 U380 ( .A(\aluResult<2> ), .B(n478), .Y(n304) );
  INVX1 U381 ( .A(n304), .Y(n305) );
  AND2X1 U382 ( .A(\aluResult<3> ), .B(n478), .Y(n306) );
  INVX1 U383 ( .A(n306), .Y(n307) );
  AND2X1 U384 ( .A(\aluResult<4> ), .B(n478), .Y(n308) );
  INVX1 U385 ( .A(n308), .Y(n309) );
  AND2X1 U386 ( .A(\aluResult<5> ), .B(n478), .Y(n310) );
  INVX1 U387 ( .A(n310), .Y(n311) );
  AND2X1 U388 ( .A(\aluResult<6> ), .B(n478), .Y(n312) );
  INVX1 U389 ( .A(n312), .Y(n313) );
  AND2X1 U390 ( .A(\aluResult<8> ), .B(n478), .Y(n314) );
  INVX1 U391 ( .A(n314), .Y(n315) );
  AND2X1 U392 ( .A(\aluResult<9> ), .B(n478), .Y(n316) );
  INVX1 U393 ( .A(n316), .Y(n317) );
  AND2X1 U394 ( .A(\aluResult<10> ), .B(n478), .Y(n318) );
  INVX1 U395 ( .A(n318), .Y(n319) );
  AND2X1 U396 ( .A(\aluResult<11> ), .B(n478), .Y(n320) );
  INVX1 U397 ( .A(n320), .Y(n321) );
  INVX1 U398 ( .A(n322), .Y(n323) );
  INVX1 U399 ( .A(n324), .Y(n325) );
  AND2X1 U400 ( .A(\aluResult<14> ), .B(n478), .Y(n326) );
  INVX1 U401 ( .A(n326), .Y(n327) );
  INVX1 U402 ( .A(\ALUOp1<12> ), .Y(n496) );
  INVX1 U403 ( .A(\ALUOp1<11> ), .Y(n495) );
  INVX1 U404 ( .A(\ALUOp1<14> ), .Y(n498) );
  INVX1 U405 ( .A(\ALUOp1<13> ), .Y(n497) );
  INVX1 U406 ( .A(\ALUOp1<5> ), .Y(n489) );
  INVX1 U407 ( .A(\ALUOp1<4> ), .Y(n488) );
  INVX1 U408 ( .A(\ALUOp1<3> ), .Y(n487) );
  INVX1 U409 ( .A(\ALUOp1<2> ), .Y(n486) );
  OR2X2 U410 ( .A(n43), .B(n429), .Y(n329) );
  INVX1 U411 ( .A(n329), .Y(n330) );
  INVX1 U412 ( .A(n331), .Y(n332) );
  INVX1 U413 ( .A(n186), .Y(n333) );
  OR2X2 U414 ( .A(n47), .B(n433), .Y(n334) );
  INVX1 U415 ( .A(n334), .Y(n335) );
  OR2X2 U416 ( .A(n48), .B(n437), .Y(n336) );
  INVX1 U417 ( .A(n336), .Y(n337) );
  OR2X1 U418 ( .A(n45), .B(n427), .Y(n338) );
  INVX1 U419 ( .A(n338), .Y(n339) );
  OR2X2 U420 ( .A(n48), .B(n428), .Y(n340) );
  INVX1 U421 ( .A(n340), .Y(n341) );
  OR2X2 U422 ( .A(n46), .B(n434), .Y(n342) );
  INVX1 U423 ( .A(n342), .Y(n343) );
  INVX1 U424 ( .A(n344), .Y(n345) );
  INVX1 U425 ( .A(n346), .Y(n347) );
  AND2X1 U426 ( .A(n502), .B(n503), .Y(n348) );
  INVX1 U427 ( .A(n348), .Y(n349) );
  INVX1 U428 ( .A(n351), .Y(n350) );
  BUFX2 U429 ( .A(_7_net_), .Y(n351) );
  AND2X1 U430 ( .A(\ForwardALUOp1<1> ), .B(n502), .Y(n352) );
  AND2X1 U431 ( .A(\ForwardALUOp1<0> ), .B(n503), .Y(n353) );
  AND2X1 U432 ( .A(\ForwardALUOp2<1> ), .B(n500), .Y(n354) );
  AND2X1 U433 ( .A(\ForwardALUOp2<0> ), .B(n501), .Y(n355) );
  INVX1 U434 ( .A(n141), .Y(n479) );
  INVX1 U435 ( .A(n463), .Y(n480) );
  AND2X1 U436 ( .A(n500), .B(n501), .Y(n356) );
  INVX1 U437 ( .A(n356), .Y(n357) );
  INVX1 U438 ( .A(BranchJumpTaken), .Y(n455) );
  BUFX2 U439 ( .A(n349), .Y(n378) );
  INVX1 U440 ( .A(\OpAReg<3> ), .Y(n425) );
  OAI21X1 U441 ( .A(n461), .B(n463), .C(n462), .Y(\Result<0> ) );
  INVX1 U442 ( .A(n372), .Y(n358) );
  BUFX2 U443 ( .A(n23), .Y(n360) );
  INVX1 U444 ( .A(n368), .Y(n361) );
  INVX1 U445 ( .A(n17), .Y(n362) );
  INVX1 U446 ( .A(n17), .Y(n368) );
  NAND2X1 U447 ( .A(\DecodeIncPC<11> ), .B(n47), .Y(n364) );
  AND2X2 U448 ( .A(n364), .B(n203), .Y(n412) );
  INVX1 U449 ( .A(n33), .Y(n365) );
  INVX1 U450 ( .A(Link), .Y(n383) );
  INVX1 U451 ( .A(JumpReg), .Y(n369) );
  INVX1 U452 ( .A(JumpReg), .Y(n386) );
  INVX2 U453 ( .A(n152), .Y(n370) );
  INVX1 U454 ( .A(n6), .Y(n372) );
  NAND2X1 U455 ( .A(n363), .B(\OpAReg<1> ), .Y(n373) );
  INVX1 U456 ( .A(Link), .Y(n374) );
  MUX2X1 U457 ( .B(\ALUOp1<15> ), .A(\aluResult<15> ), .S(n375), .Y(n388) );
  XNOR2X1 U458 ( .A(\ALUOp1<15> ), .B(\ALUOp2<15> ), .Y(n375) );
  INVX1 U459 ( .A(n388), .Y(\_2_net_<0> ) );
  INVX1 U460 ( .A(Zero), .Y(n389) );
  INVX1 U461 ( .A(\setResult<0> ), .Y(n461) );
  NAND3X1 U462 ( .A(n3), .B(\DecodeIncPC<0> ), .C(n380), .Y(n390) );
  NAND3X1 U463 ( .A(n3), .B(\DecodeIncPC<1> ), .C(n367), .Y(n392) );
  NAND3X1 U464 ( .A(n359), .B(\Imm<1> ), .C(n33), .Y(n391) );
  NAND3X1 U465 ( .A(n23), .B(\DecodeIncPC<2> ), .C(n381), .Y(n393) );
  NAND2X1 U466 ( .A(n368), .B(\OpBReg<3> ), .Y(n396) );
  NAND3X1 U467 ( .A(n23), .B(\DecodeIncPC<3> ), .C(n15), .Y(n395) );
  NAND3X1 U468 ( .A(n2), .B(\Imm<4> ), .C(n361), .Y(n398) );
  NAND3X1 U469 ( .A(n5), .B(n14), .C(\DecodeIncPC<4> ), .Y(n397) );
  NAND3X1 U470 ( .A(n2), .B(\Imm<5> ), .C(n5), .Y(n400) );
  NAND3X1 U471 ( .A(n14), .B(\DecodeIncPC<5> ), .C(n5), .Y(n399) );
  NAND3X1 U472 ( .A(n23), .B(\DecodeIncPC<6> ), .C(n381), .Y(n403) );
  NAND2X1 U473 ( .A(n362), .B(\OpBReg<6> ), .Y(n402) );
  NAND3X1 U474 ( .A(n359), .B(\Imm<6> ), .C(n381), .Y(n401) );
  NAND3X1 U475 ( .A(n2), .B(\Imm<7> ), .C(n15), .Y(n405) );
  NAND3X1 U476 ( .A(n14), .B(\DecodeIncPC<7> ), .C(n361), .Y(n404) );
  INVX2 U477 ( .A(\Imm<8> ), .Y(n407) );
  AOI22X1 U478 ( .A(\DecodeIncPC<8> ), .B(n44), .C(n362), .D(\OpBReg<8> ), .Y(
        n406) );
  OAI21X1 U479 ( .A(n152), .B(n407), .C(n406), .Y(\alu_operand_b<8> ) );
  NAND3X1 U480 ( .A(n14), .B(\DecodeIncPC<9> ), .C(n5), .Y(n410) );
  NAND3X1 U481 ( .A(n384), .B(\Imm<9> ), .C(n380), .Y(n409) );
  NAND2X1 U482 ( .A(\OpBReg<9> ), .B(n358), .Y(n408) );
  NAND3X1 U483 ( .A(n2), .B(\Imm<10> ), .C(n15), .Y(n411) );
  INVX2 U484 ( .A(\Imm<11> ), .Y(n413) );
  OAI21X1 U485 ( .A(n152), .B(n413), .C(n412), .Y(\alu_operand_b<11> ) );
  AOI22X1 U486 ( .A(\DecodeIncPC<12> ), .B(n46), .C(\Imm<12> ), .D(n370), .Y(
        n414) );
  OAI21X1 U487 ( .A(n415), .B(n366), .C(n414), .Y(\alu_operand_b<12> ) );
  AOI22X1 U488 ( .A(\DecodeIncPC<13> ), .B(n47), .C(\Imm<13> ), .D(n370), .Y(
        n416) );
  OAI21X1 U489 ( .A(n417), .B(n366), .C(n416), .Y(\alu_operand_b<13> ) );
  AOI22X1 U490 ( .A(\DecodeIncPC<14> ), .B(n45), .C(\Imm<14> ), .D(n370), .Y(
        n418) );
  OAI21X1 U491 ( .A(n419), .B(n366), .C(n418), .Y(\alu_operand_b<14> ) );
  AOI22X1 U492 ( .A(\DecodeIncPC<15> ), .B(n46), .C(\Imm<15> ), .D(n370), .Y(
        n420) );
  OAI21X1 U493 ( .A(n421), .B(n366), .C(n420), .Y(\alu_operand_b<15> ) );
  NAND2X1 U494 ( .A(\OpAReg<1> ), .B(n359), .Y(n423) );
  NAND2X1 U495 ( .A(n360), .B(n146), .Y(BranchJumpTaken) );
  AOI22X1 U496 ( .A(\IncPC<0> ), .B(n455), .C(\offsetAddr<0> ), .D(n454), .Y(
        n439) );
  OAI21X1 U497 ( .A(n360), .B(n482), .C(n439), .Y(\NextPC<0> ) );
  AOI22X1 U498 ( .A(\IncPC<1> ), .B(n455), .C(\offsetAddr<1> ), .D(n454), .Y(
        n440) );
  OAI21X1 U499 ( .A(n360), .B(n483), .C(n440), .Y(\NextPC<1> ) );
  AOI22X1 U500 ( .A(\IncPC<2> ), .B(n455), .C(\offsetAddr<2> ), .D(n454), .Y(
        n441) );
  AOI22X1 U501 ( .A(\IncPC<3> ), .B(n455), .C(\offsetAddr<3> ), .D(n454), .Y(
        n442) );
  AOI22X1 U502 ( .A(\IncPC<4> ), .B(n455), .C(\offsetAddr<4> ), .D(n454), .Y(
        n443) );
  AOI22X1 U503 ( .A(\IncPC<5> ), .B(n455), .C(\offsetAddr<5> ), .D(n454), .Y(
        n444) );
  AOI22X1 U504 ( .A(\IncPC<6> ), .B(n455), .C(\offsetAddr<6> ), .D(n454), .Y(
        n445) );
  AOI22X1 U505 ( .A(\IncPC<7> ), .B(n455), .C(\offsetAddr<7> ), .D(n454), .Y(
        n446) );
  AOI22X1 U506 ( .A(\IncPC<8> ), .B(n455), .C(\offsetAddr<8> ), .D(n454), .Y(
        n447) );
  AOI22X1 U507 ( .A(\IncPC<9> ), .B(n455), .C(\offsetAddr<9> ), .D(n454), .Y(
        n448) );
  AOI22X1 U508 ( .A(\IncPC<10> ), .B(n455), .C(\offsetAddr<10> ), .D(n454), 
        .Y(n449) );
  AOI22X1 U509 ( .A(\IncPC<11> ), .B(n455), .C(\offsetAddr<11> ), .D(n454), 
        .Y(n450) );
  AOI22X1 U510 ( .A(\IncPC<12> ), .B(n455), .C(\offsetAddr<12> ), .D(n454), 
        .Y(n451) );
  AOI22X1 U511 ( .A(\IncPC<13> ), .B(n455), .C(\offsetAddr<13> ), .D(n454), 
        .Y(n452) );
  AOI22X1 U512 ( .A(\IncPC<14> ), .B(n455), .C(\offsetAddr<14> ), .D(n454), 
        .Y(n453) );
  NAND2X1 U513 ( .A(n25), .B(\aluResult<15> ), .Y(n457) );
  AOI22X1 U514 ( .A(\IncPC<15> ), .B(n455), .C(\offsetAddr<15> ), .D(n454), 
        .Y(n456) );
  NOR3X1 U515 ( .A(Btr), .B(n25), .C(Set), .Y(n478) );
  OAI21X1 U516 ( .A(n141), .B(n458), .C(n299), .Y(n459) );
  AOI21X1 U517 ( .A(\ALUOp1<15> ), .B(Btr), .C(n459), .Y(n462) );
  NAND2X1 U518 ( .A(n460), .B(Set), .Y(n463) );
  AOI22X1 U519 ( .A(\ALUOp1<13> ), .B(Btr), .C(\setResult<2> ), .D(n480), .Y(
        n464) );
  NAND3X1 U520 ( .A(n233), .B(n464), .C(n305), .Y(n507) );
  AOI22X1 U521 ( .A(\ALUOp1<12> ), .B(Btr), .C(\setResult<3> ), .D(n480), .Y(
        n465) );
  NAND3X1 U522 ( .A(n235), .B(n465), .C(n307), .Y(\Result<3> ) );
  AOI22X1 U523 ( .A(\ALUOp1<11> ), .B(Btr), .C(\setResult<4> ), .D(n480), .Y(
        n466) );
  NAND3X1 U524 ( .A(n237), .B(n466), .C(n309), .Y(n506) );
  AOI22X1 U525 ( .A(\ALUOp1<10> ), .B(Btr), .C(\setResult<5> ), .D(n480), .Y(
        n467) );
  NAND3X1 U526 ( .A(n239), .B(n467), .C(n311), .Y(n505) );
  AOI22X1 U527 ( .A(\ALUOp1<9> ), .B(Btr), .C(\setResult<6> ), .D(n480), .Y(
        n468) );
  NAND3X1 U528 ( .A(n241), .B(n468), .C(n313), .Y(\Result<6> ) );
  AOI22X1 U529 ( .A(\ALUOp1<8> ), .B(Btr), .C(\setResult<7> ), .D(n480), .Y(
        n469) );
  AOI22X1 U530 ( .A(\ALUOp1<7> ), .B(Btr), .C(\setResult<8> ), .D(n480), .Y(
        n470) );
  NAND3X1 U531 ( .A(n243), .B(n470), .C(n315), .Y(\Result<8> ) );
  AOI22X1 U532 ( .A(\ALUOp1<6> ), .B(Btr), .C(\setResult<9> ), .D(n480), .Y(
        n471) );
  NAND3X1 U533 ( .A(n245), .B(n471), .C(n317), .Y(n504) );
  AOI22X1 U534 ( .A(\ALUOp1<5> ), .B(Btr), .C(\setResult<10> ), .D(n480), .Y(
        n472) );
  NAND3X1 U535 ( .A(n247), .B(n472), .C(n319), .Y(\Result<10> ) );
  AOI22X1 U536 ( .A(\ALUOp1<4> ), .B(Btr), .C(\setResult<11> ), .D(n480), .Y(
        n473) );
  NAND3X1 U537 ( .A(n249), .B(n473), .C(n321), .Y(\Result<11> ) );
  AOI22X1 U538 ( .A(\ALUOp1<3> ), .B(Btr), .C(\setResult<12> ), .D(n480), .Y(
        n474) );
  NAND3X1 U539 ( .A(n251), .B(n474), .C(n323), .Y(\Result<12> ) );
  AOI22X1 U540 ( .A(\ALUOp1<2> ), .B(Btr), .C(\setResult<13> ), .D(n480), .Y(
        n475) );
  NAND3X1 U541 ( .A(n253), .B(n475), .C(n325), .Y(\Result<13> ) );
  AOI22X1 U542 ( .A(\ALUOp1<1> ), .B(Btr), .C(\setResult<14> ), .D(n480), .Y(
        n476) );
  NAND3X1 U543 ( .A(n255), .B(n476), .C(n327), .Y(\Result<14> ) );
  AOI22X1 U544 ( .A(\ALUOp1<0> ), .B(Btr), .C(\setResult<15> ), .D(n480), .Y(
        n477) );
  AOI22X1 U545 ( .A(\DecodeIncPC<1> ), .B(n479), .C(\aluResult<1> ), .D(n478), 
        .Y(n114) );
endmodule


module pipe_em ( Stall, rst, clk, .Result({\Result<15> , \Result<14> , 
        \Result<13> , \Result<12> , \Result<11> , \Result<10> , \Result<9> , 
        \Result<8> , \Result<7> , \Result<6> , \Result<5> , \Result<4> , 
        \Result<3> , \Result<2> , \Result<1> , \Result<0> }), MemRead, 
        MemWrite, MemToReg, Halt, .ALUOp2({\ALUOp2<15> , \ALUOp2<14> , 
        \ALUOp2<13> , \ALUOp2<12> , \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , 
        \ALUOp2<8> , \ALUOp2<7> , \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , 
        \ALUOp2<3> , \ALUOp2<2> , \ALUOp2<1> , \ALUOp2<0> }), RegFileWrEn, 
    .Rs({\Rs<2> , \Rs<1> , \Rs<0> }), .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({
        \Rd<2> , \Rd<1> , \Rd<0> }), .WriteReg({\WriteReg<2> , \WriteReg<1> , 
        \WriteReg<0> }), .Address({\Address<15> , \Address<14> , \Address<13> , 
        \Address<12> , \Address<11> , \Address<10> , \Address<9> , 
        \Address<8> , \Address<7> , \Address<6> , \Address<5> , \Address<4> , 
        \Address<3> , \Address<2> , \Address<1> , \Address<0> }), MemRead_Out, 
        MemWrite_Out, MemToReg_Out, Halt_Out, .WriteData({\WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), RegFileWrEn_Out, 
    .Rs_Out({\Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> }), .Rt_Out({\Rt_Out<2> , 
        \Rt_Out<1> , \Rt_Out<0> }), .Rd_Out({\Rd_Out<2> , \Rd_Out<1> , 
        \Rd_Out<0> }), .WriteReg_Out({\WriteReg_Out<2> , \WriteReg_Out<1> , 
        \WriteReg_Out<0> }) );
  input Stall, rst, clk, \Result<15> , \Result<14> , \Result<13> ,
         \Result<12> , \Result<11> , \Result<10> , \Result<9> , \Result<8> ,
         \Result<7> , \Result<6> , \Result<5> , \Result<4> , \Result<3> ,
         \Result<2> , \Result<1> , \Result<0> , MemRead, MemWrite, MemToReg,
         Halt, \ALUOp2<15> , \ALUOp2<14> , \ALUOp2<13> , \ALUOp2<12> ,
         \ALUOp2<11> , \ALUOp2<10> , \ALUOp2<9> , \ALUOp2<8> , \ALUOp2<7> ,
         \ALUOp2<6> , \ALUOp2<5> , \ALUOp2<4> , \ALUOp2<3> , \ALUOp2<2> ,
         \ALUOp2<1> , \ALUOp2<0> , RegFileWrEn, \Rs<2> , \Rs<1> , \Rs<0> ,
         \Rt<2> , \Rt<1> , \Rt<0> , \Rd<2> , \Rd<1> , \Rd<0> , \WriteReg<2> ,
         \WriteReg<1> , \WriteReg<0> ;
  output \Address<15> , \Address<14> , \Address<13> , \Address<12> ,
         \Address<11> , \Address<10> , \Address<9> , \Address<8> ,
         \Address<7> , \Address<6> , \Address<5> , \Address<4> , \Address<3> ,
         \Address<2> , \Address<1> , \Address<0> , MemRead_Out, MemWrite_Out,
         MemToReg_Out, Halt_Out, \WriteData<15> , \WriteData<14> ,
         \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> ,
         \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> ,
         \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> ,
         \WriteData<1> , \WriteData<0> , RegFileWrEn_Out, \Rs_Out<2> ,
         \Rs_Out<1> , \Rs_Out<0> , \Rt_Out<2> , \Rt_Out<1> , \Rt_Out<0> ,
         \Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> , \WriteReg_Out<2> ,
         \WriteReg_Out<1> , \WriteReg_Out<0> ;
  wire   n121, n122, n123, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n77, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n2, n4, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n69, n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82,
         n83, n84, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120;

  AOI22X1 U51 ( .A(\WriteReg<2> ), .B(n37), .C(\WriteReg_Out<2> ), .D(Stall), 
        .Y(n52) );
  AOI22X1 U52 ( .A(\WriteReg<1> ), .B(n37), .C(\WriteReg_Out<1> ), .D(Stall), 
        .Y(n53) );
  AOI22X1 U53 ( .A(\WriteReg<0> ), .B(n37), .C(\WriteReg_Out<0> ), .D(Stall), 
        .Y(n54) );
  AOI22X1 U54 ( .A(\Rt<2> ), .B(n37), .C(\Rt_Out<2> ), .D(Stall), .Y(n55) );
  AOI22X1 U55 ( .A(\Rt<1> ), .B(n37), .C(\Rt_Out<1> ), .D(Stall), .Y(n56) );
  AOI22X1 U56 ( .A(\Rt<0> ), .B(n37), .C(\Rt_Out<0> ), .D(Stall), .Y(n57) );
  AOI22X1 U57 ( .A(\Rs<2> ), .B(n37), .C(\Rs_Out<2> ), .D(Stall), .Y(n58) );
  AOI22X1 U58 ( .A(\Rs<1> ), .B(n37), .C(\Rs_Out<1> ), .D(Stall), .Y(n59) );
  AOI22X1 U59 ( .A(\Rs<0> ), .B(n37), .C(\Rs_Out<0> ), .D(Stall), .Y(n60) );
  AOI22X1 U60 ( .A(RegFileWrEn), .B(n37), .C(RegFileWrEn_Out), .D(Stall), .Y(
        n61) );
  AOI22X1 U61 ( .A(\Rd<2> ), .B(n37), .C(\Rd_Out<2> ), .D(Stall), .Y(n62) );
  AOI22X1 U62 ( .A(\Rd<1> ), .B(n37), .C(\Rd_Out<1> ), .D(Stall), .Y(n63) );
  AOI22X1 U63 ( .A(\Rd<0> ), .B(n37), .C(\Rd_Out<0> ), .D(Stall), .Y(n64) );
  AOI22X1 U64 ( .A(MemWrite), .B(n37), .C(MemWrite_Out), .D(Stall), .Y(n65) );
  AOI22X1 U65 ( .A(MemToReg), .B(n37), .C(MemToReg_Out), .D(Stall), .Y(n66) );
  AOI22X1 U66 ( .A(MemRead), .B(n37), .C(MemRead_Out), .D(Stall), .Y(n67) );
  AOI22X1 U67 ( .A(Halt), .B(n37), .C(Halt_Out), .D(Stall), .Y(n68) );
  AOI22X1 U76 ( .A(\Address<1> ), .B(Stall), .C(\Result<1> ), .D(n37), .Y(n77)
         );
  AOI22X1 U84 ( .A(\ALUOp2<9> ), .B(n37), .C(\WriteData<9> ), .D(Stall), .Y(
        n85) );
  AOI22X1 U85 ( .A(\ALUOp2<8> ), .B(n37), .C(\WriteData<8> ), .D(Stall), .Y(
        n86) );
  AOI22X1 U86 ( .A(\ALUOp2<7> ), .B(n37), .C(\WriteData<7> ), .D(Stall), .Y(
        n87) );
  AOI22X1 U87 ( .A(\ALUOp2<6> ), .B(n37), .C(\WriteData<6> ), .D(Stall), .Y(
        n88) );
  AOI22X1 U88 ( .A(\ALUOp2<5> ), .B(n37), .C(\WriteData<5> ), .D(Stall), .Y(
        n89) );
  AOI22X1 U89 ( .A(\ALUOp2<4> ), .B(n37), .C(\WriteData<4> ), .D(Stall), .Y(
        n90) );
  AOI22X1 U90 ( .A(\ALUOp2<3> ), .B(n37), .C(\WriteData<3> ), .D(Stall), .Y(
        n91) );
  AOI22X1 U91 ( .A(\ALUOp2<2> ), .B(n37), .C(\WriteData<2> ), .D(Stall), .Y(
        n92) );
  AOI22X1 U92 ( .A(\ALUOp2<1> ), .B(n37), .C(\WriteData<1> ), .D(Stall), .Y(
        n93) );
  AOI22X1 U93 ( .A(\ALUOp2<15> ), .B(n37), .C(\WriteData<15> ), .D(Stall), .Y(
        n94) );
  AOI22X1 U94 ( .A(\ALUOp2<14> ), .B(n37), .C(\WriteData<14> ), .D(Stall), .Y(
        n95) );
  AOI22X1 U95 ( .A(\ALUOp2<13> ), .B(n37), .C(\WriteData<13> ), .D(Stall), .Y(
        n96) );
  AOI22X1 U96 ( .A(\ALUOp2<12> ), .B(n37), .C(\WriteData<12> ), .D(Stall), .Y(
        n97) );
  AOI22X1 U97 ( .A(\ALUOp2<11> ), .B(n37), .C(\WriteData<11> ), .D(Stall), .Y(
        n98) );
  AOI22X1 U98 ( .A(\ALUOp2<10> ), .B(n37), .C(\WriteData<10> ), .D(Stall), .Y(
        n99) );
  AOI22X1 U99 ( .A(\ALUOp2<0> ), .B(n37), .C(\WriteData<0> ), .D(Stall), .Y(
        n100) );
  dff_215 \WriteReg_reg[0]  ( .q(\WriteReg_Out<0> ), .d(n71), .clk(clk), .rst(
        n8) );
  dff_216 \WriteReg_reg[1]  ( .q(\WriteReg_Out<1> ), .d(n72), .clk(clk), .rst(
        n8) );
  dff_217 \WriteReg_reg[2]  ( .q(\WriteReg_Out<2> ), .d(n73), .clk(clk), .rst(
        n8) );
  dff_212 \rs_reg[0]  ( .q(\Rs_Out<0> ), .d(n75), .clk(clk), .rst(n8) );
  dff_213 \rs_reg[1]  ( .q(\Rs_Out<1> ), .d(n76), .clk(clk), .rst(n8) );
  dff_214 \rs_reg[2]  ( .q(\Rs_Out<2> ), .d(n78), .clk(clk), .rst(n8) );
  dff_209 \rt_reg[0]  ( .q(\Rt_Out<0> ), .d(n79), .clk(clk), .rst(n8) );
  dff_210 \rt_reg[1]  ( .q(\Rt_Out<1> ), .d(n80), .clk(clk), .rst(n8) );
  dff_211 \rt_reg[2]  ( .q(\Rt_Out<2> ), .d(n81), .clk(clk), .rst(n8) );
  dff_206 \rd_reg[0]  ( .q(\Rd_Out<0> ), .d(n82), .clk(clk), .rst(n8) );
  dff_207 \rd_reg[1]  ( .q(\Rd_Out<1> ), .d(n83), .clk(clk), .rst(n8) );
  dff_208 \rd_reg[2]  ( .q(\Rd_Out<2> ), .d(n84), .clk(clk), .rst(n8) );
  dff_222 rf_wr_en_reg ( .q(RegFileWrEn_Out), .d(n74), .clk(clk), .rst(n8) );
  dff_190 \address_reg[0]  ( .q(\Address<0> ), .d(n38), .clk(clk), .rst(n7) );
  dff_191 \address_reg[1]  ( .q(\Address<1> ), .d(n70), .clk(clk), .rst(n8) );
  dff_192 \address_reg[2]  ( .q(n123), .d(n39), .clk(clk), .rst(n7) );
  dff_193 \address_reg[3]  ( .q(n122), .d(n40), .clk(clk), .rst(n7) );
  dff_194 \address_reg[4]  ( .q(n121), .d(n41), .clk(clk), .rst(n7) );
  dff_195 \address_reg[5]  ( .q(\Address<5> ), .d(n42), .clk(clk), .rst(n7) );
  dff_196 \address_reg[6]  ( .q(\Address<6> ), .d(n43), .clk(clk), .rst(n7) );
  dff_197 \address_reg[7]  ( .q(\Address<7> ), .d(n44), .clk(clk), .rst(n7) );
  dff_198 \address_reg[8]  ( .q(\Address<8> ), .d(n45), .clk(clk), .rst(n8) );
  dff_199 \address_reg[9]  ( .q(\Address<9> ), .d(n46), .clk(clk), .rst(n7) );
  dff_200 \address_reg[10]  ( .q(\Address<10> ), .d(n47), .clk(clk), .rst(n8)
         );
  dff_201 \address_reg[11]  ( .q(\Address<11> ), .d(n48), .clk(clk), .rst(n7)
         );
  dff_202 \address_reg[12]  ( .q(\Address<12> ), .d(n49), .clk(clk), .rst(n7)
         );
  dff_203 \address_reg[13]  ( .q(\Address<13> ), .d(n50), .clk(clk), .rst(n7)
         );
  dff_204 \address_reg[14]  ( .q(\Address<14> ), .d(n51), .clk(clk), .rst(n8)
         );
  dff_205 \address_reg[15]  ( .q(\Address<15> ), .d(n69), .clk(clk), .rst(n7)
         );
  dff_221 memread_reg ( .q(MemRead_Out), .d(n118), .clk(clk), .rst(n8) );
  dff_220 memwrite_reg ( .q(MemWrite_Out), .d(n117), .clk(clk), .rst(n8) );
  dff_219 memtoreg_reg ( .q(MemToReg_Out), .d(n119), .clk(clk), .rst(n8) );
  dff_174 \writedata_reg[0]  ( .q(\WriteData<0> ), .d(n101), .clk(clk), .rst(
        n8) );
  dff_175 \writedata_reg[1]  ( .q(\WriteData<1> ), .d(n102), .clk(clk), .rst(
        n8) );
  dff_176 \writedata_reg[2]  ( .q(\WriteData<2> ), .d(n103), .clk(clk), .rst(
        n8) );
  dff_177 \writedata_reg[3]  ( .q(\WriteData<3> ), .d(n104), .clk(clk), .rst(
        n8) );
  dff_178 \writedata_reg[4]  ( .q(\WriteData<4> ), .d(n105), .clk(clk), .rst(
        n8) );
  dff_179 \writedata_reg[5]  ( .q(\WriteData<5> ), .d(n106), .clk(clk), .rst(
        n8) );
  dff_180 \writedata_reg[6]  ( .q(\WriteData<6> ), .d(n107), .clk(clk), .rst(
        n8) );
  dff_181 \writedata_reg[7]  ( .q(\WriteData<7> ), .d(n108), .clk(clk), .rst(
        n8) );
  dff_182 \writedata_reg[8]  ( .q(\WriteData<8> ), .d(n109), .clk(clk), .rst(
        n8) );
  dff_183 \writedata_reg[9]  ( .q(\WriteData<9> ), .d(n110), .clk(clk), .rst(
        n8) );
  dff_184 \writedata_reg[10]  ( .q(\WriteData<10> ), .d(n111), .clk(clk), 
        .rst(n8) );
  dff_185 \writedata_reg[11]  ( .q(\WriteData<11> ), .d(n112), .clk(clk), 
        .rst(n8) );
  dff_186 \writedata_reg[12]  ( .q(\WriteData<12> ), .d(n113), .clk(clk), 
        .rst(n8) );
  dff_187 \writedata_reg[13]  ( .q(\WriteData<13> ), .d(n114), .clk(clk), 
        .rst(n8) );
  dff_188 \writedata_reg[14]  ( .q(\WriteData<14> ), .d(n115), .clk(clk), 
        .rst(n8) );
  dff_189 \writedata_reg[15]  ( .q(\WriteData<15> ), .d(n116), .clk(clk), 
        .rst(n8) );
  dff_218 halt_reg ( .q(Halt_Out), .d(n120), .clk(clk), .rst(n8) );
  INVX1 U1 ( .A(rst), .Y(n9) );
  INVX1 U2 ( .A(n121), .Y(n6) );
  INVX1 U3 ( .A(n9), .Y(n7) );
  INVX1 U4 ( .A(\Address<10> ), .Y(n20) );
  INVX1 U5 ( .A(n123), .Y(n2) );
  INVX1 U6 ( .A(n122), .Y(n4) );
  INVX1 U7 ( .A(n6), .Y(\Address<4> ) );
  INVX1 U8 ( .A(\Address<5> ), .Y(n30) );
  INVX1 U9 ( .A(\Address<6> ), .Y(n28) );
  INVX1 U10 ( .A(\Address<7> ), .Y(n26) );
  INVX1 U11 ( .A(\Address<8> ), .Y(n24) );
  INVX1 U12 ( .A(\Address<9> ), .Y(n22) );
  INVX1 U13 ( .A(\Address<11> ), .Y(n18) );
  INVX1 U14 ( .A(\Address<12> ), .Y(n16) );
  INVX1 U15 ( .A(\Address<13> ), .Y(n14) );
  INVX1 U16 ( .A(\Address<14> ), .Y(n12) );
  INVX1 U17 ( .A(\Address<15> ), .Y(n10) );
  INVX1 U18 ( .A(Stall), .Y(n37) );
  INVX1 U19 ( .A(n9), .Y(n8) );
  INVX1 U20 ( .A(n100), .Y(n101) );
  INVX1 U21 ( .A(n99), .Y(n111) );
  INVX1 U22 ( .A(n98), .Y(n112) );
  INVX1 U23 ( .A(n97), .Y(n113) );
  INVX1 U24 ( .A(n96), .Y(n114) );
  INVX1 U25 ( .A(n95), .Y(n115) );
  INVX1 U26 ( .A(n94), .Y(n116) );
  INVX1 U27 ( .A(n93), .Y(n102) );
  INVX1 U28 ( .A(n92), .Y(n103) );
  INVX1 U29 ( .A(n91), .Y(n104) );
  INVX1 U30 ( .A(n90), .Y(n105) );
  INVX1 U31 ( .A(n89), .Y(n106) );
  INVX1 U32 ( .A(n88), .Y(n107) );
  INVX1 U33 ( .A(n87), .Y(n108) );
  INVX1 U34 ( .A(n86), .Y(n109) );
  INVX1 U35 ( .A(n85), .Y(n110) );
  INVX1 U36 ( .A(n77), .Y(n70) );
  INVX1 U37 ( .A(n68), .Y(n120) );
  INVX1 U38 ( .A(n67), .Y(n118) );
  INVX1 U39 ( .A(n66), .Y(n119) );
  INVX1 U40 ( .A(n65), .Y(n117) );
  INVX1 U41 ( .A(n64), .Y(n82) );
  INVX1 U42 ( .A(n63), .Y(n83) );
  INVX1 U43 ( .A(n62), .Y(n84) );
  INVX1 U44 ( .A(n61), .Y(n74) );
  INVX1 U45 ( .A(n60), .Y(n75) );
  INVX1 U46 ( .A(n59), .Y(n76) );
  INVX1 U47 ( .A(n58), .Y(n78) );
  INVX1 U48 ( .A(n57), .Y(n79) );
  INVX1 U49 ( .A(n56), .Y(n80) );
  INVX1 U50 ( .A(n55), .Y(n81) );
  INVX1 U68 ( .A(n54), .Y(n71) );
  INVX1 U69 ( .A(n53), .Y(n72) );
  INVX1 U70 ( .A(n52), .Y(n73) );
  INVX1 U71 ( .A(n2), .Y(\Address<2> ) );
  INVX1 U72 ( .A(n4), .Y(\Address<3> ) );
  INVX1 U73 ( .A(\Result<2> ), .Y(n34) );
  INVX1 U74 ( .A(\Result<3> ), .Y(n33) );
  INVX1 U75 ( .A(\Result<4> ), .Y(n32) );
  INVX1 U77 ( .A(\Result<5> ), .Y(n31) );
  INVX1 U78 ( .A(\Result<6> ), .Y(n29) );
  INVX1 U79 ( .A(\Result<7> ), .Y(n27) );
  INVX1 U80 ( .A(\Result<8> ), .Y(n25) );
  INVX1 U81 ( .A(\Result<9> ), .Y(n23) );
  INVX1 U82 ( .A(\Result<10> ), .Y(n21) );
  INVX1 U83 ( .A(\Result<11> ), .Y(n19) );
  INVX1 U100 ( .A(\Result<12> ), .Y(n17) );
  INVX1 U101 ( .A(\Result<13> ), .Y(n15) );
  INVX1 U102 ( .A(\Result<14> ), .Y(n13) );
  INVX1 U103 ( .A(\Result<15> ), .Y(n11) );
  OAI21X1 U104 ( .A(n36), .B(Stall), .C(n35), .Y(n38) );
  INVX1 U105 ( .A(\Result<0> ), .Y(n36) );
  MUX2X1 U106 ( .B(n11), .A(n10), .S(Stall), .Y(n69) );
  MUX2X1 U107 ( .B(n13), .A(n12), .S(Stall), .Y(n51) );
  MUX2X1 U108 ( .B(n15), .A(n14), .S(Stall), .Y(n50) );
  MUX2X1 U109 ( .B(n17), .A(n16), .S(Stall), .Y(n49) );
  MUX2X1 U110 ( .B(n19), .A(n18), .S(Stall), .Y(n48) );
  MUX2X1 U111 ( .B(n21), .A(n20), .S(Stall), .Y(n47) );
  MUX2X1 U112 ( .B(n23), .A(n22), .S(Stall), .Y(n46) );
  MUX2X1 U113 ( .B(n25), .A(n24), .S(Stall), .Y(n45) );
  MUX2X1 U114 ( .B(n27), .A(n26), .S(Stall), .Y(n44) );
  MUX2X1 U115 ( .B(n29), .A(n28), .S(Stall), .Y(n43) );
  MUX2X1 U116 ( .B(n31), .A(n30), .S(Stall), .Y(n42) );
  MUX2X1 U117 ( .B(n32), .A(n6), .S(Stall), .Y(n41) );
  MUX2X1 U118 ( .B(n33), .A(n4), .S(Stall), .Y(n40) );
  MUX2X1 U119 ( .B(n34), .A(n2), .S(Stall), .Y(n39) );
  NAND2X1 U120 ( .A(\Address<0> ), .B(Stall), .Y(n35) );
endmodule


module memory ( MemRead, MemWrite, halt, clk, rst, .Address({\Address<15> , 
        \Address<14> , \Address<13> , \Address<12> , \Address<11> , 
        \Address<10> , \Address<9> , \Address<8> , \Address<7> , \Address<6> , 
        \Address<5> , \Address<4> , \Address<3> , \Address<2> , \Address<1> , 
        \Address<0> }), .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }), .ReadData({\ReadData<15> , 
        \ReadData<14> , \ReadData<13> , \ReadData<12> , \ReadData<11> , 
        \ReadData<10> , \ReadData<9> , \ReadData<8> , \ReadData<7> , 
        \ReadData<6> , \ReadData<5> , \ReadData<4> , \ReadData<3> , 
        \ReadData<2> , \ReadData<1> , \ReadData<0> }) );
  input MemRead, MemWrite, halt, clk, rst, \Address<15> , \Address<14> ,
         \Address<13> , \Address<12> , \Address<11> , \Address<10> ,
         \Address<9> , \Address<8> , \Address<7> , \Address<6> , \Address<5> ,
         \Address<4> , \Address<3> , \Address<2> , \Address<1> , \Address<0> ,
         \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ;
  output \ReadData<15> , \ReadData<14> , \ReadData<13> , \ReadData<12> ,
         \ReadData<11> , \ReadData<10> , \ReadData<9> , \ReadData<8> ,
         \ReadData<7> , \ReadData<6> , \ReadData<5> , \ReadData<4> ,
         \ReadData<3> , \ReadData<2> , \ReadData<1> , \ReadData<0> ;
  wire   n1;

  memory2c_0 data_mem ( .data_out({\ReadData<15> , \ReadData<14> , 
        \ReadData<13> , \ReadData<12> , \ReadData<11> , \ReadData<10> , 
        \ReadData<9> , \ReadData<8> , \ReadData<7> , \ReadData<6> , 
        \ReadData<5> , \ReadData<4> , \ReadData<3> , \ReadData<2> , 
        \ReadData<1> , \ReadData<0> }), .data_in({\WriteData<15> , 
        \WriteData<14> , \WriteData<13> , \WriteData<12> , \WriteData<11> , 
        \WriteData<10> , \WriteData<9> , \WriteData<8> , \WriteData<7> , 
        \WriteData<6> , \WriteData<5> , \WriteData<4> , \WriteData<3> , 
        \WriteData<2> , \WriteData<1> , \WriteData<0> }), .addr({\Address<15> , 
        \Address<14> , \Address<13> , \Address<12> , \Address<11> , 
        \Address<10> , \Address<9> , \Address<8> , \Address<7> , \Address<6> , 
        \Address<5> , \Address<4> , \Address<3> , \Address<2> , \Address<1> , 
        \Address<0> }), .enable(n1), .wr(MemWrite), .createdump(halt), .clk(
        clk), .rst(rst) );
  INVX1 U1 ( .A(halt), .Y(n1) );
endmodule


module pipe_mw ( Stall, rst, clk, .ExecuteOut({\ExecuteOut<15> , 
        \ExecuteOut<14> , \ExecuteOut<13> , \ExecuteOut<12> , \ExecuteOut<11> , 
        \ExecuteOut<10> , \ExecuteOut<9> , \ExecuteOut<8> , \ExecuteOut<7> , 
        \ExecuteOut<6> , \ExecuteOut<5> , \ExecuteOut<4> , \ExecuteOut<3> , 
        \ExecuteOut<2> , \ExecuteOut<1> , \ExecuteOut<0> }), .MemOut({
        \MemOut<15> , \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> , 
        \MemOut<10> , \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> , 
        \MemOut<5> , \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> , 
        \MemOut<0> }), MemToReg, RegFileWrEn, .Rs({\Rs<2> , \Rs<1> , \Rs<0> }), 
    .Rt({\Rt<2> , \Rt<1> , \Rt<0> }), .Rd({\Rd<2> , \Rd<1> , \Rd<0> }), 
    .WriteReg({\WriteReg<2> , \WriteReg<1> , \WriteReg<0> }), 
    .ExecuteOut_Out({\ExecuteOut_Out<15> , \ExecuteOut_Out<14> , 
        \ExecuteOut_Out<13> , \ExecuteOut_Out<12> , \ExecuteOut_Out<11> , 
        \ExecuteOut_Out<10> , \ExecuteOut_Out<9> , \ExecuteOut_Out<8> , 
        \ExecuteOut_Out<7> , \ExecuteOut_Out<6> , \ExecuteOut_Out<5> , 
        \ExecuteOut_Out<4> , \ExecuteOut_Out<3> , \ExecuteOut_Out<2> , 
        \ExecuteOut_Out<1> , \ExecuteOut_Out<0> }), .MemOut_Out({
        \MemOut_Out<15> , \MemOut_Out<14> , \MemOut_Out<13> , \MemOut_Out<12> , 
        \MemOut_Out<11> , \MemOut_Out<10> , \MemOut_Out<9> , \MemOut_Out<8> , 
        \MemOut_Out<7> , \MemOut_Out<6> , \MemOut_Out<5> , \MemOut_Out<4> , 
        \MemOut_Out<3> , \MemOut_Out<2> , \MemOut_Out<1> , \MemOut_Out<0> }), 
        MemToReg_Out, RegFileWrEn_Out, .WriteReg_Out({\WriteReg_Out<2> , 
        \WriteReg_Out<1> , \WriteReg_Out<0> }), .Rs_Out({\Rs_Out<2> , 
        \Rs_Out<1> , \Rs_Out<0> }), .Rt_Out({\Rt_Out<2> , \Rt_Out<1> , 
        \Rt_Out<0> }), .Rd_Out({\Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> }) );
  input Stall, rst, clk, \ExecuteOut<15> , \ExecuteOut<14> , \ExecuteOut<13> ,
         \ExecuteOut<12> , \ExecuteOut<11> , \ExecuteOut<10> , \ExecuteOut<9> ,
         \ExecuteOut<8> , \ExecuteOut<7> , \ExecuteOut<6> , \ExecuteOut<5> ,
         \ExecuteOut<4> , \ExecuteOut<3> , \ExecuteOut<2> , \ExecuteOut<1> ,
         \ExecuteOut<0> , \MemOut<15> , \MemOut<14> , \MemOut<13> ,
         \MemOut<12> , \MemOut<11> , \MemOut<10> , \MemOut<9> , \MemOut<8> ,
         \MemOut<7> , \MemOut<6> , \MemOut<5> , \MemOut<4> , \MemOut<3> ,
         \MemOut<2> , \MemOut<1> , \MemOut<0> , MemToReg, RegFileWrEn, \Rs<2> ,
         \Rs<1> , \Rs<0> , \Rt<2> , \Rt<1> , \Rt<0> , \Rd<2> , \Rd<1> ,
         \Rd<0> , \WriteReg<2> , \WriteReg<1> , \WriteReg<0> ;
  output \ExecuteOut_Out<15> , \ExecuteOut_Out<14> , \ExecuteOut_Out<13> ,
         \ExecuteOut_Out<12> , \ExecuteOut_Out<11> , \ExecuteOut_Out<10> ,
         \ExecuteOut_Out<9> , \ExecuteOut_Out<8> , \ExecuteOut_Out<7> ,
         \ExecuteOut_Out<6> , \ExecuteOut_Out<5> , \ExecuteOut_Out<4> ,
         \ExecuteOut_Out<3> , \ExecuteOut_Out<2> , \ExecuteOut_Out<1> ,
         \ExecuteOut_Out<0> , \MemOut_Out<15> , \MemOut_Out<14> ,
         \MemOut_Out<13> , \MemOut_Out<12> , \MemOut_Out<11> ,
         \MemOut_Out<10> , \MemOut_Out<9> , \MemOut_Out<8> , \MemOut_Out<7> ,
         \MemOut_Out<6> , \MemOut_Out<5> , \MemOut_Out<4> , \MemOut_Out<3> ,
         \MemOut_Out<2> , \MemOut_Out<1> , \MemOut_Out<0> , MemToReg_Out,
         RegFileWrEn_Out, \WriteReg_Out<2> , \WriteReg_Out<1> ,
         \WriteReg_Out<0> , \Rs_Out<2> , \Rs_Out<1> , \Rs_Out<0> , \Rt_Out<2> ,
         \Rt_Out<1> , \Rt_Out<0> , \Rd_Out<2> , \Rd_Out<1> , \Rd_Out<0> ;
  wire   n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n95, n96, n97;

  AOI22X1 U48 ( .A(\WriteReg<2> ), .B(n97), .C(\WriteReg_Out<2> ), .D(Stall), 
        .Y(n49) );
  AOI22X1 U49 ( .A(\WriteReg<1> ), .B(n97), .C(\WriteReg_Out<1> ), .D(Stall), 
        .Y(n50) );
  AOI22X1 U50 ( .A(\WriteReg<0> ), .B(n97), .C(\WriteReg_Out<0> ), .D(Stall), 
        .Y(n51) );
  AOI22X1 U51 ( .A(\Rt<2> ), .B(n97), .C(\Rt_Out<2> ), .D(Stall), .Y(n52) );
  AOI22X1 U52 ( .A(\Rt<1> ), .B(n97), .C(\Rt_Out<1> ), .D(Stall), .Y(n53) );
  AOI22X1 U53 ( .A(\Rt<0> ), .B(n97), .C(\Rt_Out<0> ), .D(Stall), .Y(n54) );
  AOI22X1 U54 ( .A(\Rs<2> ), .B(n97), .C(\Rs_Out<2> ), .D(Stall), .Y(n55) );
  AOI22X1 U55 ( .A(\Rs<1> ), .B(n97), .C(\Rs_Out<1> ), .D(Stall), .Y(n56) );
  AOI22X1 U56 ( .A(\Rs<0> ), .B(n97), .C(\Rs_Out<0> ), .D(Stall), .Y(n57) );
  AOI22X1 U57 ( .A(RegFileWrEn), .B(n97), .C(RegFileWrEn_Out), .D(Stall), .Y(
        n58) );
  AOI22X1 U58 ( .A(\Rd<2> ), .B(n97), .C(\Rd_Out<2> ), .D(Stall), .Y(n59) );
  AOI22X1 U59 ( .A(\Rd<1> ), .B(n97), .C(\Rd_Out<1> ), .D(Stall), .Y(n60) );
  AOI22X1 U60 ( .A(\Rd<0> ), .B(n97), .C(\Rd_Out<0> ), .D(Stall), .Y(n61) );
  AOI22X1 U61 ( .A(MemToReg), .B(n97), .C(MemToReg_Out), .D(Stall), .Y(n62) );
  AOI22X1 U62 ( .A(\MemOut<9> ), .B(n97), .C(\MemOut_Out<9> ), .D(Stall), .Y(
        n63) );
  AOI22X1 U63 ( .A(\MemOut<8> ), .B(n97), .C(\MemOut_Out<8> ), .D(Stall), .Y(
        n64) );
  AOI22X1 U64 ( .A(\MemOut<7> ), .B(n97), .C(\MemOut_Out<7> ), .D(Stall), .Y(
        n65) );
  AOI22X1 U65 ( .A(\MemOut<6> ), .B(n97), .C(\MemOut_Out<6> ), .D(Stall), .Y(
        n66) );
  AOI22X1 U66 ( .A(\MemOut<5> ), .B(n97), .C(\MemOut_Out<5> ), .D(Stall), .Y(
        n67) );
  AOI22X1 U67 ( .A(\MemOut<4> ), .B(n97), .C(\MemOut_Out<4> ), .D(Stall), .Y(
        n68) );
  AOI22X1 U68 ( .A(\MemOut<3> ), .B(n97), .C(\MemOut_Out<3> ), .D(Stall), .Y(
        n69) );
  AOI22X1 U69 ( .A(\MemOut<2> ), .B(n97), .C(\MemOut_Out<2> ), .D(Stall), .Y(
        n70) );
  AOI22X1 U70 ( .A(\MemOut<1> ), .B(n97), .C(\MemOut_Out<1> ), .D(Stall), .Y(
        n71) );
  AOI22X1 U71 ( .A(\MemOut<15> ), .B(n97), .C(\MemOut_Out<15> ), .D(Stall), 
        .Y(n72) );
  AOI22X1 U72 ( .A(\MemOut<14> ), .B(n97), .C(\MemOut_Out<14> ), .D(Stall), 
        .Y(n73) );
  AOI22X1 U73 ( .A(\MemOut<13> ), .B(n97), .C(\MemOut_Out<13> ), .D(Stall), 
        .Y(n74) );
  AOI22X1 U74 ( .A(\MemOut<12> ), .B(n97), .C(\MemOut_Out<12> ), .D(Stall), 
        .Y(n75) );
  AOI22X1 U75 ( .A(\MemOut<11> ), .B(n97), .C(\MemOut_Out<11> ), .D(Stall), 
        .Y(n76) );
  AOI22X1 U76 ( .A(\MemOut<10> ), .B(n97), .C(\MemOut_Out<10> ), .D(Stall), 
        .Y(n77) );
  AOI22X1 U77 ( .A(\MemOut<0> ), .B(n97), .C(\MemOut_Out<0> ), .D(Stall), .Y(
        n78) );
  AOI22X1 U78 ( .A(\ExecuteOut<9> ), .B(n97), .C(\ExecuteOut_Out<9> ), .D(
        Stall), .Y(n79) );
  AOI22X1 U79 ( .A(\ExecuteOut<8> ), .B(n97), .C(\ExecuteOut_Out<8> ), .D(
        Stall), .Y(n80) );
  AOI22X1 U80 ( .A(\ExecuteOut<7> ), .B(n97), .C(\ExecuteOut_Out<7> ), .D(
        Stall), .Y(n81) );
  AOI22X1 U81 ( .A(\ExecuteOut<6> ), .B(n97), .C(\ExecuteOut_Out<6> ), .D(
        Stall), .Y(n82) );
  AOI22X1 U82 ( .A(\ExecuteOut<5> ), .B(n97), .C(\ExecuteOut_Out<5> ), .D(
        Stall), .Y(n83) );
  AOI22X1 U83 ( .A(\ExecuteOut<4> ), .B(n97), .C(\ExecuteOut_Out<4> ), .D(
        Stall), .Y(n84) );
  AOI22X1 U84 ( .A(\ExecuteOut<3> ), .B(n97), .C(\ExecuteOut_Out<3> ), .D(
        Stall), .Y(n85) );
  AOI22X1 U85 ( .A(\ExecuteOut<2> ), .B(n97), .C(\ExecuteOut_Out<2> ), .D(
        Stall), .Y(n86) );
  AOI22X1 U86 ( .A(\ExecuteOut<1> ), .B(n97), .C(\ExecuteOut_Out<1> ), .D(
        Stall), .Y(n87) );
  AOI22X1 U87 ( .A(\ExecuteOut<15> ), .B(n97), .C(\ExecuteOut_Out<15> ), .D(
        Stall), .Y(n88) );
  AOI22X1 U88 ( .A(\ExecuteOut<14> ), .B(n97), .C(\ExecuteOut_Out<14> ), .D(
        Stall), .Y(n89) );
  AOI22X1 U89 ( .A(\ExecuteOut<13> ), .B(n97), .C(\ExecuteOut_Out<13> ), .D(
        Stall), .Y(n90) );
  AOI22X1 U90 ( .A(\ExecuteOut<12> ), .B(n97), .C(\ExecuteOut_Out<12> ), .D(
        Stall), .Y(n91) );
  AOI22X1 U91 ( .A(\ExecuteOut<11> ), .B(n97), .C(\ExecuteOut_Out<11> ), .D(
        Stall), .Y(n92) );
  AOI22X1 U92 ( .A(\ExecuteOut<10> ), .B(n97), .C(\ExecuteOut_Out<10> ), .D(
        Stall), .Y(n93) );
  AOI22X1 U93 ( .A(\ExecuteOut<0> ), .B(n97), .C(\ExecuteOut_Out<0> ), .D(
        Stall), .Y(n94) );
  dff_169 \WriteReg_reg[0]  ( .q(\WriteReg_Out<0> ), .d(n21), .clk(clk), .rst(
        n3) );
  dff_170 \WriteReg_reg[1]  ( .q(\WriteReg_Out<1> ), .d(n22), .clk(clk), .rst(
        n3) );
  dff_171 \WriteReg_reg[2]  ( .q(\WriteReg_Out<2> ), .d(n23), .clk(clk), .rst(
        n3) );
  dff_166 \rs_reg[0]  ( .q(\Rs_Out<0> ), .d(n24), .clk(clk), .rst(n3) );
  dff_167 \rs_reg[1]  ( .q(\Rs_Out<1> ), .d(n25), .clk(clk), .rst(n3) );
  dff_168 \rs_reg[2]  ( .q(\Rs_Out<2> ), .d(n26), .clk(clk), .rst(n3) );
  dff_163 \rt_reg[0]  ( .q(\Rt_Out<0> ), .d(n27), .clk(clk), .rst(n3) );
  dff_164 \rt_reg[1]  ( .q(\Rt_Out<1> ), .d(n28), .clk(clk), .rst(n2) );
  dff_165 \rt_reg[2]  ( .q(\Rt_Out<2> ), .d(n29), .clk(clk), .rst(n2) );
  dff_160 \rd_reg[0]  ( .q(\Rd_Out<0> ), .d(n30), .clk(clk), .rst(n2) );
  dff_161 \rd_reg[1]  ( .q(\Rd_Out<1> ), .d(n31), .clk(clk), .rst(n2) );
  dff_162 \rd_reg[2]  ( .q(\Rd_Out<2> ), .d(n32), .clk(clk), .rst(n2) );
  dff_173 rf_wr_en_reg ( .q(RegFileWrEn_Out), .d(n33), .clk(clk), .rst(n2) );
  dff_144 \executeout_reg[0]  ( .q(\ExecuteOut_Out<0> ), .d(n34), .clk(clk), 
        .rst(n2) );
  dff_145 \executeout_reg[1]  ( .q(\ExecuteOut_Out<1> ), .d(n35), .clk(clk), 
        .rst(n2) );
  dff_146 \executeout_reg[2]  ( .q(\ExecuteOut_Out<2> ), .d(n36), .clk(clk), 
        .rst(n2) );
  dff_147 \executeout_reg[3]  ( .q(\ExecuteOut_Out<3> ), .d(n37), .clk(clk), 
        .rst(n2) );
  dff_148 \executeout_reg[4]  ( .q(\ExecuteOut_Out<4> ), .d(n38), .clk(clk), 
        .rst(n2) );
  dff_149 \executeout_reg[5]  ( .q(\ExecuteOut_Out<5> ), .d(n39), .clk(clk), 
        .rst(n2) );
  dff_150 \executeout_reg[6]  ( .q(\ExecuteOut_Out<6> ), .d(n40), .clk(clk), 
        .rst(n2) );
  dff_151 \executeout_reg[7]  ( .q(\ExecuteOut_Out<7> ), .d(n41), .clk(clk), 
        .rst(n1) );
  dff_152 \executeout_reg[8]  ( .q(\ExecuteOut_Out<8> ), .d(n42), .clk(clk), 
        .rst(n1) );
  dff_153 \executeout_reg[9]  ( .q(\ExecuteOut_Out<9> ), .d(n43), .clk(clk), 
        .rst(n1) );
  dff_154 \executeout_reg[10]  ( .q(\ExecuteOut_Out<10> ), .d(n44), .clk(clk), 
        .rst(n1) );
  dff_155 \executeout_reg[11]  ( .q(\ExecuteOut_Out<11> ), .d(n45), .clk(clk), 
        .rst(n1) );
  dff_156 \executeout_reg[12]  ( .q(\ExecuteOut_Out<12> ), .d(n46), .clk(clk), 
        .rst(n1) );
  dff_157 \executeout_reg[13]  ( .q(\ExecuteOut_Out<13> ), .d(n47), .clk(clk), 
        .rst(n1) );
  dff_158 \executeout_reg[14]  ( .q(\ExecuteOut_Out<14> ), .d(n48), .clk(clk), 
        .rst(n1) );
  dff_159 \executeout_reg[15]  ( .q(\ExecuteOut_Out<15> ), .d(n95), .clk(clk), 
        .rst(n1) );
  dff_128 \memout_reg[0]  ( .q(\MemOut_Out<0> ), .d(n20), .clk(clk), .rst(n1)
         );
  dff_129 \memout_reg[1]  ( .q(\MemOut_Out<1> ), .d(n18), .clk(clk), .rst(n1)
         );
  dff_130 \memout_reg[2]  ( .q(\MemOut_Out<2> ), .d(n16), .clk(clk), .rst(n1)
         );
  dff_131 \memout_reg[3]  ( .q(\MemOut_Out<3> ), .d(n14), .clk(clk), .rst(n1)
         );
  dff_132 \memout_reg[4]  ( .q(\MemOut_Out<4> ), .d(n12), .clk(clk), .rst(n3)
         );
  dff_133 \memout_reg[5]  ( .q(\MemOut_Out<5> ), .d(n10), .clk(clk), .rst(n3)
         );
  dff_134 \memout_reg[6]  ( .q(\MemOut_Out<6> ), .d(n8), .clk(clk), .rst(n3)
         );
  dff_135 \memout_reg[7]  ( .q(\MemOut_Out<7> ), .d(n6), .clk(clk), .rst(n3)
         );
  dff_136 \memout_reg[8]  ( .q(\MemOut_Out<8> ), .d(n19), .clk(clk), .rst(n3)
         );
  dff_137 \memout_reg[9]  ( .q(\MemOut_Out<9> ), .d(n17), .clk(clk), .rst(n3)
         );
  dff_138 \memout_reg[10]  ( .q(\MemOut_Out<10> ), .d(n15), .clk(clk), .rst(
        rst) );
  dff_139 \memout_reg[11]  ( .q(\MemOut_Out<11> ), .d(n13), .clk(clk), .rst(
        rst) );
  dff_140 \memout_reg[12]  ( .q(\MemOut_Out<12> ), .d(n11), .clk(clk), .rst(
        rst) );
  dff_141 \memout_reg[13]  ( .q(\MemOut_Out<13> ), .d(n9), .clk(clk), .rst(rst) );
  dff_142 \memout_reg[14]  ( .q(\MemOut_Out<14> ), .d(n7), .clk(clk), .rst(rst) );
  dff_143 \memout_reg[15]  ( .q(\MemOut_Out<15> ), .d(n5), .clk(clk), .rst(rst) );
  dff_172 memtoreg_reg ( .q(MemToReg_Out), .d(n96), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(Stall), .Y(n97) );
  INVX1 U2 ( .A(n64), .Y(n19) );
  INVX1 U3 ( .A(n63), .Y(n17) );
  INVX1 U4 ( .A(n77), .Y(n15) );
  INVX1 U5 ( .A(n76), .Y(n13) );
  INVX1 U6 ( .A(n75), .Y(n11) );
  INVX1 U7 ( .A(n74), .Y(n9) );
  INVX1 U8 ( .A(n73), .Y(n7) );
  INVX1 U9 ( .A(n72), .Y(n5) );
  INVX1 U10 ( .A(rst), .Y(n4) );
  INVX1 U11 ( .A(n4), .Y(n1) );
  INVX1 U12 ( .A(n4), .Y(n2) );
  INVX1 U13 ( .A(n4), .Y(n3) );
  INVX1 U14 ( .A(n94), .Y(n34) );
  INVX1 U15 ( .A(n93), .Y(n44) );
  INVX1 U16 ( .A(n92), .Y(n45) );
  INVX1 U17 ( .A(n91), .Y(n46) );
  INVX1 U18 ( .A(n90), .Y(n47) );
  INVX1 U19 ( .A(n89), .Y(n48) );
  INVX1 U20 ( .A(n88), .Y(n95) );
  INVX1 U21 ( .A(n87), .Y(n35) );
  INVX1 U22 ( .A(n86), .Y(n36) );
  INVX1 U23 ( .A(n85), .Y(n37) );
  INVX1 U24 ( .A(n84), .Y(n38) );
  INVX1 U25 ( .A(n83), .Y(n39) );
  INVX1 U26 ( .A(n82), .Y(n40) );
  INVX1 U27 ( .A(n81), .Y(n41) );
  INVX1 U28 ( .A(n80), .Y(n42) );
  INVX1 U29 ( .A(n79), .Y(n43) );
  INVX1 U30 ( .A(n78), .Y(n20) );
  INVX1 U31 ( .A(n71), .Y(n18) );
  INVX1 U32 ( .A(n70), .Y(n16) );
  INVX1 U33 ( .A(n69), .Y(n14) );
  INVX1 U34 ( .A(n68), .Y(n12) );
  INVX1 U35 ( .A(n67), .Y(n10) );
  INVX1 U36 ( .A(n66), .Y(n8) );
  INVX1 U37 ( .A(n65), .Y(n6) );
  INVX1 U38 ( .A(n62), .Y(n96) );
  INVX1 U39 ( .A(n61), .Y(n30) );
  INVX1 U40 ( .A(n60), .Y(n31) );
  INVX1 U41 ( .A(n59), .Y(n32) );
  INVX1 U42 ( .A(n58), .Y(n33) );
  INVX1 U43 ( .A(n57), .Y(n24) );
  INVX1 U44 ( .A(n56), .Y(n25) );
  INVX1 U45 ( .A(n55), .Y(n26) );
  INVX1 U46 ( .A(n54), .Y(n27) );
  INVX1 U47 ( .A(n53), .Y(n28) );
  INVX1 U94 ( .A(n52), .Y(n29) );
  INVX1 U95 ( .A(n51), .Y(n21) );
  INVX1 U96 ( .A(n50), .Y(n22) );
  INVX1 U97 ( .A(n49), .Y(n23) );
endmodule


module writeback ( .ExecuteOut({\ExecuteOut<15> , \ExecuteOut<14> , 
        \ExecuteOut<13> , \ExecuteOut<12> , \ExecuteOut<11> , \ExecuteOut<10> , 
        \ExecuteOut<9> , \ExecuteOut<8> , \ExecuteOut<7> , \ExecuteOut<6> , 
        \ExecuteOut<5> , \ExecuteOut<4> , \ExecuteOut<3> , \ExecuteOut<2> , 
        \ExecuteOut<1> , \ExecuteOut<0> }), .MemOut({\MemOut<15> , 
        \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> , \MemOut<10> , 
        \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> , \MemOut<5> , 
        \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> , \MemOut<0> }), 
        MemToReg, .WriteData({\WriteData<15> , \WriteData<14> , 
        \WriteData<13> , \WriteData<12> , \WriteData<11> , \WriteData<10> , 
        \WriteData<9> , \WriteData<8> , \WriteData<7> , \WriteData<6> , 
        \WriteData<5> , \WriteData<4> , \WriteData<3> , \WriteData<2> , 
        \WriteData<1> , \WriteData<0> }) );
  input \ExecuteOut<15> , \ExecuteOut<14> , \ExecuteOut<13> , \ExecuteOut<12> ,
         \ExecuteOut<11> , \ExecuteOut<10> , \ExecuteOut<9> , \ExecuteOut<8> ,
         \ExecuteOut<7> , \ExecuteOut<6> , \ExecuteOut<5> , \ExecuteOut<4> ,
         \ExecuteOut<3> , \ExecuteOut<2> , \ExecuteOut<1> , \ExecuteOut<0> ,
         \MemOut<15> , \MemOut<14> , \MemOut<13> , \MemOut<12> , \MemOut<11> ,
         \MemOut<10> , \MemOut<9> , \MemOut<8> , \MemOut<7> , \MemOut<6> ,
         \MemOut<5> , \MemOut<4> , \MemOut<3> , \MemOut<2> , \MemOut<1> ,
         \MemOut<0> , MemToReg;
  output \WriteData<15> , \WriteData<14> , \WriteData<13> , \WriteData<12> ,
         \WriteData<11> , \WriteData<10> , \WriteData<9> , \WriteData<8> ,
         \WriteData<7> , \WriteData<6> , \WriteData<5> , \WriteData<4> ,
         \WriteData<3> , \WriteData<2> , \WriteData<1> , \WriteData<0> ;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n17;

  AOI22X1 U18 ( .A(\ExecuteOut<9> ), .B(n17), .C(MemToReg), .D(\MemOut<9> ), 
        .Y(n19) );
  AOI22X1 U19 ( .A(\ExecuteOut<8> ), .B(n17), .C(\MemOut<8> ), .D(MemToReg), 
        .Y(n20) );
  AOI22X1 U20 ( .A(\ExecuteOut<7> ), .B(n17), .C(\MemOut<7> ), .D(MemToReg), 
        .Y(n21) );
  AOI22X1 U21 ( .A(\ExecuteOut<6> ), .B(n17), .C(\MemOut<6> ), .D(MemToReg), 
        .Y(n22) );
  AOI22X1 U22 ( .A(\ExecuteOut<5> ), .B(n17), .C(\MemOut<5> ), .D(MemToReg), 
        .Y(n23) );
  AOI22X1 U23 ( .A(\ExecuteOut<4> ), .B(n17), .C(\MemOut<4> ), .D(MemToReg), 
        .Y(n24) );
  AOI22X1 U24 ( .A(\ExecuteOut<3> ), .B(n17), .C(\MemOut<3> ), .D(MemToReg), 
        .Y(n25) );
  AOI22X1 U25 ( .A(\ExecuteOut<2> ), .B(n17), .C(\MemOut<2> ), .D(MemToReg), 
        .Y(n26) );
  AOI22X1 U26 ( .A(\ExecuteOut<1> ), .B(n17), .C(\MemOut<1> ), .D(MemToReg), 
        .Y(n27) );
  AOI22X1 U27 ( .A(\ExecuteOut<15> ), .B(n17), .C(\MemOut<15> ), .D(MemToReg), 
        .Y(n28) );
  AOI22X1 U28 ( .A(\ExecuteOut<14> ), .B(n17), .C(\MemOut<14> ), .D(MemToReg), 
        .Y(n29) );
  AOI22X1 U29 ( .A(\ExecuteOut<13> ), .B(n17), .C(\MemOut<13> ), .D(MemToReg), 
        .Y(n30) );
  AOI22X1 U30 ( .A(\ExecuteOut<12> ), .B(n17), .C(\MemOut<12> ), .D(MemToReg), 
        .Y(n31) );
  AOI22X1 U31 ( .A(\ExecuteOut<11> ), .B(n17), .C(\MemOut<11> ), .D(MemToReg), 
        .Y(n32) );
  AOI22X1 U32 ( .A(\ExecuteOut<10> ), .B(n17), .C(\MemOut<10> ), .D(MemToReg), 
        .Y(n33) );
  AOI22X1 U33 ( .A(\ExecuteOut<0> ), .B(n17), .C(\MemOut<0> ), .D(MemToReg), 
        .Y(n34) );
  INVX1 U1 ( .A(n34), .Y(\WriteData<0> ) );
  INVX1 U2 ( .A(n33), .Y(\WriteData<10> ) );
  INVX1 U3 ( .A(n32), .Y(\WriteData<11> ) );
  INVX1 U4 ( .A(n31), .Y(\WriteData<12> ) );
  INVX1 U5 ( .A(n30), .Y(\WriteData<13> ) );
  INVX1 U6 ( .A(n29), .Y(\WriteData<14> ) );
  INVX1 U7 ( .A(n28), .Y(\WriteData<15> ) );
  INVX1 U8 ( .A(n27), .Y(\WriteData<1> ) );
  INVX1 U9 ( .A(n26), .Y(\WriteData<2> ) );
  INVX1 U10 ( .A(n25), .Y(\WriteData<3> ) );
  INVX1 U11 ( .A(n24), .Y(\WriteData<4> ) );
  INVX1 U12 ( .A(n23), .Y(\WriteData<5> ) );
  INVX1 U13 ( .A(n22), .Y(\WriteData<6> ) );
  INVX1 U14 ( .A(n21), .Y(\WriteData<7> ) );
  INVX1 U15 ( .A(n20), .Y(\WriteData<8> ) );
  INVX1 U16 ( .A(n19), .Y(\WriteData<9> ) );
  INVX1 U17 ( .A(MemToReg), .Y(n17) );
endmodule


module proc ( err, clk, rst );
  input clk, rst;
  output err;
  wire   E_BranchJumpTaken, D_RsValid, PDE_RegFileWrEn, \PDE_WriteReg<2> ,
         \PDE_WriteReg<1> , \PDE_WriteReg<0> , \D_Rs<2> , \D_Rs<1> , \D_Rs<0> ,
         D_RtValid, \D_Rt<2> , \D_Rt<1> , \D_Rt<0> , PEM_RegFileWrEn,
         \PEM_WriteReg<2> , \PEM_WriteReg<1> , \PEM_WriteReg<0> , D_RdValid,
         D_Store, \D_Rd<2> , \D_Rd<1> , \D_Rd<0> , \E_BranchPC<15> ,
         \E_BranchPC<14> , \E_BranchPC<13> , \E_BranchPC<12> ,
         \E_BranchPC<11> , \E_BranchPC<10> , \E_BranchPC<9> , \E_BranchPC<8> ,
         \E_BranchPC<7> , \E_BranchPC<6> , \E_BranchPC<5> , \E_BranchPC<4> ,
         \E_BranchPC<3> , \E_BranchPC<2> , \E_BranchPC<1> , \E_BranchPC<0> ,
         PEM_Halt, D_Exception, D_Rti, \F_Instr<15> , \F_Instr<14> ,
         \F_Instr<13> , \F_Instr<12> , \F_Instr<11> , \F_Instr<10> ,
         \F_Instr<9> , \F_Instr<8> , \F_Instr<7> , \F_Instr<6> , \F_Instr<5> ,
         \F_Instr<4> , \F_Instr<3> , \F_Instr<2> , \F_Instr<1> , \F_Instr<0> ,
         \F_IncPC<15> , \F_IncPC<14> , \F_IncPC<13> , \F_IncPC<12> ,
         \F_IncPC<11> , \F_IncPC<10> , \F_IncPC<9> , \F_IncPC<8> ,
         \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , \F_IncPC<4> , \F_IncPC<3> ,
         \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> , _2_net_, \PFD_Instr<15> ,
         \PFD_Instr<14> , \PFD_Instr<13> , \PFD_Instr<12> , \PFD_Instr<11> ,
         \PFD_Instr<10> , \PFD_Instr<9> , \PFD_Instr<8> , \PFD_Instr<7> ,
         \PFD_Instr<6> , \PFD_Instr<5> , \PFD_Instr<4> , \PFD_Instr<3> ,
         \PFD_Instr<2> , \PFD_Instr<1> , \PFD_Instr<0> , \PFD_IncPC<15> ,
         \PFD_IncPC<14> , \PFD_IncPC<13> , \PFD_IncPC<12> , \PFD_IncPC<11> ,
         \PFD_IncPC<10> , \PFD_IncPC<9> , \PFD_IncPC<8> , \PFD_IncPC<7> ,
         \PFD_IncPC<6> , \PFD_IncPC<5> , \PFD_IncPC<4> , \PFD_IncPC<3> ,
         \PFD_IncPC<2> , \PFD_IncPC<1> , \PFD_IncPC<0> , PFD_CPUActive,
         \W_WriteData<15> , \W_WriteData<14> , \W_WriteData<13> ,
         \W_WriteData<12> , \W_WriteData<11> , \W_WriteData<10> ,
         \W_WriteData<9> , \W_WriteData<8> , \W_WriteData<7> ,
         \W_WriteData<6> , \W_WriteData<5> , \W_WriteData<4> ,
         \W_WriteData<3> , \W_WriteData<2> , \W_WriteData<1> ,
         \W_WriteData<0> , \D_ALUOp1<15> , \D_ALUOp1<14> , \D_ALUOp1<13> ,
         \D_ALUOp1<12> , \D_ALUOp1<11> , \D_ALUOp1<10> , \D_ALUOp1<9> ,
         \D_ALUOp1<8> , \D_ALUOp1<7> , \D_ALUOp1<6> , \D_ALUOp1<5> ,
         \D_ALUOp1<4> , \D_ALUOp1<3> , \D_ALUOp1<2> , \D_ALUOp1<1> ,
         \D_ALUOp1<0> , \D_ALUOp2<15> , \D_ALUOp2<14> , \D_ALUOp2<13> ,
         \D_ALUOp2<12> , \D_ALUOp2<11> , \D_ALUOp2<10> , \D_ALUOp2<9> ,
         \D_ALUOp2<8> , \D_ALUOp2<7> , \D_ALUOp2<6> , \D_ALUOp2<5> ,
         \D_ALUOp2<4> , \D_ALUOp2<3> , \D_ALUOp2<2> , \D_ALUOp2<1> ,
         \D_ALUOp2<0> , D_ALUSrc, D_Branch, D_Jump, D_JumpReg, D_Set, D_Btr,
         \D_ALUOpcode<2> , \D_ALUOpcode<1> , \D_ALUOpcode<0> , \D_Func<1> ,
         \D_Func<0> , D_MemWrite, D_MemRead, D_MemToReg, D_Halt,
         \D_Immediate<15> , \D_Immediate<14> , \D_Immediate<13> ,
         \D_Immediate<12> , \D_Immediate<11> , \D_Immediate<10> ,
         \D_Immediate<9> , \D_Immediate<8> , \D_Immediate<7> ,
         \D_Immediate<6> , \D_Immediate<5> , \D_Immediate<4> ,
         \D_Immediate<3> , \D_Immediate<2> , \D_Immediate<1> ,
         \D_Immediate<0> , D_InvA, D_InvB, D_Cin, PMW_RegFileWrEn,
         D_RegFileWrEn, \PMW_WriteReg<2> , \PMW_WriteReg<1> ,
         \PMW_WriteReg<0> , \D_WriteReg<2> , \D_WriteReg<1> , \D_WriteReg<0> ,
         D_Link, _3_net_, \_5_net_<0> , _6_net_, _7_net_, _8_net_, _9_net_,
         _10_net_, _11_net_, _12_net_, _14_net_, _15_net_, _16_net_, _17_net_,
         _18_net_, \PDE_IncPC<15> , \PDE_IncPC<14> , \PDE_IncPC<13> ,
         \PDE_IncPC<12> , \PDE_IncPC<11> , \PDE_IncPC<10> , \PDE_IncPC<9> ,
         \PDE_IncPC<8> , \PDE_IncPC<7> , \PDE_IncPC<6> , \PDE_IncPC<5> ,
         \PDE_IncPC<4> , \PDE_IncPC<3> , \PDE_IncPC<2> , \PDE_IncPC<1> ,
         \PDE_IncPC<0> , \PDE_ALUOp1<15> , \PDE_ALUOp1<14> , \PDE_ALUOp1<13> ,
         \PDE_ALUOp1<12> , \PDE_ALUOp1<11> , \PDE_ALUOp1<10> , \PDE_ALUOp1<9> ,
         \PDE_ALUOp1<8> , \PDE_ALUOp1<7> , \PDE_ALUOp1<6> , \PDE_ALUOp1<5> ,
         \PDE_ALUOp1<4> , \PDE_ALUOp1<3> , \PDE_ALUOp1<2> , \PDE_ALUOp1<1> ,
         \PDE_ALUOp1<0> , \PDE_ALUOp2<15> , \PDE_ALUOp2<14> , \PDE_ALUOp2<13> ,
         \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , \PDE_ALUOp2<10> , \PDE_ALUOp2<9> ,
         \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , \PDE_ALUOp2<6> , \PDE_ALUOp2<5> ,
         \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , \PDE_ALUOp2<2> , \PDE_ALUOp2<1> ,
         \PDE_ALUOp2<0> , \PDE_Immediate<15> , \PDE_Immediate<14> ,
         \PDE_Immediate<13> , \PDE_Immediate<12> , \PDE_Immediate<11> ,
         \PDE_Immediate<10> , \PDE_Immediate<9> , \PDE_Immediate<8> ,
         \PDE_Immediate<7> , \PDE_Immediate<6> , \PDE_Immediate<5> ,
         \PDE_Immediate<4> , \PDE_Immediate<3> , \PDE_Immediate<2> ,
         \PDE_Immediate<1> , \PDE_Immediate<0> , \PDE_ALUOpcode<2> ,
         \PDE_ALUOpcode<1> , \PDE_ALUOpcode<0> , \PDE_Func<1> , \PDE_Func<0> ,
         PDE_ALUSrc, PDE_Branch, PDE_Jump, PDE_JumpReg, PDE_Set, PDE_Btr,
         PDE_MemWrite, PDE_MemRead, PDE_MemToReg, PDE_Halt, PDE_InvA, PDE_InvB,
         PDE_Cin, _19_net_, \PDE_Rs<2> , \PDE_Rs<1> , \PDE_Rs<0> , \PDE_Rt<2> ,
         \PDE_Rt<1> , \PDE_Rt<0> , \PDE_Rd<2> , \PDE_Rd<1> , \PDE_Rd<0> ,
         _20_net_, \PDE_DecodeIncPC<15> , \PDE_DecodeIncPC<14> ,
         \PDE_DecodeIncPC<13> , \PDE_DecodeIncPC<12> , \PDE_DecodeIncPC<11> ,
         \PDE_DecodeIncPC<10> , \PDE_DecodeIncPC<9> , \PDE_DecodeIncPC<8> ,
         \PDE_DecodeIncPC<7> , \PDE_DecodeIncPC<6> , \PDE_DecodeIncPC<5> ,
         \PDE_DecodeIncPC<4> , \PDE_DecodeIncPC<3> , \PDE_DecodeIncPC<2> ,
         \PDE_DecodeIncPC<1> , \PDE_DecodeIncPC<0> , PDE_Link,
         \E_ExecuteResult<15> , \E_ExecuteResult<14> , \E_ExecuteResult<13> ,
         \E_ExecuteResult<12> , \E_ExecuteResult<11> , \E_ExecuteResult<10> ,
         \E_ExecuteResult<9> , \E_ExecuteResult<8> , \E_ExecuteResult<7> ,
         \E_ExecuteResult<6> , \E_ExecuteResult<5> , \E_ExecuteResult<4> ,
         \E_ExecuteResult<3> , \E_ExecuteResult<2> , \E_ExecuteResult<1> ,
         \E_ExecuteResult<0> , \PEM_Address<15> , \PEM_Address<14> ,
         \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> ,
         \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> ,
         \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> ,
         \PEM_Address<4> , \PEM_Address<3> , \PEM_Address<2> ,
         \PEM_Address<1> , \PEM_Address<0> , \PMW_ExecuteOut<15> ,
         \PMW_ExecuteOut<14> , \PMW_ExecuteOut<13> , \PMW_ExecuteOut<12> ,
         \PMW_ExecuteOut<11> , \PMW_ExecuteOut<10> , \PMW_ExecuteOut<9> ,
         \PMW_ExecuteOut<8> , \PMW_ExecuteOut<7> , \PMW_ExecuteOut<6> ,
         \PMW_ExecuteOut<5> , \PMW_ExecuteOut<4> , \PMW_ExecuteOut<3> ,
         \PMW_ExecuteOut<2> , \PMW_ExecuteOut<1> , \PMW_ExecuteOut<0> ,
         PEM_MemRead, PEM_MemWrite, PEM_MemToReg, \PEM_WriteData<15> ,
         \PEM_WriteData<14> , \PEM_WriteData<13> , \PEM_WriteData<12> ,
         \PEM_WriteData<11> , \PEM_WriteData<10> , \PEM_WriteData<9> ,
         \PEM_WriteData<8> , \PEM_WriteData<7> , \PEM_WriteData<6> ,
         \PEM_WriteData<5> , \PEM_WriteData<4> , \PEM_WriteData<3> ,
         \PEM_WriteData<2> , \PEM_WriteData<1> , \PEM_WriteData<0> ,
         \PEM_Rs<2> , \PEM_Rs<1> , \PEM_Rs<0> , \PEM_Rt<2> , \PEM_Rt<1> ,
         \PEM_Rt<0> , \PEM_Rd<2> , \PEM_Rd<1> , \PEM_Rd<0> , \M_ReadData<15> ,
         \M_ReadData<14> , \M_ReadData<13> , \M_ReadData<12> ,
         \M_ReadData<11> , \M_ReadData<10> , \M_ReadData<9> , \M_ReadData<8> ,
         \M_ReadData<7> , \M_ReadData<6> , \M_ReadData<5> , \M_ReadData<4> ,
         \M_ReadData<3> , \M_ReadData<2> , \M_ReadData<1> , \M_ReadData<0> ,
         \PMW_MemOut<15> , \PMW_MemOut<14> , \PMW_MemOut<13> ,
         \PMW_MemOut<12> , \PMW_MemOut<11> , \PMW_MemOut<10> , \PMW_MemOut<9> ,
         \PMW_MemOut<8> , \PMW_MemOut<7> , \PMW_MemOut<6> , \PMW_MemOut<5> ,
         \PMW_MemOut<4> , \PMW_MemOut<3> , \PMW_MemOut<2> , \PMW_MemOut<1> ,
         \PMW_MemOut<0> , PMW_MemToReg, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30,
         n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  OR2X2 U7 ( .A(n62), .B(_2_net_), .Y(_3_net_) );
  AND2X2 U9 ( .A(D_RtValid), .B(n7), .Y(_19_net_) );
  OR2X2 U19 ( .A(n46), .B(n65), .Y(_2_net_) );
  NOR3X1 U26 ( .A(n62), .B(n65), .C(n68), .Y(_15_net_) );
  AOI22X1 U27 ( .A(PDE_RegFileWrEn), .B(n43), .C(PEM_RegFileWrEn), .D(n44), 
        .Y(n8) );
  NAND3X1 U28 ( .A(n48), .B(n51), .C(n53), .Y(n10) );
  NAND3X1 U29 ( .A(n14), .B(n15), .C(n61), .Y(n13) );
  XOR2X1 U31 ( .A(\PEM_WriteReg<2> ), .B(\D_Rs<2> ), .Y(n17) );
  XNOR2X1 U32 ( .A(\D_Rs<1> ), .B(\PEM_WriteReg<1> ), .Y(n15) );
  XNOR2X1 U33 ( .A(\D_Rs<0> ), .B(\PEM_WriteReg<0> ), .Y(n14) );
  NAND3X1 U34 ( .A(n18), .B(n19), .C(n20), .Y(n12) );
  NOR3X1 U35 ( .A(n21), .B(n69), .C(n71), .Y(n20) );
  XOR2X1 U36 ( .A(\PEM_WriteReg<2> ), .B(\D_Rd<2> ), .Y(n21) );
  XNOR2X1 U37 ( .A(\D_Rd<1> ), .B(\PEM_WriteReg<1> ), .Y(n19) );
  XNOR2X1 U38 ( .A(\D_Rd<0> ), .B(\PEM_WriteReg<0> ), .Y(n18) );
  NAND3X1 U39 ( .A(n22), .B(n23), .C(n59), .Y(n11) );
  XOR2X1 U41 ( .A(\PEM_WriteReg<2> ), .B(\D_Rt<2> ), .Y(n25) );
  XNOR2X1 U42 ( .A(\D_Rt<1> ), .B(\PEM_WriteReg<1> ), .Y(n23) );
  XNOR2X1 U43 ( .A(\D_Rt<0> ), .B(\PEM_WriteReg<0> ), .Y(n22) );
  NAND3X1 U44 ( .A(n42), .B(n50), .C(n47), .Y(n9) );
  NAND3X1 U45 ( .A(n29), .B(n30), .C(n57), .Y(n28) );
  XOR2X1 U47 ( .A(\PDE_WriteReg<2> ), .B(\D_Rs<2> ), .Y(n32) );
  XNOR2X1 U48 ( .A(\D_Rs<1> ), .B(\PDE_WriteReg<1> ), .Y(n30) );
  XNOR2X1 U49 ( .A(\D_Rs<0> ), .B(\PDE_WriteReg<0> ), .Y(n29) );
  NAND3X1 U50 ( .A(n33), .B(n34), .C(n35), .Y(n27) );
  NOR3X1 U51 ( .A(n36), .B(n69), .C(n71), .Y(n35) );
  XOR2X1 U52 ( .A(\PDE_WriteReg<2> ), .B(\D_Rd<2> ), .Y(n36) );
  XNOR2X1 U53 ( .A(\D_Rd<1> ), .B(\PDE_WriteReg<1> ), .Y(n34) );
  XNOR2X1 U54 ( .A(\D_Rd<0> ), .B(\PDE_WriteReg<0> ), .Y(n33) );
  NAND3X1 U55 ( .A(n37), .B(n38), .C(n55), .Y(n26) );
  XOR2X1 U57 ( .A(\PDE_WriteReg<2> ), .B(\D_Rt<2> ), .Y(n40) );
  XNOR2X1 U58 ( .A(\D_Rt<1> ), .B(\PDE_WriteReg<1> ), .Y(n38) );
  XNOR2X1 U59 ( .A(\D_Rt<0> ), .B(\PDE_WriteReg<0> ), .Y(n37) );
  fetch f ( .BranchPC({\E_BranchPC<15> , \E_BranchPC<14> , \E_BranchPC<13> , 
        \E_BranchPC<12> , \E_BranchPC<11> , \E_BranchPC<10> , \E_BranchPC<9> , 
        \E_BranchPC<8> , \E_BranchPC<7> , \E_BranchPC<6> , \E_BranchPC<5> , 
        \E_BranchPC<4> , \E_BranchPC<3> , \E_BranchPC<2> , \E_BranchPC<1> , 
        \E_BranchPC<0> }), .BranchJumpTaken(n46), .clk(clk), .rst(n65), .Halt(
        PEM_Halt), .Rti(D_Rti), .Exception(D_Exception), .Stall(n62), .Instr({
        \F_Instr<15> , \F_Instr<14> , \F_Instr<13> , \F_Instr<12> , 
        \F_Instr<11> , \F_Instr<10> , \F_Instr<9> , \F_Instr<8> , \F_Instr<7> , 
        \F_Instr<6> , \F_Instr<5> , \F_Instr<4> , \F_Instr<3> , \F_Instr<2> , 
        \F_Instr<1> , \F_Instr<0> }), .IncPC({\F_IncPC<15> , \F_IncPC<14> , 
        \F_IncPC<13> , \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , 
        \F_IncPC<9> , \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , 
        \F_IncPC<4> , \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> })
         );
  pipe_fd fd ( .Stall(n62), .Flush(_2_net_), .rst(_2_net_), .clk(clk), .Instr(
        {\F_Instr<15> , \F_Instr<14> , \F_Instr<13> , \F_Instr<12> , 
        \F_Instr<11> , \F_Instr<10> , \F_Instr<9> , \F_Instr<8> , \F_Instr<7> , 
        \F_Instr<6> , \F_Instr<5> , \F_Instr<4> , \F_Instr<3> , \F_Instr<2> , 
        \F_Instr<1> , \F_Instr<0> }), .IncPC({\F_IncPC<15> , \F_IncPC<14> , 
        \F_IncPC<13> , \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , 
        \F_IncPC<9> , \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , 
        \F_IncPC<4> , \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> }), 
        .Instr_Out({\PFD_Instr<15> , \PFD_Instr<14> , \PFD_Instr<13> , 
        \PFD_Instr<12> , \PFD_Instr<11> , \PFD_Instr<10> , \PFD_Instr<9> , 
        \PFD_Instr<8> , \PFD_Instr<7> , \PFD_Instr<6> , \PFD_Instr<5> , 
        \PFD_Instr<4> , \PFD_Instr<3> , \PFD_Instr<2> , \PFD_Instr<1> , 
        \PFD_Instr<0> }), .IncPC_Out({\PFD_IncPC<15> , \PFD_IncPC<14> , 
        \PFD_IncPC<13> , \PFD_IncPC<12> , \PFD_IncPC<11> , \PFD_IncPC<10> , 
        \PFD_IncPC<9> , \PFD_IncPC<8> , \PFD_IncPC<7> , \PFD_IncPC<6> , 
        \PFD_IncPC<5> , \PFD_IncPC<4> , \PFD_IncPC<3> , \PFD_IncPC<2> , 
        \PFD_IncPC<1> , \PFD_IncPC<0> }), .CPUActive(PFD_CPUActive) );
  decode d ( .clk(clk), .rst(n65), .Stall(n62), .Instr({\PFD_Instr<15> , 
        \PFD_Instr<14> , \PFD_Instr<13> , \PFD_Instr<12> , \PFD_Instr<11> , 
        \PFD_Instr<10> , \PFD_Instr<9> , \PFD_Instr<8> , \PFD_Instr<7> , 
        \PFD_Instr<6> , \PFD_Instr<5> , \PFD_Instr<4> , \PFD_Instr<3> , 
        \PFD_Instr<2> , \PFD_Instr<1> , \PFD_Instr<0> }), .WriteData({
        \W_WriteData<15> , \W_WriteData<14> , \W_WriteData<13> , 
        \W_WriteData<12> , \W_WriteData<11> , \W_WriteData<10> , 
        \W_WriteData<9> , \W_WriteData<8> , \W_WriteData<7> , \W_WriteData<6> , 
        \W_WriteData<5> , \W_WriteData<4> , \W_WriteData<3> , \W_WriteData<2> , 
        \W_WriteData<1> , \W_WriteData<0> }), .IncPC({\PFD_IncPC<15> , 
        \PFD_IncPC<14> , \PFD_IncPC<13> , \PFD_IncPC<12> , \PFD_IncPC<11> , 
        \PFD_IncPC<10> , \PFD_IncPC<9> , \PFD_IncPC<8> , \PFD_IncPC<7> , 
        \PFD_IncPC<6> , \PFD_IncPC<5> , \PFD_IncPC<4> , \PFD_IncPC<3> , 
        \PFD_IncPC<2> , \PFD_IncPC<1> , \PFD_IncPC<0> }), .ALUOp1({
        \D_ALUOp1<15> , \D_ALUOp1<14> , \D_ALUOp1<13> , \D_ALUOp1<12> , 
        \D_ALUOp1<11> , \D_ALUOp1<10> , \D_ALUOp1<9> , \D_ALUOp1<8> , 
        \D_ALUOp1<7> , \D_ALUOp1<6> , \D_ALUOp1<5> , \D_ALUOp1<4> , 
        \D_ALUOp1<3> , \D_ALUOp1<2> , \D_ALUOp1<1> , \D_ALUOp1<0> }), .ALUOp2(
        {\D_ALUOp2<15> , \D_ALUOp2<14> , \D_ALUOp2<13> , \D_ALUOp2<12> , 
        \D_ALUOp2<11> , \D_ALUOp2<10> , \D_ALUOp2<9> , \D_ALUOp2<8> , 
        \D_ALUOp2<7> , \D_ALUOp2<6> , \D_ALUOp2<5> , \D_ALUOp2<4> , 
        \D_ALUOp2<3> , \D_ALUOp2<2> , \D_ALUOp2<1> , \D_ALUOp2<0> }), .ALUSrc(
        D_ALUSrc), .Immediate({\D_Immediate<15> , \D_Immediate<14> , 
        \D_Immediate<13> , \D_Immediate<12> , \D_Immediate<11> , 
        \D_Immediate<10> , \D_Immediate<9> , \D_Immediate<8> , 
        \D_Immediate<7> , \D_Immediate<6> , \D_Immediate<5> , \D_Immediate<4> , 
        \D_Immediate<3> , \D_Immediate<2> , \D_Immediate<1> , \D_Immediate<0> }), .Branch(D_Branch), .Jump(D_Jump), .JumpReg(D_JumpReg), .Set(D_Set), .Btr(
        D_Btr), .InvA(D_InvA), .InvB(D_InvB), .Cin(D_Cin), .ALUOpcode({
        \D_ALUOpcode<2> , \D_ALUOpcode<1> , \D_ALUOpcode<0> }), .Func({
        \D_Func<1> , \D_Func<0> }), .MemWrite(D_MemWrite), .MemRead(D_MemRead), 
        .MemToReg(D_MemToReg), .Halt(D_Halt), .Exception(D_Exception), .Err(), 
        .Rti(D_Rti), .Rs({\D_Rs<2> , \D_Rs<1> , \D_Rs<0> }), .Rt({\D_Rt<2> , 
        \D_Rt<1> , \D_Rt<0> }), .Rd({\D_Rd<2> , \D_Rd<1> , \D_Rd<0> }), 
        .RegFileWrEn(PMW_RegFileWrEn), .RegFileWrEn_Out(D_RegFileWrEn), 
        .WriteReg({\PMW_WriteReg<2> , \PMW_WriteReg<1> , \PMW_WriteReg<0> }), 
        .WriteReg_Out({\D_WriteReg<2> , \D_WriteReg<1> , \D_WriteReg<0> }), 
        .RtValid(D_RtValid), .RsValid(D_RsValid), .RdValid(D_RdValid), .Link(
        D_Link), .Store(D_Store) );
  pipe_de pde ( .clk(clk), .rst(_3_net_), .Stall(1'b0), .Flush(_2_net_), 
        .ALUOp1({\D_ALUOp1<15> , \D_ALUOp1<14> , \D_ALUOp1<13> , 
        \D_ALUOp1<12> , \D_ALUOp1<11> , \D_ALUOp1<10> , \D_ALUOp1<9> , 
        \D_ALUOp1<8> , \D_ALUOp1<7> , \D_ALUOp1<6> , \D_ALUOp1<5> , 
        \D_ALUOp1<4> , \D_ALUOp1<3> , \D_ALUOp1<2> , \D_ALUOp1<1> , 
        \D_ALUOp1<0> }), .ALUOp2({\D_ALUOp2<15> , \D_ALUOp2<14> , 
        \D_ALUOp2<13> , \D_ALUOp2<12> , \D_ALUOp2<11> , \D_ALUOp2<10> , 
        \D_ALUOp2<9> , \D_ALUOp2<8> , \D_ALUOp2<7> , \D_ALUOp2<6> , 
        \D_ALUOp2<5> , \D_ALUOp2<4> , \D_ALUOp2<3> , \D_ALUOp2<2> , 
        \D_ALUOp2<1> , \D_ALUOp2<0> }), .Immediate({\D_Immediate<15> , 
        \D_Immediate<14> , \D_Immediate<13> , \D_Immediate<12> , 
        \D_Immediate<11> , \D_Immediate<10> , \D_Immediate<9> , 
        \D_Immediate<8> , \D_Immediate<7> , \D_Immediate<6> , \D_Immediate<5> , 
        \D_Immediate<4> , \D_Immediate<3> , \D_Immediate<2> , \D_Immediate<1> , 
        \D_Immediate<0> }), .ALUOpcode({\D_ALUOpcode<2> , \D_ALUOpcode<1> , 
        \D_ALUOpcode<0> }), .Func({\D_Func<1> , \_5_net_<0> }), .ALUSrc(
        _6_net_), .Branch(_7_net_), .Jump(_8_net_), .JumpReg(_9_net_), .Set(
        _10_net_), .Btr(_11_net_), .MemWrite(_12_net_), .MemRead(_14_net_), 
        .MemToReg(_14_net_), .Halt(_15_net_), .InvA(_16_net_), .InvB(_17_net_), 
        .Cin(_18_net_), .IncPC({\F_IncPC<15> , \F_IncPC<14> , \F_IncPC<13> , 
        \F_IncPC<12> , \F_IncPC<11> , \F_IncPC<10> , \F_IncPC<9> , 
        \F_IncPC<8> , \F_IncPC<7> , \F_IncPC<6> , \F_IncPC<5> , \F_IncPC<4> , 
        \F_IncPC<3> , \F_IncPC<2> , \F_IncPC<1> , \F_IncPC<0> }), .CPUActive(
        PFD_CPUActive), .ALUOp1_Out({\PDE_ALUOp1<15> , \PDE_ALUOp1<14> , 
        \PDE_ALUOp1<13> , \PDE_ALUOp1<12> , \PDE_ALUOp1<11> , \PDE_ALUOp1<10> , 
        \PDE_ALUOp1<9> , \PDE_ALUOp1<8> , \PDE_ALUOp1<7> , \PDE_ALUOp1<6> , 
        \PDE_ALUOp1<5> , \PDE_ALUOp1<4> , \PDE_ALUOp1<3> , \PDE_ALUOp1<2> , 
        \PDE_ALUOp1<1> , \PDE_ALUOp1<0> }), .ALUOp2_Out({\PDE_ALUOp2<15> , 
        \PDE_ALUOp2<14> , \PDE_ALUOp2<13> , \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , 
        \PDE_ALUOp2<10> , \PDE_ALUOp2<9> , \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , 
        \PDE_ALUOp2<6> , \PDE_ALUOp2<5> , \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , 
        \PDE_ALUOp2<2> , \PDE_ALUOp2<1> , \PDE_ALUOp2<0> }), .Immediate_Out({
        \PDE_Immediate<15> , \PDE_Immediate<14> , \PDE_Immediate<13> , 
        \PDE_Immediate<12> , \PDE_Immediate<11> , \PDE_Immediate<10> , 
        \PDE_Immediate<9> , \PDE_Immediate<8> , \PDE_Immediate<7> , 
        \PDE_Immediate<6> , \PDE_Immediate<5> , \PDE_Immediate<4> , 
        \PDE_Immediate<3> , \PDE_Immediate<2> , \PDE_Immediate<1> , 
        \PDE_Immediate<0> }), .ALUOpcode_Out({\PDE_ALUOpcode<2> , 
        \PDE_ALUOpcode<1> , \PDE_ALUOpcode<0> }), .Func_Out({\PDE_Func<1> , 
        \PDE_Func<0> }), .ALUSrc_Out(PDE_ALUSrc), .Branch_Out(PDE_Branch), 
        .Jump_Out(PDE_Jump), .JumpReg_Out(PDE_JumpReg), .Set_Out(PDE_Set), 
        .Btr_Out(PDE_Btr), .MemWrite_Out(PDE_MemWrite), .MemRead_Out(
        PDE_MemRead), .MemToReg_Out(PDE_MemToReg), .Halt_Out(PDE_Halt), 
        .InvA_Out(PDE_InvA), .InvB_Out(PDE_InvB), .Cin_Out(PDE_Cin), .Rs({
        \D_Rs<2> , \D_Rs<1> , \D_Rs<0> }), .Rt({\D_Rt<2> , \D_Rt<1> , 
        \D_Rt<0> }), .Rd({\D_Rd<2> , \D_Rd<1> , \D_Rd<0> }), .Rs_Out({
        \PDE_Rs<2> , \PDE_Rs<1> , \PDE_Rs<0> }), .Rt_Out({\PDE_Rt<2> , 
        \PDE_Rt<1> , \PDE_Rt<0> }), .Rd_Out({\PDE_Rd<2> , \PDE_Rd<1> , 
        \PDE_Rd<0> }), .RegFileWrEn(_20_net_), .RegFileWrEn_Out(
        PDE_RegFileWrEn), .IncPC_Out({\PDE_IncPC<15> , \PDE_IncPC<14> , 
        \PDE_IncPC<13> , \PDE_IncPC<12> , \PDE_IncPC<11> , \PDE_IncPC<10> , 
        \PDE_IncPC<9> , \PDE_IncPC<8> , \PDE_IncPC<7> , \PDE_IncPC<6> , 
        \PDE_IncPC<5> , \PDE_IncPC<4> , \PDE_IncPC<3> , \PDE_IncPC<2> , 
        \PDE_IncPC<1> , \PDE_IncPC<0> }), .WriteReg({\D_WriteReg<2> , 
        \D_WriteReg<1> , \D_WriteReg<0> }), .WriteReg_Out({\PDE_WriteReg<2> , 
        \PDE_WriteReg<1> , \PDE_WriteReg<0> }), .RtValid(_19_net_), 
        .RtValid_Out(), .CPUActive_Out(), .RsValid(D_RsValid), .RdValid(
        D_RdValid), .RsValid_Out(), .RdValid_Out(), .DecodeIncPC({
        \PFD_IncPC<15> , \PFD_IncPC<14> , \PFD_IncPC<13> , \PFD_IncPC<12> , 
        \PFD_IncPC<11> , \PFD_IncPC<10> , \PFD_IncPC<9> , \PFD_IncPC<8> , 
        \PFD_IncPC<7> , \PFD_IncPC<6> , \PFD_IncPC<5> , \PFD_IncPC<4> , 
        \PFD_IncPC<3> , \PFD_IncPC<2> , \PFD_IncPC<1> , \PFD_IncPC<0> }), 
        .DecodeIncPC_Out({\PDE_DecodeIncPC<15> , \PDE_DecodeIncPC<14> , 
        \PDE_DecodeIncPC<13> , \PDE_DecodeIncPC<12> , \PDE_DecodeIncPC<11> , 
        \PDE_DecodeIncPC<10> , \PDE_DecodeIncPC<9> , \PDE_DecodeIncPC<8> , 
        \PDE_DecodeIncPC<7> , \PDE_DecodeIncPC<6> , \PDE_DecodeIncPC<5> , 
        \PDE_DecodeIncPC<4> , \PDE_DecodeIncPC<3> , \PDE_DecodeIncPC<2> , 
        \PDE_DecodeIncPC<1> , \PDE_DecodeIncPC<0> }), .Link(D_Link), 
        .Link_Out(PDE_Link) );
  execute e ( .ALUOp1({\PDE_ALUOp1<15> , \PDE_ALUOp1<14> , \PDE_ALUOp1<13> , 
        \PDE_ALUOp1<12> , \PDE_ALUOp1<11> , \PDE_ALUOp1<10> , \PDE_ALUOp1<9> , 
        \PDE_ALUOp1<8> , \PDE_ALUOp1<7> , \PDE_ALUOp1<6> , \PDE_ALUOp1<5> , 
        \PDE_ALUOp1<4> , \PDE_ALUOp1<3> , \PDE_ALUOp1<2> , \PDE_ALUOp1<1> , 
        \PDE_ALUOp1<0> }), .ALUOp2({\PDE_ALUOp2<15> , \PDE_ALUOp2<14> , 
        \PDE_ALUOp2<13> , \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , \PDE_ALUOp2<10> , 
        \PDE_ALUOp2<9> , \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , \PDE_ALUOp2<6> , 
        \PDE_ALUOp2<5> , \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , \PDE_ALUOp2<2> , 
        \PDE_ALUOp2<1> , \PDE_ALUOp2<0> }), .Opcode({\PDE_ALUOpcode<2> , 
        \PDE_ALUOpcode<1> , \PDE_ALUOpcode<0> }), .IncPC({\PDE_IncPC<15> , 
        \PDE_IncPC<14> , \PDE_IncPC<13> , \PDE_IncPC<12> , \PDE_IncPC<11> , 
        \PDE_IncPC<10> , \PDE_IncPC<9> , \PDE_IncPC<8> , \PDE_IncPC<7> , 
        \PDE_IncPC<6> , \PDE_IncPC<5> , \PDE_IncPC<4> , \PDE_IncPC<3> , 
        \PDE_IncPC<2> , \PDE_IncPC<1> , \PDE_IncPC<0> }), .Jump(PDE_Jump), 
        .Branch(PDE_Branch), .JumpReg(PDE_JumpReg), .Set(PDE_Set), .InvA(
        PDE_InvA), .InvB(PDE_InvB), .Cin(PDE_Cin), .Btr(PDE_Btr), .Func({
        \PDE_Func<1> , \PDE_Func<0> }), .Imm({\PDE_Immediate<15> , 
        \PDE_Immediate<14> , \PDE_Immediate<13> , \PDE_Immediate<12> , 
        \PDE_Immediate<11> , \PDE_Immediate<10> , \PDE_Immediate<9> , 
        \PDE_Immediate<8> , \PDE_Immediate<7> , \PDE_Immediate<6> , 
        \PDE_Immediate<5> , \PDE_Immediate<4> , \PDE_Immediate<3> , 
        \PDE_Immediate<2> , \PDE_Immediate<1> , \PDE_Immediate<0> }), .ALUSrc(
        PDE_ALUSrc), .Result({\E_ExecuteResult<15> , \E_ExecuteResult<14> , 
        \E_ExecuteResult<13> , \E_ExecuteResult<12> , \E_ExecuteResult<11> , 
        \E_ExecuteResult<10> , \E_ExecuteResult<9> , \E_ExecuteResult<8> , 
        \E_ExecuteResult<7> , \E_ExecuteResult<6> , \E_ExecuteResult<5> , 
        \E_ExecuteResult<4> , \E_ExecuteResult<3> , \E_ExecuteResult<2> , 
        \E_ExecuteResult<1> , \E_ExecuteResult<0> }), .NextPC({
        \E_BranchPC<15> , \E_BranchPC<14> , \E_BranchPC<13> , \E_BranchPC<12> , 
        \E_BranchPC<11> , \E_BranchPC<10> , \E_BranchPC<9> , \E_BranchPC<8> , 
        \E_BranchPC<7> , \E_BranchPC<6> , \E_BranchPC<5> , \E_BranchPC<4> , 
        \E_BranchPC<3> , \E_BranchPC<2> , \E_BranchPC<1> , \E_BranchPC<0> }), 
        .Err(), .BranchJumpTaken(E_BranchJumpTaken), .rst(n65), .DecodeIncPC({
        \PDE_DecodeIncPC<15> , \PDE_DecodeIncPC<14> , \PDE_DecodeIncPC<13> , 
        \PDE_DecodeIncPC<12> , \PDE_DecodeIncPC<11> , \PDE_DecodeIncPC<10> , 
        \PDE_DecodeIncPC<9> , \PDE_DecodeIncPC<8> , \PDE_DecodeIncPC<7> , 
        \PDE_DecodeIncPC<6> , \PDE_DecodeIncPC<5> , \PDE_DecodeIncPC<4> , 
        \PDE_DecodeIncPC<3> , \PDE_DecodeIncPC<2> , \PDE_DecodeIncPC<1> , 
        \PDE_DecodeIncPC<0> }), .Link(PDE_Link), .ForwardALUOp1({1'b0, 1'b0}), 
        .ForwardALUOp2({1'b0, 1'b0}), .PipeMW_Result({\PMW_ExecuteOut<15> , 
        \PMW_ExecuteOut<14> , \PMW_ExecuteOut<13> , \PMW_ExecuteOut<12> , 
        \PMW_ExecuteOut<11> , \PMW_ExecuteOut<10> , \PMW_ExecuteOut<9> , 
        \PMW_ExecuteOut<8> , \PMW_ExecuteOut<7> , \PMW_ExecuteOut<6> , 
        \PMW_ExecuteOut<5> , \PMW_ExecuteOut<4> , \PMW_ExecuteOut<3> , 
        \PMW_ExecuteOut<2> , \PMW_ExecuteOut<1> , \PMW_ExecuteOut<0> }), 
        .PipeEM_Result({\PEM_Address<15> , \PEM_Address<14> , 
        \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> , 
        \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> , 
        \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> , n63, 
        \PEM_Address<3> , \PEM_Address<2> , \PEM_Address<1> , \PEM_Address<0> }) );
  pipe_em pem ( .Stall(1'b0), .rst(n65), .clk(clk), .Result({
        \E_ExecuteResult<15> , \E_ExecuteResult<14> , \E_ExecuteResult<13> , 
        \E_ExecuteResult<12> , \E_ExecuteResult<11> , \E_ExecuteResult<10> , 
        \E_ExecuteResult<9> , \E_ExecuteResult<8> , \E_ExecuteResult<7> , 
        \E_ExecuteResult<6> , \E_ExecuteResult<5> , \E_ExecuteResult<4> , 
        \E_ExecuteResult<3> , \E_ExecuteResult<2> , \E_ExecuteResult<1> , 
        \E_ExecuteResult<0> }), .MemRead(PDE_MemRead), .MemWrite(PDE_MemWrite), 
        .MemToReg(PDE_MemToReg), .Halt(PDE_Halt), .ALUOp2({\PDE_ALUOp2<15> , 
        \PDE_ALUOp2<14> , \PDE_ALUOp2<13> , \PDE_ALUOp2<12> , \PDE_ALUOp2<11> , 
        \PDE_ALUOp2<10> , \PDE_ALUOp2<9> , \PDE_ALUOp2<8> , \PDE_ALUOp2<7> , 
        \PDE_ALUOp2<6> , \PDE_ALUOp2<5> , \PDE_ALUOp2<4> , \PDE_ALUOp2<3> , 
        \PDE_ALUOp2<2> , \PDE_ALUOp2<1> , \PDE_ALUOp2<0> }), .RegFileWrEn(
        PDE_RegFileWrEn), .Rs({\PDE_Rs<2> , \PDE_Rs<1> , \PDE_Rs<0> }), .Rt({
        \PDE_Rt<2> , \PDE_Rt<1> , \PDE_Rt<0> }), .Rd({\PDE_Rd<2> , \PDE_Rd<1> , 
        \PDE_Rd<0> }), .WriteReg({\PDE_WriteReg<2> , \PDE_WriteReg<1> , 
        \PDE_WriteReg<0> }), .Address({\PEM_Address<15> , \PEM_Address<14> , 
        \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> , 
        \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> , 
        \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> , \PEM_Address<4> , 
        \PEM_Address<3> , \PEM_Address<2> , \PEM_Address<1> , \PEM_Address<0> }), .MemRead_Out(PEM_MemRead), .MemWrite_Out(PEM_MemWrite), .MemToReg_Out(
        PEM_MemToReg), .Halt_Out(PEM_Halt), .WriteData({\PEM_WriteData<15> , 
        \PEM_WriteData<14> , \PEM_WriteData<13> , \PEM_WriteData<12> , 
        \PEM_WriteData<11> , \PEM_WriteData<10> , \PEM_WriteData<9> , 
        \PEM_WriteData<8> , \PEM_WriteData<7> , \PEM_WriteData<6> , 
        \PEM_WriteData<5> , \PEM_WriteData<4> , \PEM_WriteData<3> , 
        \PEM_WriteData<2> , \PEM_WriteData<1> , \PEM_WriteData<0> }), 
        .RegFileWrEn_Out(PEM_RegFileWrEn), .Rs_Out({\PEM_Rs<2> , \PEM_Rs<1> , 
        \PEM_Rs<0> }), .Rt_Out({\PEM_Rt<2> , \PEM_Rt<1> , \PEM_Rt<0> }), 
        .Rd_Out({\PEM_Rd<2> , \PEM_Rd<1> , \PEM_Rd<0> }), .WriteReg_Out({
        \PEM_WriteReg<2> , \PEM_WriteReg<1> , \PEM_WriteReg<0> }) );
  memory m ( .MemRead(PEM_MemRead), .MemWrite(PEM_MemWrite), .halt(PEM_Halt), 
        .clk(clk), .rst(n65), .Address({\PEM_Address<15> , \PEM_Address<14> , 
        \PEM_Address<13> , \PEM_Address<12> , \PEM_Address<11> , 
        \PEM_Address<10> , \PEM_Address<9> , \PEM_Address<8> , 
        \PEM_Address<7> , \PEM_Address<6> , \PEM_Address<5> , n63, 
        \PEM_Address<3> , \PEM_Address<2> , \PEM_Address<1> , \PEM_Address<0> }), .WriteData({\PEM_WriteData<15> , \PEM_WriteData<14> , \PEM_WriteData<13> , 
        \PEM_WriteData<12> , \PEM_WriteData<11> , \PEM_WriteData<10> , 
        \PEM_WriteData<9> , \PEM_WriteData<8> , \PEM_WriteData<7> , 
        \PEM_WriteData<6> , \PEM_WriteData<5> , \PEM_WriteData<4> , 
        \PEM_WriteData<3> , \PEM_WriteData<2> , \PEM_WriteData<1> , 
        \PEM_WriteData<0> }), .ReadData({\M_ReadData<15> , \M_ReadData<14> , 
        \M_ReadData<13> , \M_ReadData<12> , \M_ReadData<11> , \M_ReadData<10> , 
        \M_ReadData<9> , \M_ReadData<8> , \M_ReadData<7> , \M_ReadData<6> , 
        \M_ReadData<5> , \M_ReadData<4> , \M_ReadData<3> , \M_ReadData<2> , 
        \M_ReadData<1> , \M_ReadData<0> }) );
  pipe_mw pmw ( .Stall(1'b0), .rst(n65), .clk(clk), .ExecuteOut({
        \PEM_Address<15> , \PEM_Address<14> , \PEM_Address<13> , 
        \PEM_Address<12> , \PEM_Address<11> , \PEM_Address<10> , 
        \PEM_Address<9> , \PEM_Address<8> , \PEM_Address<7> , \PEM_Address<6> , 
        \PEM_Address<5> , n63, \PEM_Address<3> , \PEM_Address<2> , 
        \PEM_Address<1> , \PEM_Address<0> }), .MemOut({\M_ReadData<15> , 
        \M_ReadData<14> , \M_ReadData<13> , \M_ReadData<12> , \M_ReadData<11> , 
        \M_ReadData<10> , \M_ReadData<9> , \M_ReadData<8> , \M_ReadData<7> , 
        \M_ReadData<6> , \M_ReadData<5> , \M_ReadData<4> , \M_ReadData<3> , 
        \M_ReadData<2> , \M_ReadData<1> , \M_ReadData<0> }), .MemToReg(
        PEM_MemToReg), .RegFileWrEn(PEM_RegFileWrEn), .Rs({\PEM_Rs<2> , 
        \PEM_Rs<1> , \PEM_Rs<0> }), .Rt({\PEM_Rt<2> , \PEM_Rt<1> , \PEM_Rt<0> }), .Rd({\PEM_Rd<2> , \PEM_Rd<1> , \PEM_Rd<0> }), .WriteReg({\PEM_WriteReg<2> , 
        \PEM_WriteReg<1> , \PEM_WriteReg<0> }), .ExecuteOut_Out({
        \PMW_ExecuteOut<15> , \PMW_ExecuteOut<14> , \PMW_ExecuteOut<13> , 
        \PMW_ExecuteOut<12> , \PMW_ExecuteOut<11> , \PMW_ExecuteOut<10> , 
        \PMW_ExecuteOut<9> , \PMW_ExecuteOut<8> , \PMW_ExecuteOut<7> , 
        \PMW_ExecuteOut<6> , \PMW_ExecuteOut<5> , \PMW_ExecuteOut<4> , 
        \PMW_ExecuteOut<3> , \PMW_ExecuteOut<2> , \PMW_ExecuteOut<1> , 
        \PMW_ExecuteOut<0> }), .MemOut_Out({\PMW_MemOut<15> , \PMW_MemOut<14> , 
        \PMW_MemOut<13> , \PMW_MemOut<12> , \PMW_MemOut<11> , \PMW_MemOut<10> , 
        \PMW_MemOut<9> , \PMW_MemOut<8> , \PMW_MemOut<7> , \PMW_MemOut<6> , 
        \PMW_MemOut<5> , \PMW_MemOut<4> , \PMW_MemOut<3> , \PMW_MemOut<2> , 
        \PMW_MemOut<1> , \PMW_MemOut<0> }), .MemToReg_Out(PMW_MemToReg), 
        .RegFileWrEn_Out(PMW_RegFileWrEn), .WriteReg_Out({\PMW_WriteReg<2> , 
        \PMW_WriteReg<1> , \PMW_WriteReg<0> }), .Rs_Out(), .Rt_Out(), 
        .Rd_Out() );
  writeback w ( .ExecuteOut({\PMW_ExecuteOut<15> , \PMW_ExecuteOut<14> , 
        \PMW_ExecuteOut<13> , \PMW_ExecuteOut<12> , \PMW_ExecuteOut<11> , 
        \PMW_ExecuteOut<10> , \PMW_ExecuteOut<9> , \PMW_ExecuteOut<8> , 
        \PMW_ExecuteOut<7> , \PMW_ExecuteOut<6> , \PMW_ExecuteOut<5> , 
        \PMW_ExecuteOut<4> , \PMW_ExecuteOut<3> , \PMW_ExecuteOut<2> , 
        \PMW_ExecuteOut<1> , \PMW_ExecuteOut<0> }), .MemOut({\PMW_MemOut<15> , 
        \PMW_MemOut<14> , \PMW_MemOut<13> , \PMW_MemOut<12> , \PMW_MemOut<11> , 
        \PMW_MemOut<10> , \PMW_MemOut<9> , \PMW_MemOut<8> , \PMW_MemOut<7> , 
        \PMW_MemOut<6> , \PMW_MemOut<5> , \PMW_MemOut<4> , \PMW_MemOut<3> , 
        \PMW_MemOut<2> , \PMW_MemOut<1> , \PMW_MemOut<0> }), .MemToReg(
        PMW_MemToReg), .WriteData({\W_WriteData<15> , \W_WriteData<14> , 
        \W_WriteData<13> , \W_WriteData<12> , \W_WriteData<11> , 
        \W_WriteData<10> , \W_WriteData<9> , \W_WriteData<8> , 
        \W_WriteData<7> , \W_WriteData<6> , \W_WriteData<5> , \W_WriteData<4> , 
        \W_WriteData<3> , \W_WriteData<2> , \W_WriteData<1> , \W_WriteData<0> }) );
  AND2X1 U60 ( .A(D_RegFileWrEn), .B(n7), .Y(_20_net_) );
  AND2X1 U61 ( .A(\D_Func<0> ), .B(n7), .Y(\_5_net_<0> ) );
  AND2X1 U62 ( .A(D_ALUSrc), .B(n7), .Y(_6_net_) );
  AND2X1 U63 ( .A(D_Branch), .B(n7), .Y(_7_net_) );
  AND2X1 U64 ( .A(D_Jump), .B(n7), .Y(_8_net_) );
  AND2X1 U65 ( .A(D_JumpReg), .B(n7), .Y(_9_net_) );
  AND2X1 U66 ( .A(D_Set), .B(n7), .Y(_10_net_) );
  AND2X1 U67 ( .A(D_Btr), .B(n7), .Y(_11_net_) );
  AND2X1 U68 ( .A(D_InvA), .B(n7), .Y(_16_net_) );
  AND2X1 U69 ( .A(D_InvB), .B(n7), .Y(_17_net_) );
  AND2X1 U70 ( .A(D_Cin), .B(n7), .Y(_18_net_) );
  INVX1 U71 ( .A(rst), .Y(n66) );
  INVX1 U72 ( .A(\PEM_Address<4> ), .Y(n64) );
  INVX1 U73 ( .A(D_RtValid), .Y(n70) );
  INVX1 U74 ( .A(D_RsValid), .Y(n67) );
  INVX1 U75 ( .A(D_Store), .Y(n71) );
  AND2X1 U76 ( .A(D_MemWrite), .B(n7), .Y(_12_net_) );
  AND2X1 U77 ( .A(D_MemToReg), .B(n7), .Y(_14_net_) );
  INVX1 U78 ( .A(D_Halt), .Y(n68) );
  INVX2 U79 ( .A(n66), .Y(n65) );
  OR2X2 U80 ( .A(n8), .B(_2_net_), .Y(n41) );
  BUFX2 U81 ( .A(n28), .Y(n42) );
  BUFX2 U82 ( .A(n9), .Y(n43) );
  BUFX2 U83 ( .A(n10), .Y(n44) );
  INVX2 U84 ( .A(n41), .Y(n62) );
  INVX1 U85 ( .A(E_BranchJumpTaken), .Y(n45) );
  INVX1 U86 ( .A(n45), .Y(n46) );
  BUFX2 U87 ( .A(n26), .Y(n47) );
  BUFX2 U88 ( .A(n11), .Y(n48) );
  INVX1 U89 ( .A(n27), .Y(n49) );
  INVX1 U90 ( .A(n49), .Y(n50) );
  BUFX2 U91 ( .A(n12), .Y(n51) );
  INVX1 U92 ( .A(n13), .Y(n52) );
  INVX1 U93 ( .A(n52), .Y(n53) );
  OR2X1 U94 ( .A(n70), .B(n40), .Y(n54) );
  INVX1 U95 ( .A(n54), .Y(n55) );
  OR2X1 U96 ( .A(n67), .B(n32), .Y(n56) );
  INVX1 U97 ( .A(n56), .Y(n57) );
  OR2X1 U98 ( .A(n70), .B(n25), .Y(n58) );
  INVX1 U99 ( .A(n58), .Y(n59) );
  OR2X1 U100 ( .A(n67), .B(n17), .Y(n60) );
  INVX1 U101 ( .A(n60), .Y(n61) );
  INVX1 U102 ( .A(n64), .Y(n63) );
  INVX1 U103 ( .A(n62), .Y(n7) );
  INVX2 U104 ( .A(D_RdValid), .Y(n69) );
endmodule

