
module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memc_Size16_7 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n214, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1162), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1161), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1160), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1159), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1158), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1157), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1156), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1155), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1154), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1153), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1152), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1151), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1150), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1149), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1148), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1147), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1146), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1145), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1144), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1143), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1142), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1141), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1140), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1139), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1138), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1137), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1136), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1135), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1134), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1133), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1132), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1131), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1130), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1129), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1128), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1127), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1126), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1125), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1124), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1123), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1122), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1121), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1120), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1119), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1118), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1117), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1116), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1115), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1114), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1113), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1112), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1111), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1110), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1109), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1108), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1107), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1106), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1105), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1104), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1103), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1102), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1101), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1100), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1099), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1098), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1097), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1096), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1095), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1094), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1093), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1092), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1091), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1090), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1089), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1088), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1087), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1085), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1083), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1082), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1081), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1080), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1079), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1078), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1077), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1076), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1075), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1074), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1073), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1072), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1071), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1070), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1069), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1068), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1067), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1066), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1065), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1064), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1063), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1062), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1061), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1060), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1059), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1058), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1057), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1056), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1055), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1054), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1053), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1052), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1051), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1050), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1049), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1048), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1047), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1046), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1045), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1044), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1043), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1042), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1041), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1040), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1039), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1038), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1037), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1036), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1035), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1034), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1033), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1032), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1031), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1030), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1029), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1028), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1027), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1026), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1025), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1024), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1023), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1022), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1021), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1020), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1019), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1018), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1017), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1016), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1015), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1014), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1013), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1012), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1011), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1010), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1009), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1008), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1007), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1006), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1005), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1004), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1003), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1002), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1001), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1000), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n999), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n998), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n997), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n996), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n995), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n994), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n993), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n992), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n991), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n990), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n989), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n988), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n987), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n986), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n985), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n984), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n983), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n982), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n981), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n980), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n979), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n978), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n977), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n976), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n975), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n974), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n973), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n972), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n971), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n970), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n969), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n968), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n967), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n966), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n965), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n964), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n963), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n962), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n961), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n960), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n959), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n958), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n957), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n956), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n955), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n954), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n953), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n952), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n951), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n950), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n949), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n948), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n947), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n946), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n945), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n944), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n943), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n942), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n941), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n940), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n939), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n938), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n937), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n936), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n935), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n934), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n933), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n932), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n931), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n930), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n929), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n928), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n927), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n926), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n925), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n924), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n923), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n922), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n921), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n920), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n919), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n918), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n917), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n916), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n915), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n914), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n913), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n912), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n911), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n910), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n909), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n908), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n907), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n906), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n905), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n904), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n903), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n902), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n901), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n900), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n899), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n898), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n897), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n896), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n895), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n894), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n893), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n892), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n891), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n890), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n889), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n888), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n887), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n886), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n885), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n884), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n883), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n882), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n881), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n880), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n879), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n878), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n877), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n876), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n875), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n874), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n873), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n872), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n871), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n870), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n869), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n868), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n867), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n866), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n865), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n864), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n863), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n862), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n861), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n860), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n859), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n858), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n857), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n856), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n855), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n854), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n853), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n852), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n851), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n850), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n849), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n848), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n847), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n846), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n845), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n844), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n843), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n842), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n841), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n840), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n839), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n838), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n837), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n836), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n835), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n834), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n833), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n832), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n831), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n830), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n829), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n828), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n827), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n826), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n825), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n824), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n823), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n822), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n821), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n820), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n819), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n818), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n817), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n816), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n815), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n814), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n813), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n812), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n811), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n810), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n809), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n808), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n807), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n806), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n805), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n804), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n803), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n802), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n801), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n800), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n799), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n798), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n797), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n796), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n795), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n794), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n793), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n792), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n791), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n790), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n789), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n788), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n787), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n786), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n785), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n784), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n783), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n782), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n781), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n780), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n779), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n778), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n777), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n776), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n775), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n774), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n773), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n772), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n771), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n770), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n769), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n768), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n767), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n766), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n765), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n764), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n763), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n762), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n761), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n760), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n759), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n758), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n757), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n756), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n755), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n754), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n753), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n752), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n751), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n750), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n749), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n748), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n747), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n746), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n745), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n744), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n743), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n742), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n741), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n740), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n739), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n738), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n737), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n736), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n735), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n734), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n733), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n732), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n731), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n730), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n729), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n728), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n727), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n726), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n725), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n724), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n723), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n722), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n721), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n720), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n719), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n718), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n717), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n716), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n715), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n714), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n713), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n712), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n711), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n710), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n709), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n708), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n707), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n706), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n705), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n704), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n703), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n702), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n701), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n700), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n699), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n698), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n697), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n696), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n695), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n694), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n693), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n692), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n691), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n690), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n689), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n688), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n687), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n686), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n685), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n684), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n683), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n682), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n681), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n680), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n679), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n678), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n677), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n676), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n675), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n674), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n673), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n672), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n671), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n670), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n669), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n668), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n667), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n666), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n665), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n664), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n663), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n662), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n661), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n660), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n659), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n658), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n657), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n656), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n655), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n654), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n653), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n652), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n651), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n214) );
  INVX1 U2 ( .A(n1204), .Y(n1214) );
  INVX1 U3 ( .A(n1203), .Y(n1215) );
  INVX1 U4 ( .A(n1323), .Y(n1186) );
  INVX1 U5 ( .A(n1323), .Y(n1184) );
  INVX1 U6 ( .A(n1164), .Y(N31) );
  INVX1 U7 ( .A(n1204), .Y(n1205) );
  INVX1 U8 ( .A(n1204), .Y(n1206) );
  INVX1 U9 ( .A(n1200), .Y(n1189) );
  INVX1 U10 ( .A(n1204), .Y(n1207) );
  INVX1 U11 ( .A(n1200), .Y(n1190) );
  INVX1 U12 ( .A(n1200), .Y(n1191) );
  INVX1 U13 ( .A(n1203), .Y(n1208) );
  INVX1 U14 ( .A(n1188), .Y(n1192) );
  INVX1 U15 ( .A(n1203), .Y(n1209) );
  INVX1 U16 ( .A(n1188), .Y(n1193) );
  INVX1 U17 ( .A(n1202), .Y(n1210) );
  INVX1 U18 ( .A(n1188), .Y(n1194) );
  INVX1 U19 ( .A(n1201), .Y(n1212) );
  INVX1 U20 ( .A(n1187), .Y(n1195) );
  INVX1 U21 ( .A(n1203), .Y(n1213) );
  INVX1 U22 ( .A(n1187), .Y(n1196) );
  INVX1 U23 ( .A(n1187), .Y(n1197) );
  INVX1 U24 ( .A(n1201), .Y(n1216) );
  INVX1 U25 ( .A(n1201), .Y(n1217) );
  INVX1 U26 ( .A(n1188), .Y(n1198) );
  INVX1 U27 ( .A(n1201), .Y(n1218) );
  INVX2 U28 ( .A(n1201), .Y(n1219) );
  INVX1 U29 ( .A(n1187), .Y(n1199) );
  INVX1 U30 ( .A(n1165), .Y(N30) );
  INVX1 U31 ( .A(n1169), .Y(N26) );
  INVX1 U32 ( .A(n1163), .Y(N32) );
  INVX1 U33 ( .A(n1166), .Y(N29) );
  INVX1 U34 ( .A(n1167), .Y(N28) );
  INVX1 U35 ( .A(n1168), .Y(N27) );
  INVX1 U36 ( .A(n1170), .Y(N25) );
  INVX1 U37 ( .A(n1171), .Y(N24) );
  INVX1 U38 ( .A(n1172), .Y(N23) );
  INVX1 U39 ( .A(n1173), .Y(N22) );
  INVX1 U40 ( .A(n1174), .Y(N21) );
  INVX1 U41 ( .A(n1175), .Y(N20) );
  INVX1 U42 ( .A(n1176), .Y(N19) );
  INVX1 U43 ( .A(n1177), .Y(N18) );
  INVX1 U44 ( .A(n1178), .Y(N17) );
  INVX1 U45 ( .A(N14), .Y(n1327) );
  INVX1 U46 ( .A(n1320), .Y(n1220) );
  INVX1 U47 ( .A(n1323), .Y(n1185) );
  INVX1 U48 ( .A(n1319), .Y(n1202) );
  INVX2 U49 ( .A(n1202), .Y(n1211) );
  INVX1 U50 ( .A(n1327), .Y(n1179) );
  INVX1 U51 ( .A(n1321), .Y(n1200) );
  INVX1 U52 ( .A(n1220), .Y(n1204) );
  INVX1 U53 ( .A(n1220), .Y(n1203) );
  INVX1 U54 ( .A(N12), .Y(n1323) );
  INVX1 U55 ( .A(n1323), .Y(n1182) );
  INVX1 U56 ( .A(n1323), .Y(n1183) );
  INVX1 U57 ( .A(N13), .Y(n1325) );
  INVX1 U58 ( .A(n1325), .Y(n1181) );
  INVX1 U59 ( .A(n1325), .Y(n1180) );
  INVX1 U60 ( .A(n1321), .Y(n1187) );
  INVX1 U61 ( .A(n1321), .Y(n1188) );
  INVX8 U62 ( .A(n1291), .Y(n1289) );
  INVX1 U63 ( .A(n1319), .Y(n1201) );
  INVX1 U64 ( .A(n86), .Y(n1235) );
  INVX1 U65 ( .A(n87), .Y(n1252) );
  INVX1 U66 ( .A(n88), .Y(n1269) );
  INVX1 U67 ( .A(n89), .Y(n1286) );
  INVX1 U68 ( .A(rst), .Y(n1328) );
  AND2X2 U69 ( .A(write), .B(n1328), .Y(n56) );
  BUFX2 U70 ( .A(n35), .Y(n1) );
  BUFX2 U71 ( .A(n33), .Y(n2) );
  BUFX2 U72 ( .A(n31), .Y(n3) );
  BUFX2 U73 ( .A(n29), .Y(n4) );
  BUFX2 U74 ( .A(n27), .Y(n5) );
  BUFX2 U75 ( .A(n25), .Y(n6) );
  BUFX2 U76 ( .A(n23), .Y(n7) );
  BUFX2 U77 ( .A(n19), .Y(n8) );
  BUFX2 U78 ( .A(n17), .Y(n9) );
  BUFX2 U79 ( .A(n15), .Y(n10) );
  BUFX2 U80 ( .A(n53), .Y(n11) );
  BUFX2 U81 ( .A(n21), .Y(n12) );
  INVX4 U82 ( .A(n56), .Y(n1291) );
  INVX1 U83 ( .A(n54), .Y(n13) );
  INVX4 U84 ( .A(n54), .Y(n55) );
  AND2X2 U85 ( .A(n1289), .B(n136), .Y(n14) );
  INVX1 U86 ( .A(n14), .Y(n15) );
  AND2X2 U87 ( .A(n1289), .B(n138), .Y(n16) );
  INVX1 U88 ( .A(n16), .Y(n17) );
  AND2X2 U89 ( .A(n1289), .B(n140), .Y(n18) );
  INVX1 U90 ( .A(n18), .Y(n19) );
  AND2X2 U91 ( .A(n1289), .B(n87), .Y(n20) );
  INVX1 U92 ( .A(n20), .Y(n21) );
  AND2X2 U93 ( .A(n1289), .B(n142), .Y(n22) );
  INVX1 U94 ( .A(n22), .Y(n23) );
  AND2X2 U95 ( .A(n1289), .B(n144), .Y(n24) );
  INVX1 U96 ( .A(n24), .Y(n25) );
  AND2X2 U97 ( .A(n1289), .B(n146), .Y(n26) );
  INVX1 U98 ( .A(n26), .Y(n27) );
  AND2X2 U99 ( .A(n1289), .B(n148), .Y(n28) );
  INVX1 U100 ( .A(n28), .Y(n29) );
  AND2X2 U101 ( .A(n1289), .B(n150), .Y(n30) );
  INVX1 U102 ( .A(n30), .Y(n31) );
  AND2X2 U103 ( .A(n1289), .B(n152), .Y(n32) );
  INVX1 U104 ( .A(n32), .Y(n33) );
  AND2X2 U105 ( .A(n1289), .B(n154), .Y(n34) );
  INVX1 U106 ( .A(n34), .Y(n35) );
  AND2X2 U107 ( .A(n1290), .B(n88), .Y(n36) );
  INVX1 U108 ( .A(n36), .Y(n37) );
  AND2X2 U109 ( .A(n1290), .B(n156), .Y(n38) );
  INVX1 U110 ( .A(n38), .Y(n39) );
  AND2X2 U111 ( .A(n1290), .B(n158), .Y(n40) );
  INVX1 U112 ( .A(n40), .Y(n41) );
  AND2X2 U113 ( .A(n1290), .B(n160), .Y(n42) );
  INVX1 U114 ( .A(n42), .Y(n43) );
  AND2X2 U115 ( .A(n1290), .B(n162), .Y(n44) );
  INVX1 U116 ( .A(n44), .Y(n45) );
  AND2X2 U117 ( .A(n1290), .B(n164), .Y(n46) );
  INVX1 U118 ( .A(n46), .Y(n47) );
  AND2X2 U119 ( .A(n1290), .B(n166), .Y(n48) );
  INVX1 U120 ( .A(n48), .Y(n49) );
  AND2X2 U121 ( .A(n1290), .B(n168), .Y(n50) );
  INVX1 U122 ( .A(n50), .Y(n51) );
  AND2X2 U123 ( .A(n1289), .B(n89), .Y(n52) );
  INVX1 U124 ( .A(n52), .Y(n53) );
  OR2X2 U125 ( .A(write), .B(rst), .Y(n54) );
  BUFX2 U126 ( .A(n93), .Y(n1221) );
  BUFX2 U127 ( .A(n93), .Y(n1222) );
  BUFX2 U128 ( .A(n97), .Y(n1223) );
  BUFX2 U129 ( .A(n97), .Y(n1224) );
  BUFX2 U130 ( .A(n101), .Y(n1225) );
  BUFX2 U131 ( .A(n101), .Y(n1226) );
  BUFX2 U132 ( .A(n105), .Y(n1227) );
  BUFX2 U133 ( .A(n105), .Y(n1228) );
  BUFX2 U134 ( .A(n109), .Y(n1229) );
  BUFX2 U135 ( .A(n109), .Y(n1230) );
  BUFX2 U136 ( .A(n113), .Y(n1231) );
  BUFX2 U137 ( .A(n113), .Y(n1232) );
  BUFX2 U138 ( .A(n117), .Y(n1233) );
  BUFX2 U139 ( .A(n117), .Y(n1234) );
  BUFX2 U140 ( .A(n119), .Y(n1236) );
  BUFX2 U141 ( .A(n119), .Y(n1237) );
  BUFX2 U142 ( .A(n123), .Y(n1238) );
  BUFX2 U143 ( .A(n123), .Y(n1239) );
  BUFX2 U144 ( .A(n127), .Y(n1240) );
  BUFX2 U145 ( .A(n127), .Y(n1241) );
  BUFX2 U146 ( .A(n131), .Y(n1242) );
  BUFX2 U147 ( .A(n131), .Y(n1243) );
  BUFX2 U148 ( .A(n135), .Y(n1244) );
  BUFX2 U149 ( .A(n135), .Y(n1245) );
  BUFX2 U150 ( .A(n15), .Y(n1246) );
  BUFX2 U151 ( .A(n15), .Y(n1247) );
  BUFX2 U152 ( .A(n17), .Y(n1248) );
  BUFX2 U153 ( .A(n17), .Y(n1249) );
  BUFX2 U154 ( .A(n19), .Y(n1250) );
  BUFX2 U155 ( .A(n19), .Y(n1251) );
  BUFX2 U156 ( .A(n21), .Y(n1253) );
  BUFX2 U157 ( .A(n21), .Y(n1254) );
  BUFX2 U158 ( .A(n23), .Y(n1255) );
  BUFX2 U159 ( .A(n23), .Y(n1256) );
  BUFX2 U160 ( .A(n25), .Y(n1257) );
  BUFX2 U161 ( .A(n25), .Y(n1258) );
  BUFX2 U162 ( .A(n27), .Y(n1259) );
  BUFX2 U163 ( .A(n27), .Y(n1260) );
  BUFX2 U164 ( .A(n29), .Y(n1261) );
  BUFX2 U165 ( .A(n29), .Y(n1262) );
  BUFX2 U166 ( .A(n31), .Y(n1263) );
  BUFX2 U167 ( .A(n31), .Y(n1264) );
  BUFX2 U168 ( .A(n33), .Y(n1265) );
  BUFX2 U169 ( .A(n33), .Y(n1266) );
  BUFX2 U170 ( .A(n35), .Y(n1267) );
  BUFX2 U171 ( .A(n35), .Y(n1268) );
  BUFX2 U172 ( .A(n37), .Y(n1270) );
  BUFX2 U173 ( .A(n37), .Y(n1271) );
  BUFX2 U174 ( .A(n39), .Y(n1272) );
  BUFX2 U175 ( .A(n39), .Y(n1273) );
  BUFX2 U176 ( .A(n41), .Y(n1274) );
  BUFX2 U177 ( .A(n41), .Y(n1275) );
  BUFX2 U178 ( .A(n43), .Y(n1276) );
  BUFX2 U179 ( .A(n43), .Y(n1277) );
  BUFX2 U180 ( .A(n45), .Y(n1278) );
  BUFX2 U181 ( .A(n45), .Y(n1279) );
  BUFX2 U182 ( .A(n47), .Y(n1280) );
  BUFX2 U183 ( .A(n47), .Y(n1281) );
  BUFX2 U184 ( .A(n49), .Y(n1282) );
  BUFX2 U185 ( .A(n49), .Y(n1283) );
  BUFX2 U186 ( .A(n51), .Y(n1284) );
  BUFX2 U187 ( .A(n51), .Y(n1285) );
  BUFX2 U188 ( .A(n53), .Y(n1287) );
  BUFX2 U189 ( .A(n53), .Y(n1288) );
  INVX1 U190 ( .A(n1320), .Y(n1319) );
  INVX1 U191 ( .A(n1325), .Y(n1324) );
  AND2X1 U192 ( .A(n1185), .B(n1321), .Y(n57) );
  INVX1 U193 ( .A(n1322), .Y(n1321) );
  AND2X1 U194 ( .A(n214), .B(n1326), .Y(n58) );
  INVX1 U195 ( .A(n1327), .Y(n1326) );
  BUFX2 U196 ( .A(n1361), .Y(n59) );
  INVX1 U197 ( .A(n59), .Y(n1753) );
  BUFX2 U198 ( .A(n1378), .Y(n60) );
  INVX1 U199 ( .A(n60), .Y(n1770) );
  BUFX2 U200 ( .A(n1395), .Y(n61) );
  INVX1 U201 ( .A(n61), .Y(n1787) );
  BUFX2 U202 ( .A(n1412), .Y(n62) );
  INVX1 U203 ( .A(n62), .Y(n1804) );
  BUFX2 U204 ( .A(n1429), .Y(n63) );
  INVX1 U205 ( .A(n63), .Y(n1821) );
  BUFX2 U206 ( .A(n1590), .Y(n64) );
  INVX1 U207 ( .A(n64), .Y(n1703) );
  BUFX2 U208 ( .A(n1720), .Y(n65) );
  INVX1 U209 ( .A(n65), .Y(n1838) );
  AND2X1 U210 ( .A(n1319), .B(n57), .Y(n66) );
  AND2X1 U211 ( .A(n1324), .B(n58), .Y(n67) );
  AND2X1 U212 ( .A(n1320), .B(n57), .Y(n68) );
  AND2X1 U213 ( .A(n1325), .B(n58), .Y(n69) );
  AND2X2 U214 ( .A(\data_in<0> ), .B(n1290), .Y(n70) );
  AND2X2 U215 ( .A(\data_in<1> ), .B(n1289), .Y(n71) );
  AND2X2 U216 ( .A(\data_in<2> ), .B(n1290), .Y(n72) );
  AND2X2 U217 ( .A(\data_in<3> ), .B(n1290), .Y(n73) );
  AND2X2 U218 ( .A(\data_in<4> ), .B(n1290), .Y(n74) );
  AND2X2 U219 ( .A(\data_in<5> ), .B(n1290), .Y(n75) );
  AND2X2 U220 ( .A(\data_in<6> ), .B(n1290), .Y(n76) );
  AND2X2 U221 ( .A(\data_in<7> ), .B(n1290), .Y(n77) );
  AND2X2 U222 ( .A(\data_in<8> ), .B(n1290), .Y(n78) );
  AND2X2 U223 ( .A(\data_in<9> ), .B(n1290), .Y(n79) );
  AND2X2 U224 ( .A(\data_in<10> ), .B(n1290), .Y(n80) );
  AND2X2 U225 ( .A(\data_in<11> ), .B(n1290), .Y(n81) );
  AND2X2 U226 ( .A(\data_in<12> ), .B(n1290), .Y(n82) );
  AND2X2 U227 ( .A(\data_in<13> ), .B(n1290), .Y(n83) );
  AND2X2 U228 ( .A(\data_in<14> ), .B(n1290), .Y(n84) );
  AND2X2 U229 ( .A(\data_in<15> ), .B(n1290), .Y(n85) );
  AND2X1 U230 ( .A(n67), .B(n1839), .Y(n86) );
  AND2X1 U231 ( .A(n1839), .B(n69), .Y(n87) );
  AND2X1 U232 ( .A(n1839), .B(n1703), .Y(n88) );
  AND2X1 U233 ( .A(n1839), .B(n1838), .Y(n89) );
  AND2X1 U234 ( .A(n66), .B(n67), .Y(n90) );
  INVX1 U235 ( .A(n90), .Y(n91) );
  AND2X1 U236 ( .A(n1289), .B(n90), .Y(n92) );
  INVX1 U237 ( .A(n92), .Y(n93) );
  AND2X1 U238 ( .A(n67), .B(n68), .Y(n94) );
  INVX1 U239 ( .A(n94), .Y(n95) );
  AND2X1 U240 ( .A(n1289), .B(n94), .Y(n96) );
  INVX1 U241 ( .A(n96), .Y(n97) );
  AND2X1 U242 ( .A(n67), .B(n1753), .Y(n98) );
  INVX1 U243 ( .A(n98), .Y(n99) );
  AND2X1 U244 ( .A(n1290), .B(n98), .Y(n100) );
  INVX1 U245 ( .A(n100), .Y(n101) );
  AND2X1 U246 ( .A(n67), .B(n1770), .Y(n102) );
  INVX1 U247 ( .A(n102), .Y(n103) );
  AND2X1 U248 ( .A(n1289), .B(n102), .Y(n104) );
  INVX1 U249 ( .A(n104), .Y(n105) );
  AND2X1 U250 ( .A(n67), .B(n1787), .Y(n106) );
  INVX1 U251 ( .A(n106), .Y(n107) );
  AND2X1 U252 ( .A(n1290), .B(n106), .Y(n108) );
  INVX1 U253 ( .A(n108), .Y(n109) );
  AND2X1 U254 ( .A(n67), .B(n1804), .Y(n110) );
  INVX1 U255 ( .A(n110), .Y(n111) );
  AND2X1 U256 ( .A(n1289), .B(n110), .Y(n112) );
  INVX1 U257 ( .A(n112), .Y(n113) );
  AND2X1 U258 ( .A(n67), .B(n1821), .Y(n114) );
  INVX1 U259 ( .A(n114), .Y(n115) );
  AND2X1 U260 ( .A(n1290), .B(n114), .Y(n116) );
  INVX1 U261 ( .A(n116), .Y(n117) );
  AND2X1 U262 ( .A(n1289), .B(n86), .Y(n118) );
  INVX1 U263 ( .A(n118), .Y(n119) );
  AND2X1 U264 ( .A(n66), .B(n69), .Y(n120) );
  INVX1 U265 ( .A(n120), .Y(n121) );
  AND2X1 U266 ( .A(n1289), .B(n120), .Y(n122) );
  INVX1 U267 ( .A(n122), .Y(n123) );
  AND2X1 U268 ( .A(n68), .B(n69), .Y(n124) );
  INVX1 U269 ( .A(n124), .Y(n125) );
  AND2X1 U270 ( .A(n1289), .B(n124), .Y(n126) );
  INVX1 U271 ( .A(n126), .Y(n127) );
  AND2X1 U272 ( .A(n1753), .B(n69), .Y(n128) );
  INVX1 U273 ( .A(n128), .Y(n129) );
  AND2X1 U274 ( .A(n1289), .B(n128), .Y(n130) );
  INVX1 U275 ( .A(n130), .Y(n131) );
  AND2X1 U276 ( .A(n1770), .B(n69), .Y(n132) );
  INVX1 U277 ( .A(n132), .Y(n133) );
  AND2X1 U278 ( .A(n1289), .B(n132), .Y(n134) );
  INVX1 U279 ( .A(n134), .Y(n135) );
  AND2X1 U280 ( .A(n1787), .B(n69), .Y(n136) );
  INVX1 U281 ( .A(n136), .Y(n137) );
  AND2X1 U282 ( .A(n1804), .B(n69), .Y(n138) );
  INVX1 U283 ( .A(n138), .Y(n139) );
  AND2X1 U284 ( .A(n1821), .B(n69), .Y(n140) );
  INVX1 U285 ( .A(n140), .Y(n141) );
  AND2X1 U286 ( .A(n66), .B(n1703), .Y(n142) );
  INVX1 U287 ( .A(n142), .Y(n143) );
  AND2X1 U288 ( .A(n68), .B(n1703), .Y(n144) );
  INVX1 U289 ( .A(n144), .Y(n145) );
  AND2X1 U290 ( .A(n1753), .B(n1703), .Y(n146) );
  INVX1 U291 ( .A(n146), .Y(n147) );
  AND2X1 U292 ( .A(n1770), .B(n1703), .Y(n148) );
  INVX1 U293 ( .A(n148), .Y(n149) );
  AND2X1 U294 ( .A(n1787), .B(n1703), .Y(n150) );
  INVX1 U295 ( .A(n150), .Y(n151) );
  AND2X1 U296 ( .A(n1804), .B(n1703), .Y(n152) );
  INVX1 U297 ( .A(n152), .Y(n153) );
  AND2X1 U298 ( .A(n1821), .B(n1703), .Y(n154) );
  INVX1 U299 ( .A(n154), .Y(n155) );
  AND2X1 U300 ( .A(n66), .B(n1838), .Y(n156) );
  INVX1 U301 ( .A(n156), .Y(n157) );
  AND2X1 U302 ( .A(n68), .B(n1838), .Y(n158) );
  INVX1 U303 ( .A(n158), .Y(n159) );
  AND2X1 U304 ( .A(n1753), .B(n1838), .Y(n160) );
  INVX1 U305 ( .A(n160), .Y(n161) );
  AND2X1 U306 ( .A(n1770), .B(n1838), .Y(n162) );
  INVX1 U307 ( .A(n162), .Y(n163) );
  AND2X1 U308 ( .A(n1787), .B(n1838), .Y(n164) );
  INVX1 U309 ( .A(n164), .Y(n165) );
  AND2X1 U310 ( .A(n1804), .B(n1838), .Y(n166) );
  INVX1 U311 ( .A(n166), .Y(n167) );
  AND2X1 U312 ( .A(n1821), .B(n1838), .Y(n168) );
  INVX1 U313 ( .A(n168), .Y(n169) );
  MUX2X1 U314 ( .B(n171), .A(n172), .S(n1189), .Y(n170) );
  MUX2X1 U315 ( .B(n174), .A(n175), .S(n1189), .Y(n173) );
  MUX2X1 U316 ( .B(n177), .A(n178), .S(n1189), .Y(n176) );
  MUX2X1 U317 ( .B(n180), .A(n181), .S(n1189), .Y(n179) );
  MUX2X1 U318 ( .B(n183), .A(n184), .S(n1181), .Y(n182) );
  MUX2X1 U319 ( .B(n186), .A(n187), .S(n1189), .Y(n185) );
  MUX2X1 U320 ( .B(n189), .A(n190), .S(n1189), .Y(n188) );
  MUX2X1 U321 ( .B(n192), .A(n193), .S(n1189), .Y(n191) );
  MUX2X1 U322 ( .B(n195), .A(n196), .S(n1189), .Y(n194) );
  MUX2X1 U323 ( .B(n198), .A(n199), .S(n1181), .Y(n197) );
  MUX2X1 U324 ( .B(n201), .A(n202), .S(n1190), .Y(n200) );
  MUX2X1 U325 ( .B(n204), .A(n205), .S(n1190), .Y(n203) );
  MUX2X1 U326 ( .B(n207), .A(n208), .S(n1190), .Y(n206) );
  MUX2X1 U327 ( .B(n210), .A(n211), .S(n1190), .Y(n209) );
  MUX2X1 U328 ( .B(n213), .A(n215), .S(n1181), .Y(n212) );
  MUX2X1 U329 ( .B(n217), .A(n218), .S(n1190), .Y(n216) );
  MUX2X1 U330 ( .B(n220), .A(n221), .S(n1190), .Y(n219) );
  MUX2X1 U331 ( .B(n223), .A(n224), .S(n1190), .Y(n222) );
  MUX2X1 U332 ( .B(n226), .A(n227), .S(n1190), .Y(n225) );
  MUX2X1 U333 ( .B(n229), .A(n230), .S(n1181), .Y(n228) );
  MUX2X1 U334 ( .B(n232), .A(n233), .S(n1190), .Y(n231) );
  MUX2X1 U335 ( .B(n235), .A(n236), .S(n1190), .Y(n234) );
  MUX2X1 U336 ( .B(n238), .A(n239), .S(n1190), .Y(n237) );
  MUX2X1 U337 ( .B(n241), .A(n242), .S(n1190), .Y(n240) );
  MUX2X1 U338 ( .B(n244), .A(n245), .S(n1181), .Y(n243) );
  MUX2X1 U339 ( .B(n247), .A(n248), .S(n1191), .Y(n246) );
  MUX2X1 U340 ( .B(n250), .A(n251), .S(n1191), .Y(n249) );
  MUX2X1 U341 ( .B(n253), .A(n254), .S(n1191), .Y(n252) );
  MUX2X1 U342 ( .B(n256), .A(n257), .S(n1191), .Y(n255) );
  MUX2X1 U343 ( .B(n259), .A(n260), .S(n1181), .Y(n258) );
  MUX2X1 U344 ( .B(n262), .A(n263), .S(n1191), .Y(n261) );
  MUX2X1 U345 ( .B(n265), .A(n266), .S(n1191), .Y(n264) );
  MUX2X1 U346 ( .B(n268), .A(n269), .S(n1191), .Y(n267) );
  MUX2X1 U347 ( .B(n271), .A(n272), .S(n1191), .Y(n270) );
  MUX2X1 U348 ( .B(n274), .A(n275), .S(n1181), .Y(n273) );
  MUX2X1 U349 ( .B(n277), .A(n278), .S(n1191), .Y(n276) );
  MUX2X1 U350 ( .B(n280), .A(n281), .S(n1191), .Y(n279) );
  MUX2X1 U351 ( .B(n283), .A(n284), .S(n1191), .Y(n282) );
  MUX2X1 U352 ( .B(n286), .A(n287), .S(n1191), .Y(n285) );
  MUX2X1 U353 ( .B(n289), .A(n290), .S(n1181), .Y(n288) );
  MUX2X1 U354 ( .B(n292), .A(n293), .S(n1192), .Y(n291) );
  MUX2X1 U355 ( .B(n295), .A(n296), .S(n1192), .Y(n294) );
  MUX2X1 U356 ( .B(n298), .A(n299), .S(n1192), .Y(n297) );
  MUX2X1 U357 ( .B(n301), .A(n302), .S(n1192), .Y(n300) );
  MUX2X1 U358 ( .B(n304), .A(n305), .S(n1181), .Y(n303) );
  MUX2X1 U359 ( .B(n307), .A(n308), .S(n1192), .Y(n306) );
  MUX2X1 U360 ( .B(n310), .A(n311), .S(n1192), .Y(n309) );
  MUX2X1 U361 ( .B(n313), .A(n314), .S(n1192), .Y(n312) );
  MUX2X1 U362 ( .B(n316), .A(n317), .S(n1192), .Y(n315) );
  MUX2X1 U363 ( .B(n319), .A(n320), .S(n1181), .Y(n318) );
  MUX2X1 U364 ( .B(n322), .A(n323), .S(n1192), .Y(n321) );
  MUX2X1 U365 ( .B(n325), .A(n326), .S(n1192), .Y(n324) );
  MUX2X1 U366 ( .B(n328), .A(n329), .S(n1192), .Y(n327) );
  MUX2X1 U367 ( .B(n331), .A(n332), .S(n1192), .Y(n330) );
  MUX2X1 U368 ( .B(n334), .A(n335), .S(n1181), .Y(n333) );
  MUX2X1 U369 ( .B(n337), .A(n338), .S(n1193), .Y(n336) );
  MUX2X1 U370 ( .B(n340), .A(n341), .S(n1193), .Y(n339) );
  MUX2X1 U371 ( .B(n343), .A(n344), .S(n1193), .Y(n342) );
  MUX2X1 U372 ( .B(n346), .A(n347), .S(n1193), .Y(n345) );
  MUX2X1 U373 ( .B(n349), .A(n350), .S(n1181), .Y(n348) );
  MUX2X1 U374 ( .B(n352), .A(n353), .S(n1193), .Y(n351) );
  MUX2X1 U375 ( .B(n355), .A(n356), .S(n1193), .Y(n354) );
  MUX2X1 U376 ( .B(n358), .A(n359), .S(n1193), .Y(n357) );
  MUX2X1 U377 ( .B(n361), .A(n362), .S(n1193), .Y(n360) );
  MUX2X1 U378 ( .B(n364), .A(n365), .S(n1180), .Y(n363) );
  MUX2X1 U379 ( .B(n367), .A(n368), .S(n1193), .Y(n366) );
  MUX2X1 U380 ( .B(n370), .A(n371), .S(n1193), .Y(n369) );
  MUX2X1 U381 ( .B(n373), .A(n374), .S(n1193), .Y(n372) );
  MUX2X1 U382 ( .B(n376), .A(n377), .S(n1193), .Y(n375) );
  MUX2X1 U383 ( .B(n379), .A(n380), .S(n1180), .Y(n378) );
  MUX2X1 U384 ( .B(n382), .A(n383), .S(n1194), .Y(n381) );
  MUX2X1 U385 ( .B(n385), .A(n386), .S(n1194), .Y(n384) );
  MUX2X1 U386 ( .B(n388), .A(n389), .S(n1194), .Y(n387) );
  MUX2X1 U387 ( .B(n391), .A(n392), .S(n1194), .Y(n390) );
  MUX2X1 U388 ( .B(n394), .A(n395), .S(n1180), .Y(n393) );
  MUX2X1 U389 ( .B(n397), .A(n398), .S(n1194), .Y(n396) );
  MUX2X1 U390 ( .B(n400), .A(n401), .S(n1194), .Y(n399) );
  MUX2X1 U391 ( .B(n403), .A(n404), .S(n1194), .Y(n402) );
  MUX2X1 U392 ( .B(n406), .A(n407), .S(n1194), .Y(n405) );
  MUX2X1 U393 ( .B(n409), .A(n410), .S(n1180), .Y(n408) );
  MUX2X1 U394 ( .B(n412), .A(n413), .S(n1194), .Y(n411) );
  MUX2X1 U395 ( .B(n415), .A(n416), .S(n1194), .Y(n414) );
  MUX2X1 U396 ( .B(n418), .A(n419), .S(n1194), .Y(n417) );
  MUX2X1 U397 ( .B(n421), .A(n422), .S(n1194), .Y(n420) );
  MUX2X1 U398 ( .B(n424), .A(n425), .S(n1180), .Y(n423) );
  MUX2X1 U399 ( .B(n427), .A(n428), .S(n1195), .Y(n426) );
  MUX2X1 U400 ( .B(n430), .A(n431), .S(n1195), .Y(n429) );
  MUX2X1 U401 ( .B(n433), .A(n434), .S(n1195), .Y(n432) );
  MUX2X1 U402 ( .B(n436), .A(n437), .S(n1195), .Y(n435) );
  MUX2X1 U403 ( .B(n439), .A(n440), .S(n1180), .Y(n438) );
  MUX2X1 U404 ( .B(n442), .A(n443), .S(n1195), .Y(n441) );
  MUX2X1 U405 ( .B(n445), .A(n446), .S(n1195), .Y(n444) );
  MUX2X1 U406 ( .B(n448), .A(n449), .S(n1195), .Y(n447) );
  MUX2X1 U407 ( .B(n451), .A(n452), .S(n1195), .Y(n450) );
  MUX2X1 U408 ( .B(n454), .A(n455), .S(n1180), .Y(n453) );
  MUX2X1 U409 ( .B(n457), .A(n458), .S(n1195), .Y(n456) );
  MUX2X1 U410 ( .B(n460), .A(n461), .S(n1195), .Y(n459) );
  MUX2X1 U411 ( .B(n463), .A(n464), .S(n1195), .Y(n462) );
  MUX2X1 U412 ( .B(n466), .A(n467), .S(n1195), .Y(n465) );
  MUX2X1 U413 ( .B(n469), .A(n470), .S(n1180), .Y(n468) );
  MUX2X1 U414 ( .B(n472), .A(n473), .S(n1196), .Y(n471) );
  MUX2X1 U415 ( .B(n475), .A(n476), .S(n1196), .Y(n474) );
  MUX2X1 U416 ( .B(n478), .A(n479), .S(n1196), .Y(n477) );
  MUX2X1 U417 ( .B(n481), .A(n482), .S(n1196), .Y(n480) );
  MUX2X1 U418 ( .B(n484), .A(n485), .S(n1180), .Y(n483) );
  MUX2X1 U419 ( .B(n487), .A(n488), .S(n1196), .Y(n486) );
  MUX2X1 U420 ( .B(n490), .A(n491), .S(n1196), .Y(n489) );
  MUX2X1 U421 ( .B(n493), .A(n494), .S(n1196), .Y(n492) );
  MUX2X1 U422 ( .B(n496), .A(n497), .S(n1196), .Y(n495) );
  MUX2X1 U423 ( .B(n499), .A(n500), .S(n1180), .Y(n498) );
  MUX2X1 U424 ( .B(n502), .A(n503), .S(n1196), .Y(n501) );
  MUX2X1 U425 ( .B(n505), .A(n506), .S(n1196), .Y(n504) );
  MUX2X1 U426 ( .B(n508), .A(n509), .S(n1196), .Y(n507) );
  MUX2X1 U427 ( .B(n511), .A(n512), .S(n1196), .Y(n510) );
  MUX2X1 U428 ( .B(n514), .A(n515), .S(n1180), .Y(n513) );
  MUX2X1 U429 ( .B(n517), .A(n518), .S(n1197), .Y(n516) );
  MUX2X1 U430 ( .B(n520), .A(n521), .S(n1197), .Y(n519) );
  MUX2X1 U431 ( .B(n523), .A(n524), .S(n1197), .Y(n522) );
  MUX2X1 U432 ( .B(n526), .A(n527), .S(n1197), .Y(n525) );
  MUX2X1 U433 ( .B(n529), .A(n530), .S(n1180), .Y(n528) );
  MUX2X1 U434 ( .B(n532), .A(n533), .S(n1197), .Y(n531) );
  MUX2X1 U435 ( .B(n535), .A(n536), .S(n1197), .Y(n534) );
  MUX2X1 U436 ( .B(n538), .A(n539), .S(n1197), .Y(n537) );
  MUX2X1 U437 ( .B(n541), .A(n542), .S(n1197), .Y(n540) );
  MUX2X1 U438 ( .B(n544), .A(n545), .S(n1180), .Y(n543) );
  MUX2X1 U439 ( .B(n547), .A(n548), .S(n1197), .Y(n546) );
  MUX2X1 U440 ( .B(n550), .A(n551), .S(n1197), .Y(n549) );
  MUX2X1 U441 ( .B(n553), .A(n554), .S(n1197), .Y(n552) );
  MUX2X1 U442 ( .B(n556), .A(n557), .S(n1197), .Y(n555) );
  MUX2X1 U443 ( .B(n559), .A(n560), .S(n1180), .Y(n558) );
  MUX2X1 U444 ( .B(n562), .A(n563), .S(n1198), .Y(n561) );
  MUX2X1 U445 ( .B(n565), .A(n566), .S(n1198), .Y(n564) );
  MUX2X1 U446 ( .B(n568), .A(n569), .S(n1198), .Y(n567) );
  MUX2X1 U447 ( .B(n571), .A(n572), .S(n1198), .Y(n570) );
  MUX2X1 U448 ( .B(n574), .A(n575), .S(n1181), .Y(n573) );
  MUX2X1 U449 ( .B(n577), .A(n578), .S(n1198), .Y(n576) );
  MUX2X1 U450 ( .B(n580), .A(n581), .S(n1198), .Y(n579) );
  MUX2X1 U451 ( .B(n583), .A(n584), .S(n1198), .Y(n582) );
  MUX2X1 U452 ( .B(n586), .A(n587), .S(n1198), .Y(n585) );
  MUX2X1 U453 ( .B(n589), .A(n590), .S(n1181), .Y(n588) );
  MUX2X1 U454 ( .B(n592), .A(n593), .S(n1198), .Y(n591) );
  MUX2X1 U455 ( .B(n595), .A(n596), .S(n1198), .Y(n594) );
  MUX2X1 U456 ( .B(n598), .A(n599), .S(n1198), .Y(n597) );
  MUX2X1 U457 ( .B(n601), .A(n602), .S(n1198), .Y(n600) );
  MUX2X1 U458 ( .B(n604), .A(n605), .S(n1180), .Y(n603) );
  MUX2X1 U459 ( .B(n607), .A(n608), .S(n1199), .Y(n606) );
  MUX2X1 U460 ( .B(n610), .A(n611), .S(n1199), .Y(n609) );
  MUX2X1 U461 ( .B(n613), .A(n614), .S(n1199), .Y(n612) );
  MUX2X1 U462 ( .B(n616), .A(n617), .S(n1199), .Y(n615) );
  MUX2X1 U463 ( .B(n619), .A(n620), .S(n1180), .Y(n618) );
  MUX2X1 U464 ( .B(n622), .A(n623), .S(n1199), .Y(n621) );
  MUX2X1 U465 ( .B(n625), .A(n626), .S(n1199), .Y(n624) );
  MUX2X1 U466 ( .B(n628), .A(n629), .S(n1199), .Y(n627) );
  MUX2X1 U467 ( .B(n631), .A(n632), .S(n1199), .Y(n630) );
  MUX2X1 U468 ( .B(n634), .A(n635), .S(n1181), .Y(n633) );
  MUX2X1 U469 ( .B(n637), .A(n638), .S(n1199), .Y(n636) );
  MUX2X1 U470 ( .B(n640), .A(n641), .S(n1199), .Y(n639) );
  MUX2X1 U471 ( .B(n643), .A(n644), .S(n1199), .Y(n642) );
  MUX2X1 U472 ( .B(n646), .A(n647), .S(n1199), .Y(n645) );
  MUX2X1 U473 ( .B(n649), .A(n650), .S(n1181), .Y(n648) );
  MUX2X1 U474 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1205), .Y(n172) );
  MUX2X1 U475 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1205), .Y(n171) );
  MUX2X1 U476 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1205), .Y(n175) );
  MUX2X1 U477 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1205), .Y(n174) );
  MUX2X1 U478 ( .B(n173), .A(n170), .S(n1186), .Y(n184) );
  MUX2X1 U479 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1206), .Y(n178) );
  MUX2X1 U480 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1206), .Y(n177) );
  MUX2X1 U481 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1206), .Y(n181) );
  MUX2X1 U482 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1206), .Y(n180) );
  MUX2X1 U483 ( .B(n179), .A(n176), .S(n1186), .Y(n183) );
  MUX2X1 U484 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1206), .Y(n187) );
  MUX2X1 U485 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1206), .Y(n186) );
  MUX2X1 U486 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1206), .Y(n190) );
  MUX2X1 U487 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1206), .Y(n189) );
  MUX2X1 U488 ( .B(n188), .A(n185), .S(n1186), .Y(n199) );
  MUX2X1 U489 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1206), .Y(n193) );
  MUX2X1 U490 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1206), .Y(n192) );
  MUX2X1 U491 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1206), .Y(n196) );
  MUX2X1 U492 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1206), .Y(n195) );
  MUX2X1 U493 ( .B(n194), .A(n191), .S(n1186), .Y(n198) );
  MUX2X1 U494 ( .B(n197), .A(n182), .S(n1179), .Y(n1163) );
  MUX2X1 U495 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1207), .Y(n202) );
  MUX2X1 U496 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1207), .Y(n201) );
  MUX2X1 U497 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1207), .Y(n205) );
  MUX2X1 U498 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1207), .Y(n204) );
  MUX2X1 U499 ( .B(n203), .A(n200), .S(n1186), .Y(n215) );
  MUX2X1 U500 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1207), .Y(n208) );
  MUX2X1 U501 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1207), .Y(n207) );
  MUX2X1 U502 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1207), .Y(n211) );
  MUX2X1 U503 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1207), .Y(n210) );
  MUX2X1 U504 ( .B(n209), .A(n206), .S(n1186), .Y(n213) );
  MUX2X1 U505 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1207), .Y(n218) );
  MUX2X1 U506 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1207), .Y(n217) );
  MUX2X1 U507 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1207), .Y(n221) );
  MUX2X1 U508 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1207), .Y(n220) );
  MUX2X1 U509 ( .B(n219), .A(n216), .S(n1186), .Y(n230) );
  MUX2X1 U510 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1219), .Y(n224) );
  MUX2X1 U511 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1205), .Y(n223) );
  MUX2X1 U512 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1206), .Y(n227) );
  MUX2X1 U513 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1207), .Y(n226) );
  MUX2X1 U514 ( .B(n225), .A(n222), .S(n1186), .Y(n229) );
  MUX2X1 U515 ( .B(n228), .A(n212), .S(n1179), .Y(n1164) );
  MUX2X1 U516 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1211), .Y(n233) );
  MUX2X1 U517 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1206), .Y(n232) );
  MUX2X1 U518 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1209), .Y(n236) );
  MUX2X1 U519 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1216), .Y(n235) );
  MUX2X1 U520 ( .B(n234), .A(n231), .S(n1186), .Y(n245) );
  MUX2X1 U521 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1213), .Y(n239) );
  MUX2X1 U522 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1208), .Y(n238) );
  MUX2X1 U523 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1219), .Y(n242) );
  MUX2X1 U524 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1207), .Y(n241) );
  MUX2X1 U525 ( .B(n240), .A(n237), .S(n1186), .Y(n244) );
  MUX2X1 U526 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1209), .Y(n248) );
  MUX2X1 U527 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1211), .Y(n247) );
  MUX2X1 U528 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1205), .Y(n251) );
  MUX2X1 U529 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1206), .Y(n250) );
  MUX2X1 U530 ( .B(n249), .A(n246), .S(n1186), .Y(n260) );
  MUX2X1 U531 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1205), .Y(n254) );
  MUX2X1 U532 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1213), .Y(n253) );
  MUX2X1 U533 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1219), .Y(n257) );
  MUX2X1 U534 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1219), .Y(n256) );
  MUX2X1 U535 ( .B(n255), .A(n252), .S(n1186), .Y(n259) );
  MUX2X1 U536 ( .B(n258), .A(n243), .S(n1179), .Y(n1165) );
  MUX2X1 U537 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1211), .Y(n263) );
  MUX2X1 U538 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1213), .Y(n262) );
  MUX2X1 U539 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1209), .Y(n266) );
  MUX2X1 U540 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1205), .Y(n265) );
  MUX2X1 U541 ( .B(n264), .A(n261), .S(n1185), .Y(n275) );
  MUX2X1 U542 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1211), .Y(n269) );
  MUX2X1 U543 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1207), .Y(n268) );
  MUX2X1 U544 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1219), .Y(n272) );
  MUX2X1 U545 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1208), .Y(n271) );
  MUX2X1 U546 ( .B(n270), .A(n267), .S(n1185), .Y(n274) );
  MUX2X1 U547 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1208), .Y(n278) );
  MUX2X1 U548 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1208), .Y(n277) );
  MUX2X1 U549 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1207), .Y(n281) );
  MUX2X1 U550 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1219), .Y(n280) );
  MUX2X1 U551 ( .B(n279), .A(n276), .S(n1185), .Y(n290) );
  MUX2X1 U552 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1211), .Y(n284) );
  MUX2X1 U553 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1209), .Y(n283) );
  MUX2X1 U554 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1206), .Y(n287) );
  MUX2X1 U555 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1219), .Y(n286) );
  MUX2X1 U556 ( .B(n285), .A(n282), .S(n1185), .Y(n289) );
  MUX2X1 U557 ( .B(n288), .A(n273), .S(n1179), .Y(n1166) );
  MUX2X1 U558 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1219), .Y(n293) );
  MUX2X1 U559 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1215), .Y(n292) );
  MUX2X1 U560 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1205), .Y(n296) );
  MUX2X1 U561 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1217), .Y(n295) );
  MUX2X1 U562 ( .B(n294), .A(n291), .S(n1185), .Y(n305) );
  MUX2X1 U563 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1208), .Y(n299) );
  MUX2X1 U564 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1212), .Y(n298) );
  MUX2X1 U565 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1209), .Y(n302) );
  MUX2X1 U566 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1218), .Y(n301) );
  MUX2X1 U567 ( .B(n300), .A(n297), .S(n1185), .Y(n304) );
  MUX2X1 U568 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1219), .Y(n308) );
  MUX2X1 U569 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1207), .Y(n307) );
  MUX2X1 U570 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1206), .Y(n311) );
  MUX2X1 U571 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1213), .Y(n310) );
  MUX2X1 U572 ( .B(n309), .A(n306), .S(n1185), .Y(n320) );
  MUX2X1 U573 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1208), .Y(n314) );
  MUX2X1 U574 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1208), .Y(n313) );
  MUX2X1 U575 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1208), .Y(n317) );
  MUX2X1 U576 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1208), .Y(n316) );
  MUX2X1 U577 ( .B(n315), .A(n312), .S(n1185), .Y(n319) );
  MUX2X1 U578 ( .B(n318), .A(n303), .S(n1179), .Y(n1167) );
  MUX2X1 U579 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1208), .Y(n323) );
  MUX2X1 U580 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1208), .Y(n322) );
  MUX2X1 U581 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1208), .Y(n326) );
  MUX2X1 U582 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1208), .Y(n325) );
  MUX2X1 U583 ( .B(n324), .A(n321), .S(n1185), .Y(n335) );
  MUX2X1 U584 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1208), .Y(n329) );
  MUX2X1 U585 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1208), .Y(n328) );
  MUX2X1 U586 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1208), .Y(n332) );
  MUX2X1 U587 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1208), .Y(n331) );
  MUX2X1 U588 ( .B(n330), .A(n327), .S(n1185), .Y(n334) );
  MUX2X1 U589 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1209), .Y(n338) );
  MUX2X1 U590 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1209), .Y(n337) );
  MUX2X1 U591 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1209), .Y(n341) );
  MUX2X1 U592 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1209), .Y(n340) );
  MUX2X1 U593 ( .B(n339), .A(n336), .S(n1185), .Y(n350) );
  MUX2X1 U594 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1209), .Y(n344) );
  MUX2X1 U595 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1209), .Y(n343) );
  MUX2X1 U596 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1209), .Y(n347) );
  MUX2X1 U597 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1209), .Y(n346) );
  MUX2X1 U598 ( .B(n345), .A(n342), .S(n1185), .Y(n349) );
  MUX2X1 U599 ( .B(n348), .A(n333), .S(n1179), .Y(n1168) );
  MUX2X1 U600 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1209), .Y(n353) );
  MUX2X1 U601 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1209), .Y(n352) );
  MUX2X1 U602 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1209), .Y(n356) );
  MUX2X1 U603 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1209), .Y(n355) );
  MUX2X1 U604 ( .B(n354), .A(n351), .S(n1184), .Y(n365) );
  MUX2X1 U605 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1210), .Y(n359) );
  MUX2X1 U606 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1210), .Y(n358) );
  MUX2X1 U607 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1210), .Y(n362) );
  MUX2X1 U608 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1210), .Y(n361) );
  MUX2X1 U609 ( .B(n360), .A(n357), .S(n1184), .Y(n364) );
  MUX2X1 U610 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1210), .Y(n368) );
  MUX2X1 U611 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1210), .Y(n367) );
  MUX2X1 U612 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1210), .Y(n371) );
  MUX2X1 U613 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1210), .Y(n370) );
  MUX2X1 U614 ( .B(n369), .A(n366), .S(n1184), .Y(n380) );
  MUX2X1 U615 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1210), .Y(n374) );
  MUX2X1 U616 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1210), .Y(n373) );
  MUX2X1 U617 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1210), .Y(n377) );
  MUX2X1 U618 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1210), .Y(n376) );
  MUX2X1 U619 ( .B(n375), .A(n372), .S(n1184), .Y(n379) );
  MUX2X1 U620 ( .B(n378), .A(n363), .S(n1179), .Y(n1169) );
  MUX2X1 U621 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1211), .Y(n383) );
  MUX2X1 U622 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1211), .Y(n382) );
  MUX2X1 U623 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1211), .Y(n386) );
  MUX2X1 U624 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1211), .Y(n385) );
  MUX2X1 U625 ( .B(n384), .A(n381), .S(n1184), .Y(n395) );
  MUX2X1 U626 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1211), .Y(n389) );
  MUX2X1 U627 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1211), .Y(n388) );
  MUX2X1 U628 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1211), .Y(n392) );
  MUX2X1 U629 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1211), .Y(n391) );
  MUX2X1 U630 ( .B(n390), .A(n387), .S(n1184), .Y(n394) );
  MUX2X1 U631 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1211), .Y(n398) );
  MUX2X1 U632 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1211), .Y(n397) );
  MUX2X1 U633 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1211), .Y(n401) );
  MUX2X1 U634 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1211), .Y(n400) );
  MUX2X1 U635 ( .B(n399), .A(n396), .S(n1184), .Y(n410) );
  MUX2X1 U636 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1211), .Y(n404) );
  MUX2X1 U637 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1211), .Y(n403) );
  MUX2X1 U638 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1211), .Y(n407) );
  MUX2X1 U639 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1211), .Y(n406) );
  MUX2X1 U640 ( .B(n405), .A(n402), .S(n1184), .Y(n409) );
  MUX2X1 U641 ( .B(n408), .A(n393), .S(n1179), .Y(n1170) );
  MUX2X1 U642 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1211), .Y(n413) );
  MUX2X1 U643 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1211), .Y(n412) );
  MUX2X1 U644 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1211), .Y(n416) );
  MUX2X1 U645 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1211), .Y(n415) );
  MUX2X1 U646 ( .B(n414), .A(n411), .S(n1184), .Y(n425) );
  MUX2X1 U647 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1210), .Y(n419) );
  MUX2X1 U648 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1210), .Y(n418) );
  MUX2X1 U649 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1211), .Y(n422) );
  MUX2X1 U650 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1211), .Y(n421) );
  MUX2X1 U651 ( .B(n420), .A(n417), .S(n1184), .Y(n424) );
  MUX2X1 U652 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1215), .Y(n428) );
  MUX2X1 U653 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1215), .Y(n427) );
  MUX2X1 U654 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1205), .Y(n431) );
  MUX2X1 U655 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1214), .Y(n430) );
  MUX2X1 U656 ( .B(n429), .A(n426), .S(n1184), .Y(n440) );
  MUX2X1 U657 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1214), .Y(n434) );
  MUX2X1 U658 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1205), .Y(n433) );
  MUX2X1 U659 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1205), .Y(n437) );
  MUX2X1 U660 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1215), .Y(n436) );
  MUX2X1 U661 ( .B(n435), .A(n432), .S(n1184), .Y(n439) );
  MUX2X1 U662 ( .B(n438), .A(n423), .S(n1179), .Y(n1171) );
  MUX2X1 U663 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1215), .Y(n443) );
  MUX2X1 U664 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1205), .Y(n442) );
  MUX2X1 U665 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1214), .Y(n446) );
  MUX2X1 U666 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1214), .Y(n445) );
  MUX2X1 U667 ( .B(n444), .A(n441), .S(n1183), .Y(n455) );
  MUX2X1 U668 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1212), .Y(n449) );
  MUX2X1 U669 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1212), .Y(n448) );
  MUX2X1 U670 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1212), .Y(n452) );
  MUX2X1 U671 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1212), .Y(n451) );
  MUX2X1 U672 ( .B(n450), .A(n447), .S(n1183), .Y(n454) );
  MUX2X1 U673 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1212), .Y(n458) );
  MUX2X1 U674 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1212), .Y(n457) );
  MUX2X1 U675 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1212), .Y(n461) );
  MUX2X1 U676 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1212), .Y(n460) );
  MUX2X1 U677 ( .B(n459), .A(n456), .S(n1183), .Y(n470) );
  MUX2X1 U678 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1212), .Y(n464) );
  MUX2X1 U679 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1212), .Y(n463) );
  MUX2X1 U680 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1212), .Y(n467) );
  MUX2X1 U681 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1212), .Y(n466) );
  MUX2X1 U682 ( .B(n465), .A(n462), .S(n1183), .Y(n469) );
  MUX2X1 U683 ( .B(n468), .A(n453), .S(n1179), .Y(n1172) );
  MUX2X1 U684 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1213), .Y(n473) );
  MUX2X1 U685 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1213), .Y(n472) );
  MUX2X1 U686 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1213), .Y(n476) );
  MUX2X1 U687 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1213), .Y(n475) );
  MUX2X1 U688 ( .B(n474), .A(n471), .S(n1183), .Y(n485) );
  MUX2X1 U689 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1213), .Y(n479) );
  MUX2X1 U690 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1213), .Y(n478) );
  MUX2X1 U691 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1213), .Y(n482) );
  MUX2X1 U692 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1213), .Y(n481) );
  MUX2X1 U693 ( .B(n480), .A(n477), .S(n1183), .Y(n484) );
  MUX2X1 U694 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1213), .Y(n488) );
  MUX2X1 U695 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1213), .Y(n487) );
  MUX2X1 U696 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1213), .Y(n491) );
  MUX2X1 U697 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1213), .Y(n490) );
  MUX2X1 U698 ( .B(n489), .A(n486), .S(n1183), .Y(n500) );
  MUX2X1 U699 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1214), .Y(n494) );
  MUX2X1 U700 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1214), .Y(n493) );
  MUX2X1 U701 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1214), .Y(n497) );
  MUX2X1 U702 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1214), .Y(n496) );
  MUX2X1 U703 ( .B(n495), .A(n492), .S(n1183), .Y(n499) );
  MUX2X1 U704 ( .B(n498), .A(n483), .S(n1179), .Y(n1173) );
  MUX2X1 U705 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1214), .Y(n503) );
  MUX2X1 U706 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1214), .Y(n502) );
  MUX2X1 U707 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1214), .Y(n506) );
  MUX2X1 U708 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1214), .Y(n505) );
  MUX2X1 U709 ( .B(n504), .A(n501), .S(n1183), .Y(n515) );
  MUX2X1 U710 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1214), .Y(n509) );
  MUX2X1 U711 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1214), .Y(n508) );
  MUX2X1 U712 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1214), .Y(n512) );
  MUX2X1 U713 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1214), .Y(n511) );
  MUX2X1 U714 ( .B(n510), .A(n507), .S(n1183), .Y(n514) );
  MUX2X1 U715 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1215), .Y(n518) );
  MUX2X1 U716 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1215), .Y(n517) );
  MUX2X1 U717 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1215), .Y(n521) );
  MUX2X1 U718 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1215), .Y(n520) );
  MUX2X1 U719 ( .B(n519), .A(n516), .S(n1183), .Y(n530) );
  MUX2X1 U720 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1215), .Y(n524) );
  MUX2X1 U721 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1215), .Y(n523) );
  MUX2X1 U722 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1215), .Y(n527) );
  MUX2X1 U723 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1215), .Y(n526) );
  MUX2X1 U724 ( .B(n525), .A(n522), .S(n1183), .Y(n529) );
  MUX2X1 U725 ( .B(n528), .A(n513), .S(n1179), .Y(n1174) );
  MUX2X1 U726 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1215), .Y(n533) );
  MUX2X1 U727 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1215), .Y(n532) );
  MUX2X1 U728 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1215), .Y(n536) );
  MUX2X1 U729 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1215), .Y(n535) );
  MUX2X1 U730 ( .B(n534), .A(n531), .S(n1182), .Y(n545) );
  MUX2X1 U731 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1219), .Y(n539) );
  MUX2X1 U732 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1205), .Y(n538) );
  MUX2X1 U733 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1219), .Y(n542) );
  MUX2X1 U734 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1219), .Y(n541) );
  MUX2X1 U735 ( .B(n540), .A(n537), .S(n1182), .Y(n544) );
  MUX2X1 U736 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1205), .Y(n548) );
  MUX2X1 U737 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1219), .Y(n547) );
  MUX2X1 U738 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1205), .Y(n551) );
  MUX2X1 U739 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1213), .Y(n550) );
  MUX2X1 U740 ( .B(n549), .A(n546), .S(n1182), .Y(n560) );
  MUX2X1 U741 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1211), .Y(n554) );
  MUX2X1 U742 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1217), .Y(n553) );
  MUX2X1 U743 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1205), .Y(n557) );
  MUX2X1 U744 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1219), .Y(n556) );
  MUX2X1 U745 ( .B(n555), .A(n552), .S(n1182), .Y(n559) );
  MUX2X1 U746 ( .B(n558), .A(n543), .S(n1179), .Y(n1175) );
  MUX2X1 U747 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1216), .Y(n563) );
  MUX2X1 U748 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1216), .Y(n562) );
  MUX2X1 U749 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1216), .Y(n566) );
  MUX2X1 U750 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1216), .Y(n565) );
  MUX2X1 U751 ( .B(n564), .A(n561), .S(n1182), .Y(n575) );
  MUX2X1 U752 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1216), .Y(n569) );
  MUX2X1 U753 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1216), .Y(n568) );
  MUX2X1 U754 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1216), .Y(n572) );
  MUX2X1 U755 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1216), .Y(n571) );
  MUX2X1 U756 ( .B(n570), .A(n567), .S(n1182), .Y(n574) );
  MUX2X1 U757 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1216), .Y(n578) );
  MUX2X1 U758 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1216), .Y(n577) );
  MUX2X1 U759 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1216), .Y(n581) );
  MUX2X1 U760 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1216), .Y(n580) );
  MUX2X1 U761 ( .B(n579), .A(n576), .S(n1182), .Y(n590) );
  MUX2X1 U762 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1217), .Y(n584) );
  MUX2X1 U763 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1217), .Y(n583) );
  MUX2X1 U764 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1217), .Y(n587) );
  MUX2X1 U765 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1217), .Y(n586) );
  MUX2X1 U766 ( .B(n585), .A(n582), .S(n1182), .Y(n589) );
  MUX2X1 U767 ( .B(n588), .A(n573), .S(n1179), .Y(n1176) );
  MUX2X1 U768 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1217), .Y(n593) );
  MUX2X1 U769 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1217), .Y(n592) );
  MUX2X1 U770 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1217), .Y(n596) );
  MUX2X1 U771 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1217), .Y(n595) );
  MUX2X1 U772 ( .B(n594), .A(n591), .S(n1182), .Y(n605) );
  MUX2X1 U773 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1217), .Y(n599) );
  MUX2X1 U774 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1217), .Y(n598) );
  MUX2X1 U775 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1217), .Y(n602) );
  MUX2X1 U776 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1217), .Y(n601) );
  MUX2X1 U777 ( .B(n600), .A(n597), .S(n1182), .Y(n604) );
  MUX2X1 U778 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1218), .Y(n608) );
  MUX2X1 U779 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1218), .Y(n607) );
  MUX2X1 U780 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1218), .Y(n611) );
  MUX2X1 U781 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1218), .Y(n610) );
  MUX2X1 U782 ( .B(n609), .A(n606), .S(n1182), .Y(n620) );
  MUX2X1 U783 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1218), .Y(n614) );
  MUX2X1 U784 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1218), .Y(n613) );
  MUX2X1 U785 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1218), .Y(n617) );
  MUX2X1 U786 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1218), .Y(n616) );
  MUX2X1 U787 ( .B(n615), .A(n612), .S(n1182), .Y(n619) );
  MUX2X1 U788 ( .B(n618), .A(n603), .S(n1179), .Y(n1177) );
  MUX2X1 U789 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1218), .Y(n623) );
  MUX2X1 U790 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1218), .Y(n622) );
  MUX2X1 U791 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1218), .Y(n626) );
  MUX2X1 U792 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1218), .Y(n625) );
  MUX2X1 U793 ( .B(n624), .A(n621), .S(n1182), .Y(n635) );
  MUX2X1 U794 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1219), .Y(n629) );
  MUX2X1 U795 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1219), .Y(n628) );
  MUX2X1 U796 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1219), .Y(n632) );
  MUX2X1 U797 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1219), .Y(n631) );
  MUX2X1 U798 ( .B(n630), .A(n627), .S(n1183), .Y(n634) );
  MUX2X1 U799 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1219), .Y(n638) );
  MUX2X1 U800 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1219), .Y(n637) );
  MUX2X1 U801 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1219), .Y(n641) );
  MUX2X1 U802 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1219), .Y(n640) );
  MUX2X1 U803 ( .B(n639), .A(n636), .S(n1182), .Y(n650) );
  MUX2X1 U804 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1219), .Y(n644) );
  MUX2X1 U805 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1219), .Y(n643) );
  MUX2X1 U806 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1219), .Y(n647) );
  MUX2X1 U807 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1219), .Y(n646) );
  MUX2X1 U808 ( .B(n645), .A(n642), .S(n1183), .Y(n649) );
  MUX2X1 U809 ( .B(n648), .A(n633), .S(n1179), .Y(n1178) );
  INVX1 U810 ( .A(N11), .Y(n1322) );
  INVX1 U811 ( .A(N10), .Y(n1320) );
  INVX8 U812 ( .A(n1291), .Y(n1290) );
  INVX8 U813 ( .A(n70), .Y(n1292) );
  INVX8 U814 ( .A(n70), .Y(n1293) );
  INVX8 U815 ( .A(n71), .Y(n1294) );
  INVX8 U816 ( .A(n71), .Y(n1295) );
  INVX8 U817 ( .A(n72), .Y(n1296) );
  INVX8 U818 ( .A(n72), .Y(n1297) );
  INVX8 U819 ( .A(n73), .Y(n1298) );
  INVX8 U820 ( .A(n73), .Y(n1299) );
  INVX8 U821 ( .A(n74), .Y(n1300) );
  INVX8 U822 ( .A(n74), .Y(n1301) );
  INVX8 U823 ( .A(n75), .Y(n1302) );
  INVX8 U824 ( .A(n75), .Y(n1303) );
  INVX8 U825 ( .A(n76), .Y(n1304) );
  INVX8 U826 ( .A(n76), .Y(n1305) );
  INVX8 U827 ( .A(n77), .Y(n1306) );
  INVX8 U828 ( .A(n77), .Y(n1307) );
  INVX8 U829 ( .A(n78), .Y(n1308) );
  INVX8 U830 ( .A(n78), .Y(n1309) );
  INVX8 U831 ( .A(n79), .Y(n1310) );
  INVX8 U832 ( .A(n79), .Y(n1311) );
  INVX8 U833 ( .A(n80), .Y(n1312) );
  INVX8 U834 ( .A(n80), .Y(n1313) );
  INVX8 U835 ( .A(n81), .Y(n1314) );
  INVX8 U836 ( .A(n82), .Y(n1315) );
  INVX8 U837 ( .A(n83), .Y(n1316) );
  INVX8 U838 ( .A(n84), .Y(n1317) );
  INVX8 U839 ( .A(n85), .Y(n1318) );
  AND2X2 U840 ( .A(N32), .B(n55), .Y(\data_out<0> ) );
  AND2X2 U841 ( .A(n55), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U842 ( .A(n55), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U843 ( .A(N29), .B(n55), .Y(\data_out<3> ) );
  AND2X2 U844 ( .A(N28), .B(n55), .Y(\data_out<4> ) );
  AND2X2 U845 ( .A(N27), .B(n55), .Y(\data_out<5> ) );
  AND2X2 U846 ( .A(N26), .B(n55), .Y(\data_out<6> ) );
  AND2X2 U847 ( .A(N25), .B(n55), .Y(\data_out<7> ) );
  AND2X2 U848 ( .A(N24), .B(n55), .Y(\data_out<8> ) );
  AND2X2 U849 ( .A(N23), .B(n55), .Y(\data_out<9> ) );
  AND2X2 U850 ( .A(N22), .B(n13), .Y(\data_out<10> ) );
  AND2X2 U851 ( .A(N21), .B(n55), .Y(\data_out<11> ) );
  AND2X2 U852 ( .A(N20), .B(n55), .Y(\data_out<12> ) );
  AND2X2 U853 ( .A(n13), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U854 ( .A(N18), .B(n13), .Y(\data_out<14> ) );
  AND2X2 U855 ( .A(N17), .B(n55), .Y(\data_out<15> ) );
  NAND2X1 U856 ( .A(\mem<31><0> ), .B(n1221), .Y(n1329) );
  OAI21X1 U857 ( .A(n91), .B(n1292), .C(n1329), .Y(n651) );
  NAND2X1 U858 ( .A(\mem<31><1> ), .B(n1221), .Y(n1330) );
  OAI21X1 U859 ( .A(n1295), .B(n91), .C(n1330), .Y(n652) );
  NAND2X1 U860 ( .A(\mem<31><2> ), .B(n1221), .Y(n1331) );
  OAI21X1 U861 ( .A(n1297), .B(n91), .C(n1331), .Y(n653) );
  NAND2X1 U862 ( .A(\mem<31><3> ), .B(n1221), .Y(n1332) );
  OAI21X1 U863 ( .A(n1299), .B(n91), .C(n1332), .Y(n654) );
  NAND2X1 U864 ( .A(\mem<31><4> ), .B(n1221), .Y(n1333) );
  OAI21X1 U865 ( .A(n1301), .B(n91), .C(n1333), .Y(n655) );
  NAND2X1 U866 ( .A(\mem<31><5> ), .B(n1221), .Y(n1334) );
  OAI21X1 U867 ( .A(n1303), .B(n91), .C(n1334), .Y(n656) );
  NAND2X1 U868 ( .A(\mem<31><6> ), .B(n1221), .Y(n1335) );
  OAI21X1 U869 ( .A(n1305), .B(n91), .C(n1335), .Y(n657) );
  NAND2X1 U870 ( .A(\mem<31><7> ), .B(n1221), .Y(n1336) );
  OAI21X1 U871 ( .A(n1307), .B(n91), .C(n1336), .Y(n658) );
  NAND2X1 U872 ( .A(\mem<31><8> ), .B(n1222), .Y(n1337) );
  OAI21X1 U873 ( .A(n1309), .B(n91), .C(n1337), .Y(n659) );
  NAND2X1 U874 ( .A(\mem<31><9> ), .B(n1222), .Y(n1338) );
  OAI21X1 U875 ( .A(n1311), .B(n91), .C(n1338), .Y(n660) );
  NAND2X1 U876 ( .A(\mem<31><10> ), .B(n1222), .Y(n1339) );
  OAI21X1 U877 ( .A(n1313), .B(n91), .C(n1339), .Y(n661) );
  NAND2X1 U878 ( .A(\mem<31><11> ), .B(n1222), .Y(n1340) );
  OAI21X1 U879 ( .A(n1314), .B(n91), .C(n1340), .Y(n662) );
  NAND2X1 U880 ( .A(\mem<31><12> ), .B(n1222), .Y(n1341) );
  OAI21X1 U881 ( .A(n1315), .B(n91), .C(n1341), .Y(n663) );
  NAND2X1 U882 ( .A(\mem<31><13> ), .B(n1222), .Y(n1342) );
  OAI21X1 U883 ( .A(n1316), .B(n91), .C(n1342), .Y(n664) );
  NAND2X1 U884 ( .A(\mem<31><14> ), .B(n1222), .Y(n1343) );
  OAI21X1 U885 ( .A(n1317), .B(n91), .C(n1343), .Y(n665) );
  NAND2X1 U886 ( .A(\mem<31><15> ), .B(n1222), .Y(n1344) );
  OAI21X1 U887 ( .A(n1318), .B(n91), .C(n1344), .Y(n666) );
  NAND2X1 U888 ( .A(\mem<30><0> ), .B(n1223), .Y(n1345) );
  OAI21X1 U889 ( .A(n95), .B(n1292), .C(n1345), .Y(n667) );
  NAND2X1 U890 ( .A(\mem<30><1> ), .B(n1223), .Y(n1346) );
  OAI21X1 U891 ( .A(n95), .B(n1295), .C(n1346), .Y(n668) );
  NAND2X1 U892 ( .A(\mem<30><2> ), .B(n1223), .Y(n1347) );
  OAI21X1 U893 ( .A(n95), .B(n1297), .C(n1347), .Y(n669) );
  NAND2X1 U894 ( .A(\mem<30><3> ), .B(n1223), .Y(n1348) );
  OAI21X1 U895 ( .A(n95), .B(n1299), .C(n1348), .Y(n670) );
  NAND2X1 U896 ( .A(\mem<30><4> ), .B(n1223), .Y(n1349) );
  OAI21X1 U897 ( .A(n95), .B(n1301), .C(n1349), .Y(n671) );
  NAND2X1 U898 ( .A(\mem<30><5> ), .B(n1223), .Y(n1350) );
  OAI21X1 U899 ( .A(n95), .B(n1303), .C(n1350), .Y(n672) );
  NAND2X1 U900 ( .A(\mem<30><6> ), .B(n1223), .Y(n1351) );
  OAI21X1 U901 ( .A(n95), .B(n1305), .C(n1351), .Y(n673) );
  NAND2X1 U902 ( .A(\mem<30><7> ), .B(n1223), .Y(n1352) );
  OAI21X1 U903 ( .A(n95), .B(n1307), .C(n1352), .Y(n674) );
  NAND2X1 U904 ( .A(\mem<30><8> ), .B(n1224), .Y(n1353) );
  OAI21X1 U905 ( .A(n95), .B(n1308), .C(n1353), .Y(n675) );
  NAND2X1 U906 ( .A(\mem<30><9> ), .B(n1224), .Y(n1354) );
  OAI21X1 U907 ( .A(n95), .B(n1310), .C(n1354), .Y(n676) );
  NAND2X1 U908 ( .A(\mem<30><10> ), .B(n1224), .Y(n1355) );
  OAI21X1 U909 ( .A(n95), .B(n1312), .C(n1355), .Y(n677) );
  NAND2X1 U910 ( .A(\mem<30><11> ), .B(n1224), .Y(n1356) );
  OAI21X1 U911 ( .A(n95), .B(n1314), .C(n1356), .Y(n678) );
  NAND2X1 U912 ( .A(\mem<30><12> ), .B(n1224), .Y(n1357) );
  OAI21X1 U913 ( .A(n95), .B(n1315), .C(n1357), .Y(n679) );
  NAND2X1 U914 ( .A(\mem<30><13> ), .B(n1224), .Y(n1358) );
  OAI21X1 U915 ( .A(n95), .B(n1316), .C(n1358), .Y(n680) );
  NAND2X1 U916 ( .A(\mem<30><14> ), .B(n1224), .Y(n1359) );
  OAI21X1 U917 ( .A(n95), .B(n1317), .C(n1359), .Y(n681) );
  NAND2X1 U918 ( .A(\mem<30><15> ), .B(n1224), .Y(n1360) );
  OAI21X1 U919 ( .A(n95), .B(n1318), .C(n1360), .Y(n682) );
  NAND3X1 U920 ( .A(n1319), .B(n1185), .C(n1322), .Y(n1361) );
  NAND2X1 U921 ( .A(\mem<29><0> ), .B(n1225), .Y(n1362) );
  OAI21X1 U922 ( .A(n99), .B(n1292), .C(n1362), .Y(n683) );
  NAND2X1 U923 ( .A(\mem<29><1> ), .B(n1225), .Y(n1363) );
  OAI21X1 U924 ( .A(n99), .B(n1294), .C(n1363), .Y(n684) );
  NAND2X1 U925 ( .A(\mem<29><2> ), .B(n1225), .Y(n1364) );
  OAI21X1 U926 ( .A(n99), .B(n1296), .C(n1364), .Y(n685) );
  NAND2X1 U927 ( .A(\mem<29><3> ), .B(n1225), .Y(n1365) );
  OAI21X1 U928 ( .A(n99), .B(n1298), .C(n1365), .Y(n686) );
  NAND2X1 U929 ( .A(\mem<29><4> ), .B(n1225), .Y(n1366) );
  OAI21X1 U930 ( .A(n99), .B(n1300), .C(n1366), .Y(n687) );
  NAND2X1 U931 ( .A(\mem<29><5> ), .B(n1225), .Y(n1367) );
  OAI21X1 U932 ( .A(n99), .B(n1302), .C(n1367), .Y(n688) );
  NAND2X1 U933 ( .A(\mem<29><6> ), .B(n1225), .Y(n1368) );
  OAI21X1 U934 ( .A(n99), .B(n1304), .C(n1368), .Y(n689) );
  NAND2X1 U935 ( .A(\mem<29><7> ), .B(n1225), .Y(n1369) );
  OAI21X1 U936 ( .A(n99), .B(n1306), .C(n1369), .Y(n690) );
  NAND2X1 U937 ( .A(\mem<29><8> ), .B(n1226), .Y(n1370) );
  OAI21X1 U938 ( .A(n99), .B(n1309), .C(n1370), .Y(n691) );
  NAND2X1 U939 ( .A(\mem<29><9> ), .B(n1226), .Y(n1371) );
  OAI21X1 U940 ( .A(n99), .B(n1311), .C(n1371), .Y(n692) );
  NAND2X1 U941 ( .A(\mem<29><10> ), .B(n1226), .Y(n1372) );
  OAI21X1 U942 ( .A(n99), .B(n1313), .C(n1372), .Y(n693) );
  NAND2X1 U943 ( .A(\mem<29><11> ), .B(n1226), .Y(n1373) );
  OAI21X1 U944 ( .A(n99), .B(n1314), .C(n1373), .Y(n694) );
  NAND2X1 U945 ( .A(\mem<29><12> ), .B(n1226), .Y(n1374) );
  OAI21X1 U946 ( .A(n99), .B(n1315), .C(n1374), .Y(n695) );
  NAND2X1 U947 ( .A(\mem<29><13> ), .B(n1226), .Y(n1375) );
  OAI21X1 U948 ( .A(n99), .B(n1316), .C(n1375), .Y(n696) );
  NAND2X1 U949 ( .A(\mem<29><14> ), .B(n1226), .Y(n1376) );
  OAI21X1 U950 ( .A(n99), .B(n1317), .C(n1376), .Y(n697) );
  NAND2X1 U951 ( .A(\mem<29><15> ), .B(n1226), .Y(n1377) );
  OAI21X1 U952 ( .A(n99), .B(n1318), .C(n1377), .Y(n698) );
  NAND3X1 U953 ( .A(n1185), .B(n1322), .C(n1320), .Y(n1378) );
  NAND2X1 U954 ( .A(\mem<28><0> ), .B(n1227), .Y(n1379) );
  OAI21X1 U955 ( .A(n103), .B(n1292), .C(n1379), .Y(n699) );
  NAND2X1 U956 ( .A(\mem<28><1> ), .B(n1227), .Y(n1380) );
  OAI21X1 U957 ( .A(n103), .B(n1295), .C(n1380), .Y(n700) );
  NAND2X1 U958 ( .A(\mem<28><2> ), .B(n1227), .Y(n1381) );
  OAI21X1 U959 ( .A(n103), .B(n1297), .C(n1381), .Y(n701) );
  NAND2X1 U960 ( .A(\mem<28><3> ), .B(n1227), .Y(n1382) );
  OAI21X1 U961 ( .A(n103), .B(n1299), .C(n1382), .Y(n702) );
  NAND2X1 U962 ( .A(\mem<28><4> ), .B(n1227), .Y(n1383) );
  OAI21X1 U963 ( .A(n103), .B(n1301), .C(n1383), .Y(n703) );
  NAND2X1 U964 ( .A(\mem<28><5> ), .B(n1227), .Y(n1384) );
  OAI21X1 U965 ( .A(n103), .B(n1303), .C(n1384), .Y(n704) );
  NAND2X1 U966 ( .A(\mem<28><6> ), .B(n1227), .Y(n1385) );
  OAI21X1 U967 ( .A(n103), .B(n1305), .C(n1385), .Y(n705) );
  NAND2X1 U968 ( .A(\mem<28><7> ), .B(n1227), .Y(n1386) );
  OAI21X1 U969 ( .A(n103), .B(n1307), .C(n1386), .Y(n706) );
  NAND2X1 U970 ( .A(\mem<28><8> ), .B(n1228), .Y(n1387) );
  OAI21X1 U971 ( .A(n103), .B(n1308), .C(n1387), .Y(n707) );
  NAND2X1 U972 ( .A(\mem<28><9> ), .B(n1228), .Y(n1388) );
  OAI21X1 U973 ( .A(n103), .B(n1310), .C(n1388), .Y(n708) );
  NAND2X1 U974 ( .A(\mem<28><10> ), .B(n1228), .Y(n1389) );
  OAI21X1 U975 ( .A(n103), .B(n1312), .C(n1389), .Y(n709) );
  NAND2X1 U976 ( .A(\mem<28><11> ), .B(n1228), .Y(n1390) );
  OAI21X1 U977 ( .A(n103), .B(n1314), .C(n1390), .Y(n710) );
  NAND2X1 U978 ( .A(\mem<28><12> ), .B(n1228), .Y(n1391) );
  OAI21X1 U979 ( .A(n103), .B(n1315), .C(n1391), .Y(n711) );
  NAND2X1 U980 ( .A(\mem<28><13> ), .B(n1228), .Y(n1392) );
  OAI21X1 U981 ( .A(n103), .B(n1316), .C(n1392), .Y(n712) );
  NAND2X1 U982 ( .A(\mem<28><14> ), .B(n1228), .Y(n1393) );
  OAI21X1 U983 ( .A(n103), .B(n1317), .C(n1393), .Y(n713) );
  NAND2X1 U984 ( .A(\mem<28><15> ), .B(n1228), .Y(n1394) );
  OAI21X1 U985 ( .A(n103), .B(n1318), .C(n1394), .Y(n714) );
  NAND3X1 U986 ( .A(n1319), .B(n1321), .C(n1323), .Y(n1395) );
  NAND2X1 U987 ( .A(\mem<27><0> ), .B(n1229), .Y(n1396) );
  OAI21X1 U988 ( .A(n107), .B(n1292), .C(n1396), .Y(n715) );
  NAND2X1 U989 ( .A(\mem<27><1> ), .B(n1229), .Y(n1397) );
  OAI21X1 U990 ( .A(n107), .B(n1294), .C(n1397), .Y(n716) );
  NAND2X1 U991 ( .A(\mem<27><2> ), .B(n1229), .Y(n1398) );
  OAI21X1 U992 ( .A(n107), .B(n1296), .C(n1398), .Y(n717) );
  NAND2X1 U993 ( .A(\mem<27><3> ), .B(n1229), .Y(n1399) );
  OAI21X1 U994 ( .A(n107), .B(n1298), .C(n1399), .Y(n718) );
  NAND2X1 U995 ( .A(\mem<27><4> ), .B(n1229), .Y(n1400) );
  OAI21X1 U996 ( .A(n107), .B(n1300), .C(n1400), .Y(n719) );
  NAND2X1 U997 ( .A(\mem<27><5> ), .B(n1229), .Y(n1401) );
  OAI21X1 U998 ( .A(n107), .B(n1302), .C(n1401), .Y(n720) );
  NAND2X1 U999 ( .A(\mem<27><6> ), .B(n1229), .Y(n1402) );
  OAI21X1 U1000 ( .A(n107), .B(n1304), .C(n1402), .Y(n721) );
  NAND2X1 U1001 ( .A(\mem<27><7> ), .B(n1229), .Y(n1403) );
  OAI21X1 U1002 ( .A(n107), .B(n1306), .C(n1403), .Y(n722) );
  NAND2X1 U1003 ( .A(\mem<27><8> ), .B(n1230), .Y(n1404) );
  OAI21X1 U1004 ( .A(n107), .B(n1309), .C(n1404), .Y(n723) );
  NAND2X1 U1005 ( .A(\mem<27><9> ), .B(n1230), .Y(n1405) );
  OAI21X1 U1006 ( .A(n107), .B(n1311), .C(n1405), .Y(n724) );
  NAND2X1 U1007 ( .A(\mem<27><10> ), .B(n1230), .Y(n1406) );
  OAI21X1 U1008 ( .A(n107), .B(n1313), .C(n1406), .Y(n725) );
  NAND2X1 U1009 ( .A(\mem<27><11> ), .B(n1230), .Y(n1407) );
  OAI21X1 U1010 ( .A(n107), .B(n1314), .C(n1407), .Y(n726) );
  NAND2X1 U1011 ( .A(\mem<27><12> ), .B(n1230), .Y(n1408) );
  OAI21X1 U1012 ( .A(n107), .B(n1315), .C(n1408), .Y(n727) );
  NAND2X1 U1013 ( .A(\mem<27><13> ), .B(n1230), .Y(n1409) );
  OAI21X1 U1014 ( .A(n107), .B(n1316), .C(n1409), .Y(n728) );
  NAND2X1 U1015 ( .A(\mem<27><14> ), .B(n1230), .Y(n1410) );
  OAI21X1 U1016 ( .A(n107), .B(n1317), .C(n1410), .Y(n729) );
  NAND2X1 U1017 ( .A(\mem<27><15> ), .B(n1230), .Y(n1411) );
  OAI21X1 U1018 ( .A(n107), .B(n1318), .C(n1411), .Y(n730) );
  NAND3X1 U1019 ( .A(n1323), .B(n1321), .C(n1320), .Y(n1412) );
  NAND2X1 U1020 ( .A(\mem<26><0> ), .B(n1231), .Y(n1413) );
  OAI21X1 U1021 ( .A(n111), .B(n1292), .C(n1413), .Y(n731) );
  NAND2X1 U1022 ( .A(\mem<26><1> ), .B(n1231), .Y(n1414) );
  OAI21X1 U1023 ( .A(n111), .B(n1295), .C(n1414), .Y(n732) );
  NAND2X1 U1024 ( .A(\mem<26><2> ), .B(n1231), .Y(n1415) );
  OAI21X1 U1025 ( .A(n111), .B(n1297), .C(n1415), .Y(n733) );
  NAND2X1 U1026 ( .A(\mem<26><3> ), .B(n1231), .Y(n1416) );
  OAI21X1 U1027 ( .A(n111), .B(n1299), .C(n1416), .Y(n734) );
  NAND2X1 U1028 ( .A(\mem<26><4> ), .B(n1231), .Y(n1417) );
  OAI21X1 U1029 ( .A(n111), .B(n1301), .C(n1417), .Y(n735) );
  NAND2X1 U1030 ( .A(\mem<26><5> ), .B(n1231), .Y(n1418) );
  OAI21X1 U1031 ( .A(n111), .B(n1303), .C(n1418), .Y(n736) );
  NAND2X1 U1032 ( .A(\mem<26><6> ), .B(n1231), .Y(n1419) );
  OAI21X1 U1033 ( .A(n111), .B(n1305), .C(n1419), .Y(n737) );
  NAND2X1 U1034 ( .A(\mem<26><7> ), .B(n1231), .Y(n1420) );
  OAI21X1 U1035 ( .A(n111), .B(n1307), .C(n1420), .Y(n738) );
  NAND2X1 U1036 ( .A(\mem<26><8> ), .B(n1232), .Y(n1421) );
  OAI21X1 U1037 ( .A(n111), .B(n1308), .C(n1421), .Y(n739) );
  NAND2X1 U1038 ( .A(\mem<26><9> ), .B(n1232), .Y(n1422) );
  OAI21X1 U1039 ( .A(n111), .B(n1310), .C(n1422), .Y(n740) );
  NAND2X1 U1040 ( .A(\mem<26><10> ), .B(n1232), .Y(n1423) );
  OAI21X1 U1041 ( .A(n111), .B(n1312), .C(n1423), .Y(n741) );
  NAND2X1 U1042 ( .A(\mem<26><11> ), .B(n1232), .Y(n1424) );
  OAI21X1 U1043 ( .A(n111), .B(n1314), .C(n1424), .Y(n742) );
  NAND2X1 U1044 ( .A(\mem<26><12> ), .B(n1232), .Y(n1425) );
  OAI21X1 U1045 ( .A(n111), .B(n1315), .C(n1425), .Y(n743) );
  NAND2X1 U1046 ( .A(\mem<26><13> ), .B(n1232), .Y(n1426) );
  OAI21X1 U1047 ( .A(n111), .B(n1316), .C(n1426), .Y(n744) );
  NAND2X1 U1048 ( .A(\mem<26><14> ), .B(n1232), .Y(n1427) );
  OAI21X1 U1049 ( .A(n111), .B(n1317), .C(n1427), .Y(n745) );
  NAND2X1 U1050 ( .A(\mem<26><15> ), .B(n1232), .Y(n1428) );
  OAI21X1 U1051 ( .A(n111), .B(n1318), .C(n1428), .Y(n746) );
  NAND3X1 U1052 ( .A(n1319), .B(n1323), .C(n1322), .Y(n1429) );
  NAND2X1 U1053 ( .A(\mem<25><0> ), .B(n1233), .Y(n1430) );
  OAI21X1 U1054 ( .A(n115), .B(n1292), .C(n1430), .Y(n747) );
  NAND2X1 U1055 ( .A(\mem<25><1> ), .B(n1233), .Y(n1431) );
  OAI21X1 U1056 ( .A(n115), .B(n1294), .C(n1431), .Y(n748) );
  NAND2X1 U1057 ( .A(\mem<25><2> ), .B(n1233), .Y(n1432) );
  OAI21X1 U1058 ( .A(n115), .B(n1296), .C(n1432), .Y(n749) );
  NAND2X1 U1059 ( .A(\mem<25><3> ), .B(n1233), .Y(n1433) );
  OAI21X1 U1060 ( .A(n115), .B(n1298), .C(n1433), .Y(n750) );
  NAND2X1 U1061 ( .A(\mem<25><4> ), .B(n1233), .Y(n1434) );
  OAI21X1 U1062 ( .A(n115), .B(n1300), .C(n1434), .Y(n751) );
  NAND2X1 U1063 ( .A(\mem<25><5> ), .B(n1233), .Y(n1435) );
  OAI21X1 U1064 ( .A(n115), .B(n1302), .C(n1435), .Y(n752) );
  NAND2X1 U1065 ( .A(\mem<25><6> ), .B(n1233), .Y(n1436) );
  OAI21X1 U1066 ( .A(n115), .B(n1304), .C(n1436), .Y(n753) );
  NAND2X1 U1067 ( .A(\mem<25><7> ), .B(n1233), .Y(n1437) );
  OAI21X1 U1068 ( .A(n115), .B(n1306), .C(n1437), .Y(n754) );
  NAND2X1 U1069 ( .A(\mem<25><8> ), .B(n1234), .Y(n1438) );
  OAI21X1 U1070 ( .A(n115), .B(n1309), .C(n1438), .Y(n755) );
  NAND2X1 U1071 ( .A(\mem<25><9> ), .B(n1234), .Y(n1439) );
  OAI21X1 U1072 ( .A(n115), .B(n1311), .C(n1439), .Y(n756) );
  NAND2X1 U1073 ( .A(\mem<25><10> ), .B(n1234), .Y(n1440) );
  OAI21X1 U1074 ( .A(n115), .B(n1313), .C(n1440), .Y(n757) );
  NAND2X1 U1075 ( .A(\mem<25><11> ), .B(n1234), .Y(n1441) );
  OAI21X1 U1076 ( .A(n115), .B(n1314), .C(n1441), .Y(n758) );
  NAND2X1 U1077 ( .A(\mem<25><12> ), .B(n1234), .Y(n1442) );
  OAI21X1 U1078 ( .A(n115), .B(n1315), .C(n1442), .Y(n759) );
  NAND2X1 U1079 ( .A(\mem<25><13> ), .B(n1234), .Y(n1443) );
  OAI21X1 U1080 ( .A(n115), .B(n1316), .C(n1443), .Y(n760) );
  NAND2X1 U1081 ( .A(\mem<25><14> ), .B(n1234), .Y(n1444) );
  OAI21X1 U1082 ( .A(n115), .B(n1317), .C(n1444), .Y(n761) );
  NAND2X1 U1083 ( .A(\mem<25><15> ), .B(n1234), .Y(n1445) );
  OAI21X1 U1084 ( .A(n115), .B(n1318), .C(n1445), .Y(n762) );
  NOR3X1 U1085 ( .A(n1319), .B(n1321), .C(n1185), .Y(n1839) );
  NAND2X1 U1086 ( .A(\mem<24><0> ), .B(n1236), .Y(n1446) );
  OAI21X1 U1087 ( .A(n1235), .B(n1292), .C(n1446), .Y(n763) );
  NAND2X1 U1088 ( .A(\mem<24><1> ), .B(n1236), .Y(n1447) );
  OAI21X1 U1089 ( .A(n1235), .B(n1294), .C(n1447), .Y(n764) );
  NAND2X1 U1090 ( .A(\mem<24><2> ), .B(n1236), .Y(n1448) );
  OAI21X1 U1091 ( .A(n1235), .B(n1296), .C(n1448), .Y(n765) );
  NAND2X1 U1092 ( .A(\mem<24><3> ), .B(n1236), .Y(n1449) );
  OAI21X1 U1093 ( .A(n1235), .B(n1298), .C(n1449), .Y(n766) );
  NAND2X1 U1094 ( .A(\mem<24><4> ), .B(n1236), .Y(n1450) );
  OAI21X1 U1095 ( .A(n1235), .B(n1300), .C(n1450), .Y(n767) );
  NAND2X1 U1096 ( .A(\mem<24><5> ), .B(n1236), .Y(n1451) );
  OAI21X1 U1097 ( .A(n1235), .B(n1302), .C(n1451), .Y(n768) );
  NAND2X1 U1098 ( .A(\mem<24><6> ), .B(n1236), .Y(n1452) );
  OAI21X1 U1099 ( .A(n1235), .B(n1304), .C(n1452), .Y(n769) );
  NAND2X1 U1100 ( .A(\mem<24><7> ), .B(n1236), .Y(n1453) );
  OAI21X1 U1101 ( .A(n1235), .B(n1306), .C(n1453), .Y(n770) );
  NAND2X1 U1102 ( .A(\mem<24><8> ), .B(n1237), .Y(n1454) );
  OAI21X1 U1103 ( .A(n1235), .B(n1308), .C(n1454), .Y(n771) );
  NAND2X1 U1104 ( .A(\mem<24><9> ), .B(n1237), .Y(n1455) );
  OAI21X1 U1105 ( .A(n1235), .B(n1310), .C(n1455), .Y(n772) );
  NAND2X1 U1106 ( .A(\mem<24><10> ), .B(n1237), .Y(n1456) );
  OAI21X1 U1107 ( .A(n1235), .B(n1312), .C(n1456), .Y(n773) );
  NAND2X1 U1108 ( .A(\mem<24><11> ), .B(n1237), .Y(n1457) );
  OAI21X1 U1109 ( .A(n1235), .B(n1314), .C(n1457), .Y(n774) );
  NAND2X1 U1110 ( .A(\mem<24><12> ), .B(n1237), .Y(n1458) );
  OAI21X1 U1111 ( .A(n1235), .B(n1315), .C(n1458), .Y(n775) );
  NAND2X1 U1112 ( .A(\mem<24><13> ), .B(n1237), .Y(n1459) );
  OAI21X1 U1113 ( .A(n1235), .B(n1316), .C(n1459), .Y(n776) );
  NAND2X1 U1114 ( .A(\mem<24><14> ), .B(n1237), .Y(n1460) );
  OAI21X1 U1115 ( .A(n1235), .B(n1317), .C(n1460), .Y(n777) );
  NAND2X1 U1116 ( .A(\mem<24><15> ), .B(n1237), .Y(n1461) );
  OAI21X1 U1117 ( .A(n1235), .B(n1318), .C(n1461), .Y(n778) );
  NAND2X1 U1118 ( .A(\mem<23><0> ), .B(n1238), .Y(n1462) );
  OAI21X1 U1119 ( .A(n121), .B(n1292), .C(n1462), .Y(n779) );
  NAND2X1 U1120 ( .A(\mem<23><1> ), .B(n1238), .Y(n1463) );
  OAI21X1 U1121 ( .A(n121), .B(n1295), .C(n1463), .Y(n780) );
  NAND2X1 U1122 ( .A(\mem<23><2> ), .B(n1238), .Y(n1464) );
  OAI21X1 U1123 ( .A(n121), .B(n1297), .C(n1464), .Y(n781) );
  NAND2X1 U1124 ( .A(\mem<23><3> ), .B(n1238), .Y(n1465) );
  OAI21X1 U1125 ( .A(n121), .B(n1299), .C(n1465), .Y(n782) );
  NAND2X1 U1126 ( .A(\mem<23><4> ), .B(n1238), .Y(n1466) );
  OAI21X1 U1127 ( .A(n121), .B(n1301), .C(n1466), .Y(n783) );
  NAND2X1 U1128 ( .A(\mem<23><5> ), .B(n1238), .Y(n1467) );
  OAI21X1 U1129 ( .A(n121), .B(n1303), .C(n1467), .Y(n784) );
  NAND2X1 U1130 ( .A(\mem<23><6> ), .B(n1238), .Y(n1468) );
  OAI21X1 U1131 ( .A(n121), .B(n1305), .C(n1468), .Y(n785) );
  NAND2X1 U1132 ( .A(\mem<23><7> ), .B(n1238), .Y(n1469) );
  OAI21X1 U1133 ( .A(n121), .B(n1307), .C(n1469), .Y(n786) );
  NAND2X1 U1134 ( .A(\mem<23><8> ), .B(n1239), .Y(n1470) );
  OAI21X1 U1135 ( .A(n121), .B(n1309), .C(n1470), .Y(n787) );
  NAND2X1 U1136 ( .A(\mem<23><9> ), .B(n1239), .Y(n1471) );
  OAI21X1 U1137 ( .A(n121), .B(n1311), .C(n1471), .Y(n788) );
  NAND2X1 U1138 ( .A(\mem<23><10> ), .B(n1239), .Y(n1472) );
  OAI21X1 U1139 ( .A(n121), .B(n1313), .C(n1472), .Y(n789) );
  NAND2X1 U1140 ( .A(\mem<23><11> ), .B(n1239), .Y(n1473) );
  OAI21X1 U1141 ( .A(n121), .B(n1314), .C(n1473), .Y(n790) );
  NAND2X1 U1142 ( .A(\mem<23><12> ), .B(n1239), .Y(n1474) );
  OAI21X1 U1143 ( .A(n121), .B(n1315), .C(n1474), .Y(n791) );
  NAND2X1 U1144 ( .A(\mem<23><13> ), .B(n1239), .Y(n1475) );
  OAI21X1 U1145 ( .A(n121), .B(n1316), .C(n1475), .Y(n792) );
  NAND2X1 U1146 ( .A(\mem<23><14> ), .B(n1239), .Y(n1476) );
  OAI21X1 U1147 ( .A(n121), .B(n1317), .C(n1476), .Y(n793) );
  NAND2X1 U1148 ( .A(\mem<23><15> ), .B(n1239), .Y(n1477) );
  OAI21X1 U1149 ( .A(n121), .B(n1318), .C(n1477), .Y(n794) );
  NAND2X1 U1150 ( .A(\mem<22><0> ), .B(n1240), .Y(n1478) );
  OAI21X1 U1151 ( .A(n125), .B(n1292), .C(n1478), .Y(n795) );
  NAND2X1 U1152 ( .A(\mem<22><1> ), .B(n1240), .Y(n1479) );
  OAI21X1 U1153 ( .A(n125), .B(n1295), .C(n1479), .Y(n796) );
  NAND2X1 U1154 ( .A(\mem<22><2> ), .B(n1240), .Y(n1480) );
  OAI21X1 U1155 ( .A(n125), .B(n1297), .C(n1480), .Y(n797) );
  NAND2X1 U1156 ( .A(\mem<22><3> ), .B(n1240), .Y(n1481) );
  OAI21X1 U1157 ( .A(n125), .B(n1299), .C(n1481), .Y(n798) );
  NAND2X1 U1158 ( .A(\mem<22><4> ), .B(n1240), .Y(n1482) );
  OAI21X1 U1159 ( .A(n125), .B(n1301), .C(n1482), .Y(n799) );
  NAND2X1 U1160 ( .A(\mem<22><5> ), .B(n1240), .Y(n1483) );
  OAI21X1 U1161 ( .A(n125), .B(n1303), .C(n1483), .Y(n800) );
  NAND2X1 U1162 ( .A(\mem<22><6> ), .B(n1240), .Y(n1484) );
  OAI21X1 U1163 ( .A(n125), .B(n1305), .C(n1484), .Y(n801) );
  NAND2X1 U1164 ( .A(\mem<22><7> ), .B(n1240), .Y(n1485) );
  OAI21X1 U1165 ( .A(n125), .B(n1307), .C(n1485), .Y(n802) );
  NAND2X1 U1166 ( .A(\mem<22><8> ), .B(n1241), .Y(n1486) );
  OAI21X1 U1167 ( .A(n125), .B(n1309), .C(n1486), .Y(n803) );
  NAND2X1 U1168 ( .A(\mem<22><9> ), .B(n1241), .Y(n1487) );
  OAI21X1 U1169 ( .A(n125), .B(n1311), .C(n1487), .Y(n804) );
  NAND2X1 U1170 ( .A(\mem<22><10> ), .B(n1241), .Y(n1488) );
  OAI21X1 U1171 ( .A(n125), .B(n1313), .C(n1488), .Y(n805) );
  NAND2X1 U1172 ( .A(\mem<22><11> ), .B(n1241), .Y(n1489) );
  OAI21X1 U1173 ( .A(n125), .B(n1314), .C(n1489), .Y(n806) );
  NAND2X1 U1174 ( .A(\mem<22><12> ), .B(n1241), .Y(n1490) );
  OAI21X1 U1175 ( .A(n125), .B(n1315), .C(n1490), .Y(n807) );
  NAND2X1 U1177 ( .A(\mem<22><13> ), .B(n1241), .Y(n1491) );
  OAI21X1 U1178 ( .A(n125), .B(n1316), .C(n1491), .Y(n808) );
  NAND2X1 U1179 ( .A(\mem<22><14> ), .B(n1241), .Y(n1492) );
  OAI21X1 U1180 ( .A(n125), .B(n1317), .C(n1492), .Y(n809) );
  NAND2X1 U1181 ( .A(\mem<22><15> ), .B(n1241), .Y(n1493) );
  OAI21X1 U1182 ( .A(n125), .B(n1318), .C(n1493), .Y(n810) );
  NAND2X1 U1183 ( .A(\mem<21><0> ), .B(n1242), .Y(n1494) );
  OAI21X1 U1184 ( .A(n129), .B(n1292), .C(n1494), .Y(n811) );
  NAND2X1 U1185 ( .A(\mem<21><1> ), .B(n1242), .Y(n1495) );
  OAI21X1 U1186 ( .A(n129), .B(n1295), .C(n1495), .Y(n812) );
  NAND2X1 U1187 ( .A(\mem<21><2> ), .B(n1242), .Y(n1496) );
  OAI21X1 U1188 ( .A(n129), .B(n1297), .C(n1496), .Y(n813) );
  NAND2X1 U1189 ( .A(\mem<21><3> ), .B(n1242), .Y(n1497) );
  OAI21X1 U1190 ( .A(n129), .B(n1299), .C(n1497), .Y(n814) );
  NAND2X1 U1191 ( .A(\mem<21><4> ), .B(n1242), .Y(n1498) );
  OAI21X1 U1192 ( .A(n129), .B(n1301), .C(n1498), .Y(n815) );
  NAND2X1 U1193 ( .A(\mem<21><5> ), .B(n1242), .Y(n1499) );
  OAI21X1 U1194 ( .A(n129), .B(n1303), .C(n1499), .Y(n816) );
  NAND2X1 U1195 ( .A(\mem<21><6> ), .B(n1242), .Y(n1500) );
  OAI21X1 U1196 ( .A(n129), .B(n1305), .C(n1500), .Y(n817) );
  NAND2X1 U1197 ( .A(\mem<21><7> ), .B(n1242), .Y(n1501) );
  OAI21X1 U1198 ( .A(n129), .B(n1307), .C(n1501), .Y(n818) );
  NAND2X1 U1199 ( .A(\mem<21><8> ), .B(n1243), .Y(n1502) );
  OAI21X1 U1200 ( .A(n129), .B(n1309), .C(n1502), .Y(n819) );
  NAND2X1 U1201 ( .A(\mem<21><9> ), .B(n1243), .Y(n1503) );
  OAI21X1 U1202 ( .A(n129), .B(n1311), .C(n1503), .Y(n820) );
  NAND2X1 U1203 ( .A(\mem<21><10> ), .B(n1243), .Y(n1504) );
  OAI21X1 U1204 ( .A(n129), .B(n1313), .C(n1504), .Y(n821) );
  NAND2X1 U1205 ( .A(\mem<21><11> ), .B(n1243), .Y(n1505) );
  OAI21X1 U1206 ( .A(n129), .B(n1314), .C(n1505), .Y(n822) );
  NAND2X1 U1207 ( .A(\mem<21><12> ), .B(n1243), .Y(n1506) );
  OAI21X1 U1208 ( .A(n129), .B(n1315), .C(n1506), .Y(n823) );
  NAND2X1 U1209 ( .A(\mem<21><13> ), .B(n1243), .Y(n1507) );
  OAI21X1 U1210 ( .A(n129), .B(n1316), .C(n1507), .Y(n824) );
  NAND2X1 U1211 ( .A(\mem<21><14> ), .B(n1243), .Y(n1508) );
  OAI21X1 U1212 ( .A(n129), .B(n1317), .C(n1508), .Y(n825) );
  NAND2X1 U1213 ( .A(\mem<21><15> ), .B(n1243), .Y(n1509) );
  OAI21X1 U1214 ( .A(n129), .B(n1318), .C(n1509), .Y(n826) );
  NAND2X1 U1215 ( .A(\mem<20><0> ), .B(n1244), .Y(n1510) );
  OAI21X1 U1216 ( .A(n133), .B(n1292), .C(n1510), .Y(n827) );
  NAND2X1 U1217 ( .A(\mem<20><1> ), .B(n1244), .Y(n1511) );
  OAI21X1 U1218 ( .A(n133), .B(n1295), .C(n1511), .Y(n828) );
  NAND2X1 U1219 ( .A(\mem<20><2> ), .B(n1244), .Y(n1512) );
  OAI21X1 U1220 ( .A(n133), .B(n1297), .C(n1512), .Y(n829) );
  NAND2X1 U1221 ( .A(\mem<20><3> ), .B(n1244), .Y(n1513) );
  OAI21X1 U1222 ( .A(n133), .B(n1299), .C(n1513), .Y(n830) );
  NAND2X1 U1223 ( .A(\mem<20><4> ), .B(n1244), .Y(n1514) );
  OAI21X1 U1224 ( .A(n133), .B(n1301), .C(n1514), .Y(n831) );
  NAND2X1 U1225 ( .A(\mem<20><5> ), .B(n1244), .Y(n1515) );
  OAI21X1 U1226 ( .A(n133), .B(n1303), .C(n1515), .Y(n832) );
  NAND2X1 U1227 ( .A(\mem<20><6> ), .B(n1244), .Y(n1516) );
  OAI21X1 U1228 ( .A(n133), .B(n1305), .C(n1516), .Y(n833) );
  NAND2X1 U1229 ( .A(\mem<20><7> ), .B(n1244), .Y(n1517) );
  OAI21X1 U1230 ( .A(n133), .B(n1307), .C(n1517), .Y(n834) );
  NAND2X1 U1231 ( .A(\mem<20><8> ), .B(n1245), .Y(n1518) );
  OAI21X1 U1232 ( .A(n133), .B(n1309), .C(n1518), .Y(n835) );
  NAND2X1 U1233 ( .A(\mem<20><9> ), .B(n1245), .Y(n1519) );
  OAI21X1 U1234 ( .A(n133), .B(n1311), .C(n1519), .Y(n836) );
  NAND2X1 U1235 ( .A(\mem<20><10> ), .B(n1245), .Y(n1520) );
  OAI21X1 U1236 ( .A(n133), .B(n1313), .C(n1520), .Y(n837) );
  NAND2X1 U1237 ( .A(\mem<20><11> ), .B(n1245), .Y(n1521) );
  OAI21X1 U1238 ( .A(n133), .B(n1314), .C(n1521), .Y(n838) );
  NAND2X1 U1239 ( .A(\mem<20><12> ), .B(n1245), .Y(n1522) );
  OAI21X1 U1240 ( .A(n133), .B(n1315), .C(n1522), .Y(n839) );
  NAND2X1 U1241 ( .A(\mem<20><13> ), .B(n1245), .Y(n1523) );
  OAI21X1 U1242 ( .A(n133), .B(n1316), .C(n1523), .Y(n840) );
  NAND2X1 U1243 ( .A(\mem<20><14> ), .B(n1245), .Y(n1524) );
  OAI21X1 U1244 ( .A(n133), .B(n1317), .C(n1524), .Y(n841) );
  NAND2X1 U1245 ( .A(\mem<20><15> ), .B(n1245), .Y(n1525) );
  OAI21X1 U1246 ( .A(n133), .B(n1318), .C(n1525), .Y(n842) );
  NAND2X1 U1247 ( .A(\mem<19><0> ), .B(n10), .Y(n1526) );
  OAI21X1 U1248 ( .A(n137), .B(n1293), .C(n1526), .Y(n843) );
  NAND2X1 U1249 ( .A(\mem<19><1> ), .B(n10), .Y(n1527) );
  OAI21X1 U1250 ( .A(n137), .B(n1295), .C(n1527), .Y(n844) );
  NAND2X1 U1251 ( .A(\mem<19><2> ), .B(n10), .Y(n1528) );
  OAI21X1 U1252 ( .A(n137), .B(n1297), .C(n1528), .Y(n845) );
  NAND2X1 U1253 ( .A(\mem<19><3> ), .B(n1246), .Y(n1529) );
  OAI21X1 U1254 ( .A(n137), .B(n1299), .C(n1529), .Y(n846) );
  NAND2X1 U1255 ( .A(\mem<19><4> ), .B(n1247), .Y(n1530) );
  OAI21X1 U1256 ( .A(n137), .B(n1301), .C(n1530), .Y(n847) );
  NAND2X1 U1257 ( .A(\mem<19><5> ), .B(n1247), .Y(n1531) );
  OAI21X1 U1258 ( .A(n137), .B(n1303), .C(n1531), .Y(n848) );
  NAND2X1 U1259 ( .A(\mem<19><6> ), .B(n1246), .Y(n1532) );
  OAI21X1 U1260 ( .A(n137), .B(n1305), .C(n1532), .Y(n849) );
  NAND2X1 U1261 ( .A(\mem<19><7> ), .B(n10), .Y(n1533) );
  OAI21X1 U1262 ( .A(n137), .B(n1307), .C(n1533), .Y(n850) );
  NAND2X1 U1263 ( .A(\mem<19><8> ), .B(n1247), .Y(n1534) );
  OAI21X1 U1264 ( .A(n137), .B(n1309), .C(n1534), .Y(n851) );
  NAND2X1 U1265 ( .A(\mem<19><9> ), .B(n1246), .Y(n1535) );
  OAI21X1 U1266 ( .A(n137), .B(n1311), .C(n1535), .Y(n852) );
  NAND2X1 U1267 ( .A(\mem<19><10> ), .B(n10), .Y(n1536) );
  OAI21X1 U1268 ( .A(n137), .B(n1313), .C(n1536), .Y(n853) );
  NAND2X1 U1269 ( .A(\mem<19><11> ), .B(n10), .Y(n1537) );
  OAI21X1 U1270 ( .A(n137), .B(n1314), .C(n1537), .Y(n854) );
  NAND2X1 U1271 ( .A(\mem<19><12> ), .B(n1246), .Y(n1538) );
  OAI21X1 U1272 ( .A(n137), .B(n1315), .C(n1538), .Y(n855) );
  NAND2X1 U1273 ( .A(\mem<19><13> ), .B(n1247), .Y(n1539) );
  OAI21X1 U1274 ( .A(n137), .B(n1316), .C(n1539), .Y(n856) );
  NAND2X1 U1275 ( .A(\mem<19><14> ), .B(n1247), .Y(n1540) );
  OAI21X1 U1276 ( .A(n137), .B(n1317), .C(n1540), .Y(n857) );
  NAND2X1 U1277 ( .A(\mem<19><15> ), .B(n1246), .Y(n1541) );
  OAI21X1 U1278 ( .A(n137), .B(n1318), .C(n1541), .Y(n858) );
  NAND2X1 U1279 ( .A(\mem<18><0> ), .B(n9), .Y(n1542) );
  OAI21X1 U1280 ( .A(n139), .B(n1293), .C(n1542), .Y(n859) );
  NAND2X1 U1281 ( .A(\mem<18><1> ), .B(n9), .Y(n1543) );
  OAI21X1 U1282 ( .A(n139), .B(n1295), .C(n1543), .Y(n860) );
  NAND2X1 U1283 ( .A(\mem<18><2> ), .B(n9), .Y(n1544) );
  OAI21X1 U1284 ( .A(n139), .B(n1297), .C(n1544), .Y(n861) );
  NAND2X1 U1285 ( .A(\mem<18><3> ), .B(n1248), .Y(n1545) );
  OAI21X1 U1286 ( .A(n139), .B(n1299), .C(n1545), .Y(n862) );
  NAND2X1 U1287 ( .A(\mem<18><4> ), .B(n1249), .Y(n1546) );
  OAI21X1 U1288 ( .A(n139), .B(n1301), .C(n1546), .Y(n863) );
  NAND2X1 U1289 ( .A(\mem<18><5> ), .B(n1249), .Y(n1547) );
  OAI21X1 U1290 ( .A(n139), .B(n1303), .C(n1547), .Y(n864) );
  NAND2X1 U1291 ( .A(\mem<18><6> ), .B(n1248), .Y(n1548) );
  OAI21X1 U1292 ( .A(n139), .B(n1305), .C(n1548), .Y(n865) );
  NAND2X1 U1293 ( .A(\mem<18><7> ), .B(n9), .Y(n1549) );
  OAI21X1 U1294 ( .A(n139), .B(n1307), .C(n1549), .Y(n866) );
  NAND2X1 U1295 ( .A(\mem<18><8> ), .B(n1249), .Y(n1550) );
  OAI21X1 U1296 ( .A(n139), .B(n1309), .C(n1550), .Y(n867) );
  NAND2X1 U1297 ( .A(\mem<18><9> ), .B(n1248), .Y(n1551) );
  OAI21X1 U1298 ( .A(n139), .B(n1311), .C(n1551), .Y(n868) );
  NAND2X1 U1299 ( .A(\mem<18><10> ), .B(n9), .Y(n1552) );
  OAI21X1 U1300 ( .A(n139), .B(n1313), .C(n1552), .Y(n869) );
  NAND2X1 U1301 ( .A(\mem<18><11> ), .B(n9), .Y(n1553) );
  OAI21X1 U1302 ( .A(n139), .B(n1314), .C(n1553), .Y(n870) );
  NAND2X1 U1303 ( .A(\mem<18><12> ), .B(n1248), .Y(n1554) );
  OAI21X1 U1304 ( .A(n139), .B(n1315), .C(n1554), .Y(n871) );
  NAND2X1 U1305 ( .A(\mem<18><13> ), .B(n1249), .Y(n1555) );
  OAI21X1 U1306 ( .A(n139), .B(n1316), .C(n1555), .Y(n872) );
  NAND2X1 U1307 ( .A(\mem<18><14> ), .B(n1249), .Y(n1556) );
  OAI21X1 U1308 ( .A(n139), .B(n1317), .C(n1556), .Y(n873) );
  NAND2X1 U1309 ( .A(\mem<18><15> ), .B(n1248), .Y(n1557) );
  OAI21X1 U1310 ( .A(n139), .B(n1318), .C(n1557), .Y(n874) );
  NAND2X1 U1311 ( .A(\mem<17><0> ), .B(n8), .Y(n1558) );
  OAI21X1 U1312 ( .A(n141), .B(n1293), .C(n1558), .Y(n875) );
  NAND2X1 U1313 ( .A(\mem<17><1> ), .B(n8), .Y(n1559) );
  OAI21X1 U1314 ( .A(n141), .B(n1295), .C(n1559), .Y(n876) );
  NAND2X1 U1315 ( .A(\mem<17><2> ), .B(n8), .Y(n1560) );
  OAI21X1 U1316 ( .A(n141), .B(n1297), .C(n1560), .Y(n877) );
  NAND2X1 U1317 ( .A(\mem<17><3> ), .B(n1250), .Y(n1561) );
  OAI21X1 U1318 ( .A(n141), .B(n1299), .C(n1561), .Y(n878) );
  NAND2X1 U1319 ( .A(\mem<17><4> ), .B(n1251), .Y(n1562) );
  OAI21X1 U1320 ( .A(n141), .B(n1301), .C(n1562), .Y(n879) );
  NAND2X1 U1321 ( .A(\mem<17><5> ), .B(n1251), .Y(n1563) );
  OAI21X1 U1322 ( .A(n141), .B(n1303), .C(n1563), .Y(n880) );
  NAND2X1 U1323 ( .A(\mem<17><6> ), .B(n1250), .Y(n1564) );
  OAI21X1 U1324 ( .A(n141), .B(n1305), .C(n1564), .Y(n881) );
  NAND2X1 U1325 ( .A(\mem<17><7> ), .B(n8), .Y(n1565) );
  OAI21X1 U1326 ( .A(n141), .B(n1307), .C(n1565), .Y(n882) );
  NAND2X1 U1327 ( .A(\mem<17><8> ), .B(n1251), .Y(n1566) );
  OAI21X1 U1328 ( .A(n141), .B(n1309), .C(n1566), .Y(n883) );
  NAND2X1 U1329 ( .A(\mem<17><9> ), .B(n1250), .Y(n1567) );
  OAI21X1 U1330 ( .A(n141), .B(n1311), .C(n1567), .Y(n884) );
  NAND2X1 U1331 ( .A(\mem<17><10> ), .B(n8), .Y(n1568) );
  OAI21X1 U1332 ( .A(n141), .B(n1313), .C(n1568), .Y(n885) );
  NAND2X1 U1333 ( .A(\mem<17><11> ), .B(n8), .Y(n1569) );
  OAI21X1 U1334 ( .A(n141), .B(n1314), .C(n1569), .Y(n886) );
  NAND2X1 U1335 ( .A(\mem<17><12> ), .B(n1250), .Y(n1570) );
  OAI21X1 U1336 ( .A(n141), .B(n1315), .C(n1570), .Y(n887) );
  NAND2X1 U1337 ( .A(\mem<17><13> ), .B(n1251), .Y(n1571) );
  OAI21X1 U1338 ( .A(n141), .B(n1316), .C(n1571), .Y(n888) );
  NAND2X1 U1339 ( .A(\mem<17><14> ), .B(n1251), .Y(n1572) );
  OAI21X1 U1340 ( .A(n141), .B(n1317), .C(n1572), .Y(n889) );
  NAND2X1 U1341 ( .A(\mem<17><15> ), .B(n1250), .Y(n1573) );
  OAI21X1 U1342 ( .A(n141), .B(n1318), .C(n1573), .Y(n890) );
  NAND2X1 U1343 ( .A(\mem<16><0> ), .B(n1253), .Y(n1574) );
  OAI21X1 U1344 ( .A(n1252), .B(n1293), .C(n1574), .Y(n891) );
  NAND2X1 U1345 ( .A(\mem<16><1> ), .B(n12), .Y(n1575) );
  OAI21X1 U1346 ( .A(n1252), .B(n1295), .C(n1575), .Y(n892) );
  NAND2X1 U1347 ( .A(\mem<16><2> ), .B(n12), .Y(n1576) );
  OAI21X1 U1348 ( .A(n1252), .B(n1297), .C(n1576), .Y(n893) );
  NAND2X1 U1349 ( .A(\mem<16><3> ), .B(n1254), .Y(n1577) );
  OAI21X1 U1350 ( .A(n1252), .B(n1299), .C(n1577), .Y(n894) );
  NAND2X1 U1351 ( .A(\mem<16><4> ), .B(n1254), .Y(n1578) );
  OAI21X1 U1352 ( .A(n1252), .B(n1301), .C(n1578), .Y(n895) );
  NAND2X1 U1353 ( .A(\mem<16><5> ), .B(n1253), .Y(n1579) );
  OAI21X1 U1354 ( .A(n1252), .B(n1303), .C(n1579), .Y(n896) );
  NAND2X1 U1355 ( .A(\mem<16><6> ), .B(n1253), .Y(n1580) );
  OAI21X1 U1356 ( .A(n1252), .B(n1305), .C(n1580), .Y(n897) );
  NAND2X1 U1357 ( .A(\mem<16><7> ), .B(n12), .Y(n1581) );
  OAI21X1 U1358 ( .A(n1252), .B(n1307), .C(n1581), .Y(n898) );
  NAND2X1 U1359 ( .A(\mem<16><8> ), .B(n1254), .Y(n1582) );
  OAI21X1 U1360 ( .A(n1252), .B(n1309), .C(n1582), .Y(n899) );
  NAND2X1 U1361 ( .A(\mem<16><9> ), .B(n1253), .Y(n1583) );
  OAI21X1 U1362 ( .A(n1252), .B(n1311), .C(n1583), .Y(n900) );
  NAND2X1 U1363 ( .A(\mem<16><10> ), .B(n1253), .Y(n1584) );
  OAI21X1 U1364 ( .A(n1252), .B(n1313), .C(n1584), .Y(n901) );
  NAND2X1 U1365 ( .A(\mem<16><11> ), .B(n12), .Y(n1585) );
  OAI21X1 U1366 ( .A(n1252), .B(n1314), .C(n1585), .Y(n902) );
  NAND2X1 U1367 ( .A(\mem<16><12> ), .B(n12), .Y(n1586) );
  OAI21X1 U1368 ( .A(n1252), .B(n1315), .C(n1586), .Y(n903) );
  NAND2X1 U1369 ( .A(\mem<16><13> ), .B(n1254), .Y(n1587) );
  OAI21X1 U1370 ( .A(n1252), .B(n1316), .C(n1587), .Y(n904) );
  NAND2X1 U1371 ( .A(\mem<16><14> ), .B(n1254), .Y(n1588) );
  OAI21X1 U1372 ( .A(n1252), .B(n1317), .C(n1588), .Y(n905) );
  NAND2X1 U1373 ( .A(\mem<16><15> ), .B(n1253), .Y(n1589) );
  OAI21X1 U1374 ( .A(n1252), .B(n1318), .C(n1589), .Y(n906) );
  NAND3X1 U1375 ( .A(n1324), .B(n214), .C(n1327), .Y(n1590) );
  NAND2X1 U1376 ( .A(\mem<15><0> ), .B(n7), .Y(n1591) );
  OAI21X1 U1377 ( .A(n143), .B(n1293), .C(n1591), .Y(n907) );
  NAND2X1 U1378 ( .A(\mem<15><1> ), .B(n7), .Y(n1592) );
  OAI21X1 U1379 ( .A(n143), .B(n1295), .C(n1592), .Y(n908) );
  NAND2X1 U1380 ( .A(\mem<15><2> ), .B(n7), .Y(n1593) );
  OAI21X1 U1381 ( .A(n143), .B(n1297), .C(n1593), .Y(n909) );
  NAND2X1 U1382 ( .A(\mem<15><3> ), .B(n1255), .Y(n1594) );
  OAI21X1 U1383 ( .A(n143), .B(n1299), .C(n1594), .Y(n910) );
  NAND2X1 U1384 ( .A(\mem<15><4> ), .B(n1256), .Y(n1595) );
  OAI21X1 U1385 ( .A(n143), .B(n1301), .C(n1595), .Y(n911) );
  NAND2X1 U1386 ( .A(\mem<15><5> ), .B(n1256), .Y(n1596) );
  OAI21X1 U1387 ( .A(n143), .B(n1303), .C(n1596), .Y(n912) );
  NAND2X1 U1388 ( .A(\mem<15><6> ), .B(n1255), .Y(n1597) );
  OAI21X1 U1389 ( .A(n143), .B(n1305), .C(n1597), .Y(n913) );
  NAND2X1 U1390 ( .A(\mem<15><7> ), .B(n7), .Y(n1598) );
  OAI21X1 U1391 ( .A(n143), .B(n1307), .C(n1598), .Y(n914) );
  NAND2X1 U1392 ( .A(\mem<15><8> ), .B(n1256), .Y(n1599) );
  OAI21X1 U1393 ( .A(n143), .B(n1309), .C(n1599), .Y(n915) );
  NAND2X1 U1394 ( .A(\mem<15><9> ), .B(n1255), .Y(n1600) );
  OAI21X1 U1395 ( .A(n143), .B(n1311), .C(n1600), .Y(n916) );
  NAND2X1 U1396 ( .A(\mem<15><10> ), .B(n7), .Y(n1601) );
  OAI21X1 U1397 ( .A(n143), .B(n1313), .C(n1601), .Y(n917) );
  NAND2X1 U1398 ( .A(\mem<15><11> ), .B(n7), .Y(n1602) );
  OAI21X1 U1399 ( .A(n143), .B(n1314), .C(n1602), .Y(n918) );
  NAND2X1 U1400 ( .A(\mem<15><12> ), .B(n1255), .Y(n1603) );
  OAI21X1 U1401 ( .A(n143), .B(n1315), .C(n1603), .Y(n919) );
  NAND2X1 U1402 ( .A(\mem<15><13> ), .B(n1256), .Y(n1604) );
  OAI21X1 U1403 ( .A(n143), .B(n1316), .C(n1604), .Y(n920) );
  NAND2X1 U1404 ( .A(\mem<15><14> ), .B(n1256), .Y(n1605) );
  OAI21X1 U1405 ( .A(n143), .B(n1317), .C(n1605), .Y(n921) );
  NAND2X1 U1406 ( .A(\mem<15><15> ), .B(n1255), .Y(n1606) );
  OAI21X1 U1407 ( .A(n143), .B(n1318), .C(n1606), .Y(n922) );
  NAND2X1 U1408 ( .A(\mem<14><0> ), .B(n6), .Y(n1607) );
  OAI21X1 U1409 ( .A(n145), .B(n1293), .C(n1607), .Y(n923) );
  NAND2X1 U1410 ( .A(\mem<14><1> ), .B(n6), .Y(n1608) );
  OAI21X1 U1411 ( .A(n145), .B(n1295), .C(n1608), .Y(n924) );
  NAND2X1 U1412 ( .A(\mem<14><2> ), .B(n6), .Y(n1609) );
  OAI21X1 U1413 ( .A(n145), .B(n1297), .C(n1609), .Y(n925) );
  NAND2X1 U1414 ( .A(\mem<14><3> ), .B(n1257), .Y(n1610) );
  OAI21X1 U1415 ( .A(n145), .B(n1299), .C(n1610), .Y(n926) );
  NAND2X1 U1416 ( .A(\mem<14><4> ), .B(n1258), .Y(n1611) );
  OAI21X1 U1417 ( .A(n145), .B(n1301), .C(n1611), .Y(n927) );
  NAND2X1 U1418 ( .A(\mem<14><5> ), .B(n1258), .Y(n1612) );
  OAI21X1 U1419 ( .A(n145), .B(n1303), .C(n1612), .Y(n928) );
  NAND2X1 U1420 ( .A(\mem<14><6> ), .B(n1257), .Y(n1613) );
  OAI21X1 U1421 ( .A(n145), .B(n1305), .C(n1613), .Y(n929) );
  NAND2X1 U1422 ( .A(\mem<14><7> ), .B(n6), .Y(n1614) );
  OAI21X1 U1423 ( .A(n145), .B(n1307), .C(n1614), .Y(n930) );
  NAND2X1 U1424 ( .A(\mem<14><8> ), .B(n1258), .Y(n1615) );
  OAI21X1 U1425 ( .A(n145), .B(n1309), .C(n1615), .Y(n931) );
  NAND2X1 U1426 ( .A(\mem<14><9> ), .B(n1257), .Y(n1616) );
  OAI21X1 U1427 ( .A(n145), .B(n1311), .C(n1616), .Y(n932) );
  NAND2X1 U1428 ( .A(\mem<14><10> ), .B(n6), .Y(n1617) );
  OAI21X1 U1429 ( .A(n145), .B(n1313), .C(n1617), .Y(n933) );
  NAND2X1 U1430 ( .A(\mem<14><11> ), .B(n6), .Y(n1618) );
  OAI21X1 U1431 ( .A(n145), .B(n1314), .C(n1618), .Y(n934) );
  NAND2X1 U1432 ( .A(\mem<14><12> ), .B(n1257), .Y(n1619) );
  OAI21X1 U1433 ( .A(n145), .B(n1315), .C(n1619), .Y(n935) );
  NAND2X1 U1434 ( .A(\mem<14><13> ), .B(n1258), .Y(n1620) );
  OAI21X1 U1435 ( .A(n145), .B(n1316), .C(n1620), .Y(n936) );
  NAND2X1 U1436 ( .A(\mem<14><14> ), .B(n1258), .Y(n1621) );
  OAI21X1 U1437 ( .A(n145), .B(n1317), .C(n1621), .Y(n937) );
  NAND2X1 U1438 ( .A(\mem<14><15> ), .B(n1257), .Y(n1622) );
  OAI21X1 U1439 ( .A(n145), .B(n1318), .C(n1622), .Y(n938) );
  NAND2X1 U1440 ( .A(\mem<13><0> ), .B(n5), .Y(n1623) );
  OAI21X1 U1441 ( .A(n147), .B(n1293), .C(n1623), .Y(n939) );
  NAND2X1 U1442 ( .A(\mem<13><1> ), .B(n5), .Y(n1624) );
  OAI21X1 U1443 ( .A(n147), .B(n1295), .C(n1624), .Y(n940) );
  NAND2X1 U1444 ( .A(\mem<13><2> ), .B(n5), .Y(n1625) );
  OAI21X1 U1445 ( .A(n147), .B(n1297), .C(n1625), .Y(n941) );
  NAND2X1 U1446 ( .A(\mem<13><3> ), .B(n1259), .Y(n1626) );
  OAI21X1 U1447 ( .A(n147), .B(n1299), .C(n1626), .Y(n942) );
  NAND2X1 U1448 ( .A(\mem<13><4> ), .B(n1260), .Y(n1627) );
  OAI21X1 U1449 ( .A(n147), .B(n1301), .C(n1627), .Y(n943) );
  NAND2X1 U1450 ( .A(\mem<13><5> ), .B(n1260), .Y(n1628) );
  OAI21X1 U1451 ( .A(n147), .B(n1303), .C(n1628), .Y(n944) );
  NAND2X1 U1452 ( .A(\mem<13><6> ), .B(n1259), .Y(n1629) );
  OAI21X1 U1453 ( .A(n147), .B(n1305), .C(n1629), .Y(n945) );
  NAND2X1 U1454 ( .A(\mem<13><7> ), .B(n5), .Y(n1630) );
  OAI21X1 U1455 ( .A(n147), .B(n1307), .C(n1630), .Y(n946) );
  NAND2X1 U1456 ( .A(\mem<13><8> ), .B(n1260), .Y(n1631) );
  OAI21X1 U1457 ( .A(n147), .B(n1309), .C(n1631), .Y(n947) );
  NAND2X1 U1458 ( .A(\mem<13><9> ), .B(n1259), .Y(n1632) );
  OAI21X1 U1459 ( .A(n147), .B(n1311), .C(n1632), .Y(n948) );
  NAND2X1 U1460 ( .A(\mem<13><10> ), .B(n5), .Y(n1633) );
  OAI21X1 U1461 ( .A(n147), .B(n1313), .C(n1633), .Y(n949) );
  NAND2X1 U1462 ( .A(\mem<13><11> ), .B(n5), .Y(n1634) );
  OAI21X1 U1463 ( .A(n147), .B(n1314), .C(n1634), .Y(n950) );
  NAND2X1 U1464 ( .A(\mem<13><12> ), .B(n1259), .Y(n1635) );
  OAI21X1 U1465 ( .A(n147), .B(n1315), .C(n1635), .Y(n951) );
  NAND2X1 U1466 ( .A(\mem<13><13> ), .B(n1260), .Y(n1636) );
  OAI21X1 U1467 ( .A(n147), .B(n1316), .C(n1636), .Y(n952) );
  NAND2X1 U1468 ( .A(\mem<13><14> ), .B(n1260), .Y(n1637) );
  OAI21X1 U1469 ( .A(n147), .B(n1317), .C(n1637), .Y(n953) );
  NAND2X1 U1470 ( .A(\mem<13><15> ), .B(n1259), .Y(n1638) );
  OAI21X1 U1471 ( .A(n147), .B(n1318), .C(n1638), .Y(n954) );
  NAND2X1 U1472 ( .A(\mem<12><0> ), .B(n4), .Y(n1639) );
  OAI21X1 U1473 ( .A(n149), .B(n1293), .C(n1639), .Y(n955) );
  NAND2X1 U1474 ( .A(\mem<12><1> ), .B(n4), .Y(n1640) );
  OAI21X1 U1475 ( .A(n149), .B(n1295), .C(n1640), .Y(n956) );
  NAND2X1 U1476 ( .A(\mem<12><2> ), .B(n4), .Y(n1641) );
  OAI21X1 U1477 ( .A(n149), .B(n1297), .C(n1641), .Y(n957) );
  NAND2X1 U1478 ( .A(\mem<12><3> ), .B(n1261), .Y(n1642) );
  OAI21X1 U1479 ( .A(n149), .B(n1299), .C(n1642), .Y(n958) );
  NAND2X1 U1480 ( .A(\mem<12><4> ), .B(n1262), .Y(n1643) );
  OAI21X1 U1481 ( .A(n149), .B(n1301), .C(n1643), .Y(n959) );
  NAND2X1 U1482 ( .A(\mem<12><5> ), .B(n1262), .Y(n1644) );
  OAI21X1 U1483 ( .A(n149), .B(n1303), .C(n1644), .Y(n960) );
  NAND2X1 U1484 ( .A(\mem<12><6> ), .B(n1261), .Y(n1645) );
  OAI21X1 U1485 ( .A(n149), .B(n1305), .C(n1645), .Y(n961) );
  NAND2X1 U1486 ( .A(\mem<12><7> ), .B(n4), .Y(n1646) );
  OAI21X1 U1487 ( .A(n149), .B(n1307), .C(n1646), .Y(n962) );
  NAND2X1 U1488 ( .A(\mem<12><8> ), .B(n1262), .Y(n1647) );
  OAI21X1 U1489 ( .A(n149), .B(n1309), .C(n1647), .Y(n963) );
  NAND2X1 U1490 ( .A(\mem<12><9> ), .B(n1261), .Y(n1648) );
  OAI21X1 U1491 ( .A(n149), .B(n1311), .C(n1648), .Y(n964) );
  NAND2X1 U1492 ( .A(\mem<12><10> ), .B(n4), .Y(n1649) );
  OAI21X1 U1493 ( .A(n149), .B(n1313), .C(n1649), .Y(n965) );
  NAND2X1 U1494 ( .A(\mem<12><11> ), .B(n4), .Y(n1650) );
  OAI21X1 U1495 ( .A(n149), .B(n1314), .C(n1650), .Y(n966) );
  NAND2X1 U1496 ( .A(\mem<12><12> ), .B(n1261), .Y(n1651) );
  OAI21X1 U1497 ( .A(n149), .B(n1315), .C(n1651), .Y(n967) );
  NAND2X1 U1498 ( .A(\mem<12><13> ), .B(n1262), .Y(n1652) );
  OAI21X1 U1499 ( .A(n149), .B(n1316), .C(n1652), .Y(n968) );
  NAND2X1 U1500 ( .A(\mem<12><14> ), .B(n1262), .Y(n1653) );
  OAI21X1 U1501 ( .A(n149), .B(n1317), .C(n1653), .Y(n969) );
  NAND2X1 U1502 ( .A(\mem<12><15> ), .B(n1261), .Y(n1654) );
  OAI21X1 U1503 ( .A(n149), .B(n1318), .C(n1654), .Y(n970) );
  NAND2X1 U1504 ( .A(\mem<11><0> ), .B(n3), .Y(n1655) );
  OAI21X1 U1505 ( .A(n151), .B(n1293), .C(n1655), .Y(n971) );
  NAND2X1 U1506 ( .A(\mem<11><1> ), .B(n3), .Y(n1656) );
  OAI21X1 U1507 ( .A(n151), .B(n1294), .C(n1656), .Y(n972) );
  NAND2X1 U1508 ( .A(\mem<11><2> ), .B(n3), .Y(n1657) );
  OAI21X1 U1509 ( .A(n151), .B(n1296), .C(n1657), .Y(n973) );
  NAND2X1 U1510 ( .A(\mem<11><3> ), .B(n1263), .Y(n1658) );
  OAI21X1 U1511 ( .A(n151), .B(n1298), .C(n1658), .Y(n974) );
  NAND2X1 U1512 ( .A(\mem<11><4> ), .B(n1264), .Y(n1659) );
  OAI21X1 U1513 ( .A(n151), .B(n1300), .C(n1659), .Y(n975) );
  NAND2X1 U1514 ( .A(\mem<11><5> ), .B(n1264), .Y(n1660) );
  OAI21X1 U1515 ( .A(n151), .B(n1302), .C(n1660), .Y(n976) );
  NAND2X1 U1516 ( .A(\mem<11><6> ), .B(n1263), .Y(n1661) );
  OAI21X1 U1517 ( .A(n151), .B(n1304), .C(n1661), .Y(n977) );
  NAND2X1 U1518 ( .A(\mem<11><7> ), .B(n3), .Y(n1662) );
  OAI21X1 U1519 ( .A(n151), .B(n1306), .C(n1662), .Y(n978) );
  NAND2X1 U1520 ( .A(\mem<11><8> ), .B(n1264), .Y(n1663) );
  OAI21X1 U1521 ( .A(n151), .B(n1308), .C(n1663), .Y(n979) );
  NAND2X1 U1522 ( .A(\mem<11><9> ), .B(n1263), .Y(n1664) );
  OAI21X1 U1523 ( .A(n151), .B(n1310), .C(n1664), .Y(n980) );
  NAND2X1 U1524 ( .A(\mem<11><10> ), .B(n3), .Y(n1665) );
  OAI21X1 U1525 ( .A(n151), .B(n1312), .C(n1665), .Y(n981) );
  NAND2X1 U1526 ( .A(\mem<11><11> ), .B(n3), .Y(n1666) );
  OAI21X1 U1527 ( .A(n151), .B(n1314), .C(n1666), .Y(n982) );
  NAND2X1 U1528 ( .A(\mem<11><12> ), .B(n1263), .Y(n1667) );
  OAI21X1 U1529 ( .A(n151), .B(n1315), .C(n1667), .Y(n983) );
  NAND2X1 U1530 ( .A(\mem<11><13> ), .B(n1264), .Y(n1668) );
  OAI21X1 U1531 ( .A(n151), .B(n1316), .C(n1668), .Y(n984) );
  NAND2X1 U1532 ( .A(\mem<11><14> ), .B(n1264), .Y(n1669) );
  OAI21X1 U1533 ( .A(n151), .B(n1317), .C(n1669), .Y(n985) );
  NAND2X1 U1534 ( .A(\mem<11><15> ), .B(n1263), .Y(n1670) );
  OAI21X1 U1535 ( .A(n151), .B(n1318), .C(n1670), .Y(n986) );
  NAND2X1 U1536 ( .A(\mem<10><0> ), .B(n2), .Y(n1671) );
  OAI21X1 U1537 ( .A(n153), .B(n1293), .C(n1671), .Y(n987) );
  NAND2X1 U1538 ( .A(\mem<10><1> ), .B(n2), .Y(n1672) );
  OAI21X1 U1539 ( .A(n153), .B(n1294), .C(n1672), .Y(n988) );
  NAND2X1 U1540 ( .A(\mem<10><2> ), .B(n2), .Y(n1673) );
  OAI21X1 U1541 ( .A(n153), .B(n1296), .C(n1673), .Y(n989) );
  NAND2X1 U1542 ( .A(\mem<10><3> ), .B(n1265), .Y(n1674) );
  OAI21X1 U1543 ( .A(n153), .B(n1298), .C(n1674), .Y(n990) );
  NAND2X1 U1544 ( .A(\mem<10><4> ), .B(n1266), .Y(n1675) );
  OAI21X1 U1545 ( .A(n153), .B(n1300), .C(n1675), .Y(n991) );
  NAND2X1 U1546 ( .A(\mem<10><5> ), .B(n1266), .Y(n1676) );
  OAI21X1 U1547 ( .A(n153), .B(n1302), .C(n1676), .Y(n992) );
  NAND2X1 U1548 ( .A(\mem<10><6> ), .B(n1265), .Y(n1677) );
  OAI21X1 U1549 ( .A(n153), .B(n1304), .C(n1677), .Y(n993) );
  NAND2X1 U1550 ( .A(\mem<10><7> ), .B(n2), .Y(n1678) );
  OAI21X1 U1551 ( .A(n153), .B(n1306), .C(n1678), .Y(n994) );
  NAND2X1 U1552 ( .A(\mem<10><8> ), .B(n1266), .Y(n1679) );
  OAI21X1 U1553 ( .A(n153), .B(n1308), .C(n1679), .Y(n995) );
  NAND2X1 U1554 ( .A(\mem<10><9> ), .B(n1265), .Y(n1680) );
  OAI21X1 U1555 ( .A(n153), .B(n1310), .C(n1680), .Y(n996) );
  NAND2X1 U1556 ( .A(\mem<10><10> ), .B(n2), .Y(n1681) );
  OAI21X1 U1557 ( .A(n153), .B(n1312), .C(n1681), .Y(n997) );
  NAND2X1 U1558 ( .A(\mem<10><11> ), .B(n2), .Y(n1682) );
  OAI21X1 U1559 ( .A(n153), .B(n1314), .C(n1682), .Y(n998) );
  NAND2X1 U1560 ( .A(\mem<10><12> ), .B(n1265), .Y(n1683) );
  OAI21X1 U1561 ( .A(n153), .B(n1315), .C(n1683), .Y(n999) );
  NAND2X1 U1562 ( .A(\mem<10><13> ), .B(n1266), .Y(n1684) );
  OAI21X1 U1563 ( .A(n153), .B(n1316), .C(n1684), .Y(n1000) );
  NAND2X1 U1564 ( .A(\mem<10><14> ), .B(n1266), .Y(n1685) );
  OAI21X1 U1565 ( .A(n153), .B(n1317), .C(n1685), .Y(n1001) );
  NAND2X1 U1566 ( .A(\mem<10><15> ), .B(n1265), .Y(n1686) );
  OAI21X1 U1567 ( .A(n153), .B(n1318), .C(n1686), .Y(n1002) );
  NAND2X1 U1568 ( .A(\mem<9><0> ), .B(n1267), .Y(n1687) );
  OAI21X1 U1569 ( .A(n155), .B(n1293), .C(n1687), .Y(n1003) );
  NAND2X1 U1570 ( .A(\mem<9><1> ), .B(n1267), .Y(n1688) );
  OAI21X1 U1571 ( .A(n155), .B(n1294), .C(n1688), .Y(n1004) );
  NAND2X1 U1572 ( .A(\mem<9><2> ), .B(n1268), .Y(n1689) );
  OAI21X1 U1573 ( .A(n155), .B(n1296), .C(n1689), .Y(n1005) );
  NAND2X1 U1574 ( .A(\mem<9><3> ), .B(n1), .Y(n1690) );
  OAI21X1 U1575 ( .A(n155), .B(n1298), .C(n1690), .Y(n1006) );
  NAND2X1 U1576 ( .A(\mem<9><4> ), .B(n1268), .Y(n1691) );
  OAI21X1 U1577 ( .A(n155), .B(n1300), .C(n1691), .Y(n1007) );
  NAND2X1 U1578 ( .A(\mem<9><5> ), .B(n1267), .Y(n1692) );
  OAI21X1 U1579 ( .A(n155), .B(n1302), .C(n1692), .Y(n1008) );
  NAND2X1 U1580 ( .A(\mem<9><6> ), .B(n1), .Y(n1693) );
  OAI21X1 U1581 ( .A(n155), .B(n1304), .C(n1693), .Y(n1009) );
  NAND2X1 U1582 ( .A(\mem<9><7> ), .B(n1267), .Y(n1694) );
  OAI21X1 U1583 ( .A(n155), .B(n1306), .C(n1694), .Y(n1010) );
  NAND2X1 U1584 ( .A(\mem<9><8> ), .B(n1), .Y(n1695) );
  OAI21X1 U1585 ( .A(n155), .B(n1308), .C(n1695), .Y(n1011) );
  NAND2X1 U1586 ( .A(\mem<9><9> ), .B(n1268), .Y(n1696) );
  OAI21X1 U1587 ( .A(n155), .B(n1310), .C(n1696), .Y(n1012) );
  NAND2X1 U1588 ( .A(\mem<9><10> ), .B(n1267), .Y(n1697) );
  OAI21X1 U1589 ( .A(n155), .B(n1312), .C(n1697), .Y(n1013) );
  NAND2X1 U1590 ( .A(\mem<9><11> ), .B(n1), .Y(n1698) );
  OAI21X1 U1591 ( .A(n155), .B(n1314), .C(n1698), .Y(n1014) );
  NAND2X1 U1592 ( .A(\mem<9><12> ), .B(n1), .Y(n1699) );
  OAI21X1 U1593 ( .A(n155), .B(n1315), .C(n1699), .Y(n1015) );
  NAND2X1 U1594 ( .A(\mem<9><13> ), .B(n1267), .Y(n1700) );
  OAI21X1 U1595 ( .A(n155), .B(n1316), .C(n1700), .Y(n1016) );
  NAND2X1 U1596 ( .A(\mem<9><14> ), .B(n1268), .Y(n1701) );
  OAI21X1 U1597 ( .A(n155), .B(n1317), .C(n1701), .Y(n1017) );
  NAND2X1 U1598 ( .A(\mem<9><15> ), .B(n1268), .Y(n1702) );
  OAI21X1 U1599 ( .A(n155), .B(n1318), .C(n1702), .Y(n1018) );
  NAND2X1 U1600 ( .A(\mem<8><0> ), .B(n1270), .Y(n1704) );
  OAI21X1 U1601 ( .A(n1269), .B(n1293), .C(n1704), .Y(n1019) );
  NAND2X1 U1602 ( .A(\mem<8><1> ), .B(n1270), .Y(n1705) );
  OAI21X1 U1603 ( .A(n1269), .B(n1294), .C(n1705), .Y(n1020) );
  NAND2X1 U1604 ( .A(\mem<8><2> ), .B(n1270), .Y(n1706) );
  OAI21X1 U1605 ( .A(n1269), .B(n1296), .C(n1706), .Y(n1021) );
  NAND2X1 U1606 ( .A(\mem<8><3> ), .B(n1270), .Y(n1707) );
  OAI21X1 U1607 ( .A(n1269), .B(n1298), .C(n1707), .Y(n1022) );
  NAND2X1 U1608 ( .A(\mem<8><4> ), .B(n1270), .Y(n1708) );
  OAI21X1 U1609 ( .A(n1269), .B(n1300), .C(n1708), .Y(n1023) );
  NAND2X1 U1610 ( .A(\mem<8><5> ), .B(n1270), .Y(n1709) );
  OAI21X1 U1611 ( .A(n1269), .B(n1302), .C(n1709), .Y(n1024) );
  NAND2X1 U1612 ( .A(\mem<8><6> ), .B(n1270), .Y(n1710) );
  OAI21X1 U1613 ( .A(n1269), .B(n1304), .C(n1710), .Y(n1025) );
  NAND2X1 U1614 ( .A(\mem<8><7> ), .B(n1270), .Y(n1711) );
  OAI21X1 U1615 ( .A(n1269), .B(n1306), .C(n1711), .Y(n1026) );
  NAND2X1 U1616 ( .A(\mem<8><8> ), .B(n1271), .Y(n1712) );
  OAI21X1 U1617 ( .A(n1269), .B(n1308), .C(n1712), .Y(n1027) );
  NAND2X1 U1618 ( .A(\mem<8><9> ), .B(n1271), .Y(n1713) );
  OAI21X1 U1619 ( .A(n1269), .B(n1310), .C(n1713), .Y(n1028) );
  NAND2X1 U1620 ( .A(\mem<8><10> ), .B(n1271), .Y(n1714) );
  OAI21X1 U1621 ( .A(n1269), .B(n1312), .C(n1714), .Y(n1029) );
  NAND2X1 U1622 ( .A(\mem<8><11> ), .B(n1271), .Y(n1715) );
  OAI21X1 U1623 ( .A(n1269), .B(n1314), .C(n1715), .Y(n1030) );
  NAND2X1 U1624 ( .A(\mem<8><12> ), .B(n1271), .Y(n1716) );
  OAI21X1 U1625 ( .A(n1269), .B(n1315), .C(n1716), .Y(n1031) );
  NAND2X1 U1626 ( .A(\mem<8><13> ), .B(n1271), .Y(n1717) );
  OAI21X1 U1627 ( .A(n1269), .B(n1316), .C(n1717), .Y(n1032) );
  NAND2X1 U1628 ( .A(\mem<8><14> ), .B(n1271), .Y(n1718) );
  OAI21X1 U1629 ( .A(n1269), .B(n1317), .C(n1718), .Y(n1033) );
  NAND2X1 U1630 ( .A(\mem<8><15> ), .B(n1271), .Y(n1719) );
  OAI21X1 U1631 ( .A(n1269), .B(n1318), .C(n1719), .Y(n1034) );
  NAND3X1 U1632 ( .A(n1325), .B(n214), .C(n1327), .Y(n1720) );
  NAND2X1 U1633 ( .A(\mem<7><0> ), .B(n1272), .Y(n1721) );
  OAI21X1 U1634 ( .A(n157), .B(n1292), .C(n1721), .Y(n1035) );
  NAND2X1 U1635 ( .A(\mem<7><1> ), .B(n1272), .Y(n1722) );
  OAI21X1 U1636 ( .A(n157), .B(n1294), .C(n1722), .Y(n1036) );
  NAND2X1 U1637 ( .A(\mem<7><2> ), .B(n1272), .Y(n1723) );
  OAI21X1 U1638 ( .A(n157), .B(n1296), .C(n1723), .Y(n1037) );
  NAND2X1 U1639 ( .A(\mem<7><3> ), .B(n1272), .Y(n1724) );
  OAI21X1 U1640 ( .A(n157), .B(n1298), .C(n1724), .Y(n1038) );
  NAND2X1 U1641 ( .A(\mem<7><4> ), .B(n1272), .Y(n1725) );
  OAI21X1 U1642 ( .A(n157), .B(n1300), .C(n1725), .Y(n1039) );
  NAND2X1 U1643 ( .A(\mem<7><5> ), .B(n1272), .Y(n1726) );
  OAI21X1 U1644 ( .A(n157), .B(n1302), .C(n1726), .Y(n1040) );
  NAND2X1 U1645 ( .A(\mem<7><6> ), .B(n1272), .Y(n1727) );
  OAI21X1 U1646 ( .A(n157), .B(n1304), .C(n1727), .Y(n1041) );
  NAND2X1 U1647 ( .A(\mem<7><7> ), .B(n1272), .Y(n1728) );
  OAI21X1 U1648 ( .A(n157), .B(n1306), .C(n1728), .Y(n1042) );
  NAND2X1 U1649 ( .A(\mem<7><8> ), .B(n1273), .Y(n1729) );
  OAI21X1 U1650 ( .A(n157), .B(n1308), .C(n1729), .Y(n1043) );
  NAND2X1 U1651 ( .A(\mem<7><9> ), .B(n1273), .Y(n1730) );
  OAI21X1 U1652 ( .A(n157), .B(n1310), .C(n1730), .Y(n1044) );
  NAND2X1 U1653 ( .A(\mem<7><10> ), .B(n1273), .Y(n1731) );
  OAI21X1 U1654 ( .A(n157), .B(n1312), .C(n1731), .Y(n1045) );
  NAND2X1 U1655 ( .A(\mem<7><11> ), .B(n1273), .Y(n1732) );
  OAI21X1 U1656 ( .A(n157), .B(n1314), .C(n1732), .Y(n1046) );
  NAND2X1 U1657 ( .A(\mem<7><12> ), .B(n1273), .Y(n1733) );
  OAI21X1 U1658 ( .A(n157), .B(n1315), .C(n1733), .Y(n1047) );
  NAND2X1 U1659 ( .A(\mem<7><13> ), .B(n1273), .Y(n1734) );
  OAI21X1 U1660 ( .A(n157), .B(n1316), .C(n1734), .Y(n1048) );
  NAND2X1 U1661 ( .A(\mem<7><14> ), .B(n1273), .Y(n1735) );
  OAI21X1 U1662 ( .A(n157), .B(n1317), .C(n1735), .Y(n1049) );
  NAND2X1 U1663 ( .A(\mem<7><15> ), .B(n1273), .Y(n1736) );
  OAI21X1 U1664 ( .A(n157), .B(n1318), .C(n1736), .Y(n1050) );
  NAND2X1 U1665 ( .A(\mem<6><0> ), .B(n1274), .Y(n1737) );
  OAI21X1 U1666 ( .A(n159), .B(n1293), .C(n1737), .Y(n1051) );
  NAND2X1 U1667 ( .A(\mem<6><1> ), .B(n1274), .Y(n1738) );
  OAI21X1 U1668 ( .A(n159), .B(n1294), .C(n1738), .Y(n1052) );
  NAND2X1 U1669 ( .A(\mem<6><2> ), .B(n1274), .Y(n1739) );
  OAI21X1 U1670 ( .A(n159), .B(n1296), .C(n1739), .Y(n1053) );
  NAND2X1 U1671 ( .A(\mem<6><3> ), .B(n1274), .Y(n1740) );
  OAI21X1 U1672 ( .A(n159), .B(n1298), .C(n1740), .Y(n1054) );
  NAND2X1 U1673 ( .A(\mem<6><4> ), .B(n1274), .Y(n1741) );
  OAI21X1 U1674 ( .A(n159), .B(n1300), .C(n1741), .Y(n1055) );
  NAND2X1 U1675 ( .A(\mem<6><5> ), .B(n1274), .Y(n1742) );
  OAI21X1 U1676 ( .A(n159), .B(n1302), .C(n1742), .Y(n1056) );
  NAND2X1 U1677 ( .A(\mem<6><6> ), .B(n1274), .Y(n1743) );
  OAI21X1 U1678 ( .A(n159), .B(n1304), .C(n1743), .Y(n1057) );
  NAND2X1 U1679 ( .A(\mem<6><7> ), .B(n1274), .Y(n1744) );
  OAI21X1 U1680 ( .A(n159), .B(n1306), .C(n1744), .Y(n1058) );
  NAND2X1 U1681 ( .A(\mem<6><8> ), .B(n1275), .Y(n1745) );
  OAI21X1 U1682 ( .A(n159), .B(n1308), .C(n1745), .Y(n1059) );
  NAND2X1 U1683 ( .A(\mem<6><9> ), .B(n1275), .Y(n1746) );
  OAI21X1 U1684 ( .A(n159), .B(n1310), .C(n1746), .Y(n1060) );
  NAND2X1 U1685 ( .A(\mem<6><10> ), .B(n1275), .Y(n1747) );
  OAI21X1 U1686 ( .A(n159), .B(n1312), .C(n1747), .Y(n1061) );
  NAND2X1 U1687 ( .A(\mem<6><11> ), .B(n1275), .Y(n1748) );
  OAI21X1 U1688 ( .A(n159), .B(n1314), .C(n1748), .Y(n1062) );
  NAND2X1 U1689 ( .A(\mem<6><12> ), .B(n1275), .Y(n1749) );
  OAI21X1 U1690 ( .A(n159), .B(n1315), .C(n1749), .Y(n1063) );
  NAND2X1 U1691 ( .A(\mem<6><13> ), .B(n1275), .Y(n1750) );
  OAI21X1 U1692 ( .A(n159), .B(n1316), .C(n1750), .Y(n1064) );
  NAND2X1 U1693 ( .A(\mem<6><14> ), .B(n1275), .Y(n1751) );
  OAI21X1 U1694 ( .A(n159), .B(n1317), .C(n1751), .Y(n1065) );
  NAND2X1 U1695 ( .A(\mem<6><15> ), .B(n1275), .Y(n1752) );
  OAI21X1 U1696 ( .A(n159), .B(n1318), .C(n1752), .Y(n1066) );
  NAND2X1 U1697 ( .A(\mem<5><0> ), .B(n1276), .Y(n1754) );
  OAI21X1 U1698 ( .A(n161), .B(n1292), .C(n1754), .Y(n1067) );
  NAND2X1 U1699 ( .A(\mem<5><1> ), .B(n1276), .Y(n1755) );
  OAI21X1 U1700 ( .A(n161), .B(n1294), .C(n1755), .Y(n1068) );
  NAND2X1 U1701 ( .A(\mem<5><2> ), .B(n1276), .Y(n1756) );
  OAI21X1 U1702 ( .A(n161), .B(n1296), .C(n1756), .Y(n1069) );
  NAND2X1 U1703 ( .A(\mem<5><3> ), .B(n1276), .Y(n1757) );
  OAI21X1 U1704 ( .A(n161), .B(n1298), .C(n1757), .Y(n1070) );
  NAND2X1 U1705 ( .A(\mem<5><4> ), .B(n1276), .Y(n1758) );
  OAI21X1 U1706 ( .A(n161), .B(n1300), .C(n1758), .Y(n1071) );
  NAND2X1 U1707 ( .A(\mem<5><5> ), .B(n1276), .Y(n1759) );
  OAI21X1 U1708 ( .A(n161), .B(n1302), .C(n1759), .Y(n1072) );
  NAND2X1 U1709 ( .A(\mem<5><6> ), .B(n1276), .Y(n1760) );
  OAI21X1 U1710 ( .A(n161), .B(n1304), .C(n1760), .Y(n1073) );
  NAND2X1 U1711 ( .A(\mem<5><7> ), .B(n1276), .Y(n1761) );
  OAI21X1 U1712 ( .A(n161), .B(n1306), .C(n1761), .Y(n1074) );
  NAND2X1 U1713 ( .A(\mem<5><8> ), .B(n1277), .Y(n1762) );
  OAI21X1 U1714 ( .A(n161), .B(n1308), .C(n1762), .Y(n1075) );
  NAND2X1 U1715 ( .A(\mem<5><9> ), .B(n1277), .Y(n1763) );
  OAI21X1 U1716 ( .A(n161), .B(n1310), .C(n1763), .Y(n1076) );
  NAND2X1 U1717 ( .A(\mem<5><10> ), .B(n1277), .Y(n1764) );
  OAI21X1 U1718 ( .A(n161), .B(n1312), .C(n1764), .Y(n1077) );
  NAND2X1 U1719 ( .A(\mem<5><11> ), .B(n1277), .Y(n1765) );
  OAI21X1 U1720 ( .A(n161), .B(n1314), .C(n1765), .Y(n1078) );
  NAND2X1 U1721 ( .A(\mem<5><12> ), .B(n1277), .Y(n1766) );
  OAI21X1 U1722 ( .A(n161), .B(n1315), .C(n1766), .Y(n1079) );
  NAND2X1 U1723 ( .A(\mem<5><13> ), .B(n1277), .Y(n1767) );
  OAI21X1 U1724 ( .A(n161), .B(n1316), .C(n1767), .Y(n1080) );
  NAND2X1 U1725 ( .A(\mem<5><14> ), .B(n1277), .Y(n1768) );
  OAI21X1 U1726 ( .A(n161), .B(n1317), .C(n1768), .Y(n1081) );
  NAND2X1 U1727 ( .A(\mem<5><15> ), .B(n1277), .Y(n1769) );
  OAI21X1 U1728 ( .A(n161), .B(n1318), .C(n1769), .Y(n1082) );
  NAND2X1 U1729 ( .A(\mem<4><0> ), .B(n1278), .Y(n1771) );
  OAI21X1 U1730 ( .A(n163), .B(n1293), .C(n1771), .Y(n1083) );
  NAND2X1 U1731 ( .A(\mem<4><1> ), .B(n1278), .Y(n1772) );
  OAI21X1 U1732 ( .A(n163), .B(n1294), .C(n1772), .Y(n1084) );
  NAND2X1 U1733 ( .A(\mem<4><2> ), .B(n1278), .Y(n1773) );
  OAI21X1 U1734 ( .A(n163), .B(n1296), .C(n1773), .Y(n1085) );
  NAND2X1 U1735 ( .A(\mem<4><3> ), .B(n1278), .Y(n1774) );
  OAI21X1 U1736 ( .A(n163), .B(n1298), .C(n1774), .Y(n1086) );
  NAND2X1 U1737 ( .A(\mem<4><4> ), .B(n1278), .Y(n1775) );
  OAI21X1 U1738 ( .A(n163), .B(n1300), .C(n1775), .Y(n1087) );
  NAND2X1 U1739 ( .A(\mem<4><5> ), .B(n1278), .Y(n1776) );
  OAI21X1 U1740 ( .A(n163), .B(n1302), .C(n1776), .Y(n1088) );
  NAND2X1 U1741 ( .A(\mem<4><6> ), .B(n1278), .Y(n1777) );
  OAI21X1 U1742 ( .A(n163), .B(n1304), .C(n1777), .Y(n1089) );
  NAND2X1 U1743 ( .A(\mem<4><7> ), .B(n1278), .Y(n1778) );
  OAI21X1 U1744 ( .A(n163), .B(n1306), .C(n1778), .Y(n1090) );
  NAND2X1 U1745 ( .A(\mem<4><8> ), .B(n1279), .Y(n1779) );
  OAI21X1 U1746 ( .A(n163), .B(n1308), .C(n1779), .Y(n1091) );
  NAND2X1 U1747 ( .A(\mem<4><9> ), .B(n1279), .Y(n1780) );
  OAI21X1 U1748 ( .A(n163), .B(n1310), .C(n1780), .Y(n1092) );
  NAND2X1 U1749 ( .A(\mem<4><10> ), .B(n1279), .Y(n1781) );
  OAI21X1 U1750 ( .A(n163), .B(n1312), .C(n1781), .Y(n1093) );
  NAND2X1 U1751 ( .A(\mem<4><11> ), .B(n1279), .Y(n1782) );
  OAI21X1 U1752 ( .A(n163), .B(n1314), .C(n1782), .Y(n1094) );
  NAND2X1 U1753 ( .A(\mem<4><12> ), .B(n1279), .Y(n1783) );
  OAI21X1 U1754 ( .A(n163), .B(n1315), .C(n1783), .Y(n1095) );
  NAND2X1 U1755 ( .A(\mem<4><13> ), .B(n1279), .Y(n1784) );
  OAI21X1 U1756 ( .A(n163), .B(n1316), .C(n1784), .Y(n1096) );
  NAND2X1 U1757 ( .A(\mem<4><14> ), .B(n1279), .Y(n1785) );
  OAI21X1 U1758 ( .A(n163), .B(n1317), .C(n1785), .Y(n1097) );
  NAND2X1 U1759 ( .A(\mem<4><15> ), .B(n1279), .Y(n1786) );
  OAI21X1 U1760 ( .A(n163), .B(n1318), .C(n1786), .Y(n1098) );
  NAND2X1 U1761 ( .A(\mem<3><0> ), .B(n1280), .Y(n1788) );
  OAI21X1 U1762 ( .A(n165), .B(n1292), .C(n1788), .Y(n1099) );
  NAND2X1 U1763 ( .A(\mem<3><1> ), .B(n1280), .Y(n1789) );
  OAI21X1 U1764 ( .A(n165), .B(n1294), .C(n1789), .Y(n1100) );
  NAND2X1 U1765 ( .A(\mem<3><2> ), .B(n1280), .Y(n1790) );
  OAI21X1 U1766 ( .A(n165), .B(n1296), .C(n1790), .Y(n1101) );
  NAND2X1 U1767 ( .A(\mem<3><3> ), .B(n1280), .Y(n1791) );
  OAI21X1 U1768 ( .A(n165), .B(n1298), .C(n1791), .Y(n1102) );
  NAND2X1 U1769 ( .A(\mem<3><4> ), .B(n1280), .Y(n1792) );
  OAI21X1 U1770 ( .A(n165), .B(n1300), .C(n1792), .Y(n1103) );
  NAND2X1 U1771 ( .A(\mem<3><5> ), .B(n1280), .Y(n1793) );
  OAI21X1 U1772 ( .A(n165), .B(n1302), .C(n1793), .Y(n1104) );
  NAND2X1 U1773 ( .A(\mem<3><6> ), .B(n1280), .Y(n1794) );
  OAI21X1 U1774 ( .A(n165), .B(n1304), .C(n1794), .Y(n1105) );
  NAND2X1 U1775 ( .A(\mem<3><7> ), .B(n1280), .Y(n1795) );
  OAI21X1 U1776 ( .A(n165), .B(n1306), .C(n1795), .Y(n1106) );
  NAND2X1 U1777 ( .A(\mem<3><8> ), .B(n1281), .Y(n1796) );
  OAI21X1 U1778 ( .A(n165), .B(n1308), .C(n1796), .Y(n1107) );
  NAND2X1 U1779 ( .A(\mem<3><9> ), .B(n1281), .Y(n1797) );
  OAI21X1 U1780 ( .A(n165), .B(n1310), .C(n1797), .Y(n1108) );
  NAND2X1 U1781 ( .A(\mem<3><10> ), .B(n1281), .Y(n1798) );
  OAI21X1 U1782 ( .A(n165), .B(n1312), .C(n1798), .Y(n1109) );
  NAND2X1 U1783 ( .A(\mem<3><11> ), .B(n1281), .Y(n1799) );
  OAI21X1 U1784 ( .A(n165), .B(n1314), .C(n1799), .Y(n1110) );
  NAND2X1 U1785 ( .A(\mem<3><12> ), .B(n1281), .Y(n1800) );
  OAI21X1 U1786 ( .A(n165), .B(n1315), .C(n1800), .Y(n1111) );
  NAND2X1 U1787 ( .A(\mem<3><13> ), .B(n1281), .Y(n1801) );
  OAI21X1 U1788 ( .A(n165), .B(n1316), .C(n1801), .Y(n1112) );
  NAND2X1 U1789 ( .A(\mem<3><14> ), .B(n1281), .Y(n1802) );
  OAI21X1 U1790 ( .A(n165), .B(n1317), .C(n1802), .Y(n1113) );
  NAND2X1 U1791 ( .A(\mem<3><15> ), .B(n1281), .Y(n1803) );
  OAI21X1 U1792 ( .A(n165), .B(n1318), .C(n1803), .Y(n1114) );
  NAND2X1 U1793 ( .A(\mem<2><0> ), .B(n1282), .Y(n1805) );
  OAI21X1 U1794 ( .A(n167), .B(n1293), .C(n1805), .Y(n1115) );
  NAND2X1 U1795 ( .A(\mem<2><1> ), .B(n1282), .Y(n1806) );
  OAI21X1 U1796 ( .A(n167), .B(n1294), .C(n1806), .Y(n1116) );
  NAND2X1 U1797 ( .A(\mem<2><2> ), .B(n1282), .Y(n1807) );
  OAI21X1 U1798 ( .A(n167), .B(n1296), .C(n1807), .Y(n1117) );
  NAND2X1 U1799 ( .A(\mem<2><3> ), .B(n1282), .Y(n1808) );
  OAI21X1 U1800 ( .A(n167), .B(n1298), .C(n1808), .Y(n1118) );
  NAND2X1 U1801 ( .A(\mem<2><4> ), .B(n1282), .Y(n1809) );
  OAI21X1 U1802 ( .A(n167), .B(n1300), .C(n1809), .Y(n1119) );
  NAND2X1 U1803 ( .A(\mem<2><5> ), .B(n1282), .Y(n1810) );
  OAI21X1 U1804 ( .A(n167), .B(n1302), .C(n1810), .Y(n1120) );
  NAND2X1 U1805 ( .A(\mem<2><6> ), .B(n1282), .Y(n1811) );
  OAI21X1 U1806 ( .A(n167), .B(n1304), .C(n1811), .Y(n1121) );
  NAND2X1 U1807 ( .A(\mem<2><7> ), .B(n1282), .Y(n1812) );
  OAI21X1 U1808 ( .A(n167), .B(n1306), .C(n1812), .Y(n1122) );
  NAND2X1 U1809 ( .A(\mem<2><8> ), .B(n1283), .Y(n1813) );
  OAI21X1 U1810 ( .A(n167), .B(n1308), .C(n1813), .Y(n1123) );
  NAND2X1 U1811 ( .A(\mem<2><9> ), .B(n1283), .Y(n1814) );
  OAI21X1 U1812 ( .A(n167), .B(n1310), .C(n1814), .Y(n1124) );
  NAND2X1 U1813 ( .A(\mem<2><10> ), .B(n1283), .Y(n1815) );
  OAI21X1 U1814 ( .A(n167), .B(n1312), .C(n1815), .Y(n1125) );
  NAND2X1 U1815 ( .A(\mem<2><11> ), .B(n1283), .Y(n1816) );
  OAI21X1 U1816 ( .A(n167), .B(n1314), .C(n1816), .Y(n1126) );
  NAND2X1 U1817 ( .A(\mem<2><12> ), .B(n1283), .Y(n1817) );
  OAI21X1 U1818 ( .A(n167), .B(n1315), .C(n1817), .Y(n1127) );
  NAND2X1 U1819 ( .A(\mem<2><13> ), .B(n1283), .Y(n1818) );
  OAI21X1 U1820 ( .A(n167), .B(n1316), .C(n1818), .Y(n1128) );
  NAND2X1 U1821 ( .A(\mem<2><14> ), .B(n1283), .Y(n1819) );
  OAI21X1 U1822 ( .A(n167), .B(n1317), .C(n1819), .Y(n1129) );
  NAND2X1 U1823 ( .A(\mem<2><15> ), .B(n1283), .Y(n1820) );
  OAI21X1 U1824 ( .A(n167), .B(n1318), .C(n1820), .Y(n1130) );
  NAND2X1 U1825 ( .A(\mem<1><0> ), .B(n1284), .Y(n1822) );
  OAI21X1 U1826 ( .A(n169), .B(n1292), .C(n1822), .Y(n1131) );
  NAND2X1 U1827 ( .A(\mem<1><1> ), .B(n1284), .Y(n1823) );
  OAI21X1 U1828 ( .A(n169), .B(n1294), .C(n1823), .Y(n1132) );
  NAND2X1 U1829 ( .A(\mem<1><2> ), .B(n1284), .Y(n1824) );
  OAI21X1 U1830 ( .A(n169), .B(n1296), .C(n1824), .Y(n1133) );
  NAND2X1 U1831 ( .A(\mem<1><3> ), .B(n1284), .Y(n1825) );
  OAI21X1 U1832 ( .A(n169), .B(n1298), .C(n1825), .Y(n1134) );
  NAND2X1 U1833 ( .A(\mem<1><4> ), .B(n1284), .Y(n1826) );
  OAI21X1 U1834 ( .A(n169), .B(n1300), .C(n1826), .Y(n1135) );
  NAND2X1 U1835 ( .A(\mem<1><5> ), .B(n1284), .Y(n1827) );
  OAI21X1 U1836 ( .A(n169), .B(n1302), .C(n1827), .Y(n1136) );
  NAND2X1 U1837 ( .A(\mem<1><6> ), .B(n1284), .Y(n1828) );
  OAI21X1 U1838 ( .A(n169), .B(n1304), .C(n1828), .Y(n1137) );
  NAND2X1 U1839 ( .A(\mem<1><7> ), .B(n1284), .Y(n1829) );
  OAI21X1 U1840 ( .A(n169), .B(n1306), .C(n1829), .Y(n1138) );
  NAND2X1 U1841 ( .A(\mem<1><8> ), .B(n1285), .Y(n1830) );
  OAI21X1 U1842 ( .A(n169), .B(n1308), .C(n1830), .Y(n1139) );
  NAND2X1 U1843 ( .A(\mem<1><9> ), .B(n1285), .Y(n1831) );
  OAI21X1 U1844 ( .A(n169), .B(n1310), .C(n1831), .Y(n1140) );
  NAND2X1 U1845 ( .A(\mem<1><10> ), .B(n1285), .Y(n1832) );
  OAI21X1 U1846 ( .A(n169), .B(n1312), .C(n1832), .Y(n1141) );
  NAND2X1 U1847 ( .A(\mem<1><11> ), .B(n1285), .Y(n1833) );
  OAI21X1 U1848 ( .A(n169), .B(n1314), .C(n1833), .Y(n1142) );
  NAND2X1 U1849 ( .A(\mem<1><12> ), .B(n1285), .Y(n1834) );
  OAI21X1 U1850 ( .A(n169), .B(n1315), .C(n1834), .Y(n1143) );
  NAND2X1 U1851 ( .A(\mem<1><13> ), .B(n1285), .Y(n1835) );
  OAI21X1 U1852 ( .A(n169), .B(n1316), .C(n1835), .Y(n1144) );
  NAND2X1 U1853 ( .A(\mem<1><14> ), .B(n1285), .Y(n1836) );
  OAI21X1 U1854 ( .A(n169), .B(n1317), .C(n1836), .Y(n1145) );
  NAND2X1 U1855 ( .A(\mem<1><15> ), .B(n1285), .Y(n1837) );
  OAI21X1 U1856 ( .A(n169), .B(n1318), .C(n1837), .Y(n1146) );
  NAND2X1 U1857 ( .A(\mem<0><0> ), .B(n1287), .Y(n1840) );
  OAI21X1 U1858 ( .A(n1286), .B(n1293), .C(n1840), .Y(n1147) );
  NAND2X1 U1859 ( .A(\mem<0><1> ), .B(n11), .Y(n1841) );
  OAI21X1 U1860 ( .A(n1286), .B(n1294), .C(n1841), .Y(n1148) );
  NAND2X1 U1861 ( .A(\mem<0><2> ), .B(n11), .Y(n1842) );
  OAI21X1 U1862 ( .A(n1286), .B(n1296), .C(n1842), .Y(n1149) );
  NAND2X1 U1863 ( .A(\mem<0><3> ), .B(n1288), .Y(n1843) );
  OAI21X1 U1864 ( .A(n1286), .B(n1298), .C(n1843), .Y(n1150) );
  NAND2X1 U1865 ( .A(\mem<0><4> ), .B(n1288), .Y(n1844) );
  OAI21X1 U1866 ( .A(n1286), .B(n1300), .C(n1844), .Y(n1151) );
  NAND2X1 U1867 ( .A(\mem<0><5> ), .B(n1287), .Y(n1845) );
  OAI21X1 U1868 ( .A(n1286), .B(n1302), .C(n1845), .Y(n1152) );
  NAND2X1 U1869 ( .A(\mem<0><6> ), .B(n1287), .Y(n1846) );
  OAI21X1 U1870 ( .A(n1286), .B(n1304), .C(n1846), .Y(n1153) );
  NAND2X1 U1871 ( .A(\mem<0><7> ), .B(n11), .Y(n1847) );
  OAI21X1 U1872 ( .A(n1286), .B(n1306), .C(n1847), .Y(n1154) );
  NAND2X1 U1873 ( .A(\mem<0><8> ), .B(n1288), .Y(n1848) );
  OAI21X1 U1874 ( .A(n1286), .B(n1308), .C(n1848), .Y(n1155) );
  NAND2X1 U1875 ( .A(\mem<0><9> ), .B(n1287), .Y(n1849) );
  OAI21X1 U1876 ( .A(n1286), .B(n1310), .C(n1849), .Y(n1156) );
  NAND2X1 U1877 ( .A(\mem<0><10> ), .B(n1287), .Y(n1850) );
  OAI21X1 U1878 ( .A(n1286), .B(n1312), .C(n1850), .Y(n1157) );
  NAND2X1 U1879 ( .A(\mem<0><11> ), .B(n11), .Y(n1851) );
  OAI21X1 U1880 ( .A(n1286), .B(n1314), .C(n1851), .Y(n1158) );
  NAND2X1 U1881 ( .A(\mem<0><12> ), .B(n11), .Y(n1852) );
  OAI21X1 U1882 ( .A(n1286), .B(n1315), .C(n1852), .Y(n1159) );
  NAND2X1 U1883 ( .A(\mem<0><13> ), .B(n1288), .Y(n1853) );
  OAI21X1 U1884 ( .A(n1286), .B(n1316), .C(n1853), .Y(n1160) );
  NAND2X1 U1885 ( .A(\mem<0><14> ), .B(n1288), .Y(n1854) );
  OAI21X1 U1886 ( .A(n1286), .B(n1317), .C(n1854), .Y(n1161) );
  NAND2X1 U1887 ( .A(\mem<0><15> ), .B(n1287), .Y(n1855) );
  OAI21X1 U1888 ( .A(n1286), .B(n1318), .C(n1855), .Y(n1162) );
endmodule


module memc_Size16_6 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N19, N31, net59006, net59340, net59460, net59458,
         net59640, net59638, net60096, net60094, net60828, net60826, net65995,
         \C2334/net60892 , \C2334/net60452 , \C2334/net60460 ,
         \C2334/net60462 , \C2334/net60464 , \C2334/net60466 ,
         \C2334/net60468 , \C2334/net60470 , \C2334/net60472 ,
         \C2334/net60474 , \C2334/net60476 , \C2334/net60478 ,
         \C2334/net60484 , \C2334/net60490 , \C2334/net60496 ,
         \C2334/net60504 , \C2334/net60506 , \C2334/net60160 ,
         \C2334/net59908 , \C2334/net59910 , \C2334/net59912 ,
         \C2334/net59914 , \C2334/net59916 , \C2334/net59918 ,
         \C2334/net59920 , \C2334/net59922 , \C2334/net59924 ,
         \C2334/net59926 , \C2334/net59928 , \C2334/net59930 ,
         \C2334/net59934 , \C2334/net59710 , \C2334/net59712 ,
         \C2334/net59716 , \C2334/net59718 , \C2334/net59722 ,
         \C2334/net59512 , \C2334/net59514 , \C2334/net59380 ,
         \C2334/net11884 , net80056, net100591, net100598, net101601,
         net101600, net104291, net100597, \C2334/net11880 , net104441,
         net100612, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n36, n37, n40, n41, n43, n45, n48,
         n52, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n80, n82,
         n99, n101, n118, n120, n137, n139, n156, n158, n175, n177, n194, n196,
         n215, n217, n233, n235, n251, n253, n269, n271, n287, n289, n305,
         n307, n323, n325, n341, n343, n360, n362, n378, n380, n396, n398,
         n414, n416, n432, n434, n450, n452, n468, n470, n486, n488, n505,
         n507, n523, n525, n541, n543, n559, n561, n577, n579, n595, n597,
         n613, n615, n631, n633, n650, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;
  assign \data_out<6>  = net80056;
  assign \data_out<4>  = net100598;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1810), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1811), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1812), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1813), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1814), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1815), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1816), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1817), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1818), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1819), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1820), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1821), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1822), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1823), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1824), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1825), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1826), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1827), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1828), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1829), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1830), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1831), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1832), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1833), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1834), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1835), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1836), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1837), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1838), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1839), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1840), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1841), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1842), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1843), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1844), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1845), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1846), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1847), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1848), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1849), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1850), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1851), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1852), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1853), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1854), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1855), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1856), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1857), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1858), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1859), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1860), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1861), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1862), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1863), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1864), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1865), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1866), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1867), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1868), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1869), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1870), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1871), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1872), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1873), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1874), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1875), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1876), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1877), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1878), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1879), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1880), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1881), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1882), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1883), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1884), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1885), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1886), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1887), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1888), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1889), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1890), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1891), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1892), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1893), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1894), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1895), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1896), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1897), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1898), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1899), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1900), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1901), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1902), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1903), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1904), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1905), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1906), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1907), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1908), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1909), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1910), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1911), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1912), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1913), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1914), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1915), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1916), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1917), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1918), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1919), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1920), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1921), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1922), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1923), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1924), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1925), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1926), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1927), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1928), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1929), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1930), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1931), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1932), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1933), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1934), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1935), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1936), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1937), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1938), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1939), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1940), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1941), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1942), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1943), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1944), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1945), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1946), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1947), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1948), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1949), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1950), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1951), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1952), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1953), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1954), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1955), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1956), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1957), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1958), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1959), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1960), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1961), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1962), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1963), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1964), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1965), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1966), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1967), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1968), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1969), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1970), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1971), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1972), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n1973), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n1974), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n1975), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n1976), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n1977), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1978), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1979), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1980), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1981), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1982), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1983), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1984), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1985), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n1986), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n1987), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n1988), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n1989), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n1990), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n1991), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n1992), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n1993), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1994), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1995), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1996), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1997), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1998), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1999), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2000), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2001), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2002), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2003), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2004), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2005), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2006), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2007), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2008), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2009), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2010), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2011), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2012), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2013), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2014), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2015), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2016), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2017), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2018), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2019), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2020), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2021), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2022), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2023), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2024), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2025), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2026), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2027), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2028), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2029), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2030), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2031), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2032), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2033), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2034), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2035), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2036), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2037), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2038), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2039), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2040), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2041), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2042), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2043), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2044), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2045), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2046), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2047), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2048), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2049), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2050), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2051), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2052), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2053), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2054), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2055), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2056), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2057), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2058), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2059), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2060), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2061), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2062), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2063), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2064), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2065), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2066), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2067), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2068), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2069), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2070), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2071), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2072), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2073), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2074), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2075), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2076), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2077), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2078), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2079), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2080), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2081), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2082), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2083), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2084), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2085), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2086), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2087), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2088), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2089), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2090), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2091), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2092), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2093), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2094), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2095), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2096), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2097), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2098), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2099), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2100), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2101), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2102), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2103), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2104), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2105), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2106), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2107), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2108), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2109), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2110), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2111), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2112), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2113), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2114), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2115), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2116), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2117), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2118), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2119), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2120), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2121), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2122), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2123), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2124), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2125), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2126), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2127), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2128), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2129), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2130), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2131), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2132), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2133), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2134), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2135), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2136), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2137), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2138), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2139), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2140), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2141), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2142), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2143), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2144), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2145), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2146), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2147), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2148), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2149), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2150), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2151), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2152), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2153), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2154), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2155), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2156), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2157), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2158), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2159), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2160), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2161), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2162), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2163), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2164), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2165), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2166), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2167), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2168), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2169), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2170), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2171), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2172), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2173), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2174), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2175), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2176), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2177), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2178), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2179), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2180), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2181), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2182), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2183), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2184), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2185), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2186), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2187), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2188), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2189), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2190), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2191), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2192), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2193), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2194), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2195), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2196), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2197), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2198), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2199), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2200), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2201), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2202), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2203), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2204), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2205), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2206), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2207), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2208), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2209), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2210), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2211), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2212), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2213), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2214), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2215), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2216), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2217), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2218), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2219), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2220), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2221), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2222), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2223), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2224), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2225), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2226), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2227), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2228), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2229), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2230), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2231), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2232), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2233), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2234), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2235), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2236), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2237), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2238), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2239), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2240), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2241), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2242), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2243), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2244), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2245), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2246), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2247), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2248), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2249), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2250), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2251), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2252), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2253), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2254), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2255), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2256), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2257), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2258), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2259), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2260), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2261), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2262), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2263), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2264), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2265), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2266), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2267), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2268), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2269), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2270), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2271), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2272), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2273), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2274), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2275), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2276), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2277), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2278), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2279), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2280), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2281), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2282), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2283), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2284), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2285), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2286), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2287), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2288), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2289), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2290), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2291), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2292), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2293), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2294), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2295), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2296), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2297), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2298), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2299), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2300), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2301), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2302), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2303), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2304), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2305), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2306), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2307), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2308), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2309), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2310), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2311), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2312), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2313), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2314), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2315), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2316), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2317), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2318), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2319), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2320), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2321), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(net65995), .B(net59006), .Y(n2831) );
  OAI21X1 U61 ( .A(n1773), .B(n1804), .C(n2847), .Y(n2321) );
  NAND2X1 U62 ( .A(\mem<31><0> ), .B(n1775), .Y(n2847) );
  OAI21X1 U63 ( .A(n1773), .B(n1802), .C(n2846), .Y(n2320) );
  NAND2X1 U64 ( .A(\mem<31><1> ), .B(n1775), .Y(n2846) );
  OAI21X1 U65 ( .A(n1773), .B(n1800), .C(n2845), .Y(n2319) );
  NAND2X1 U66 ( .A(\mem<31><2> ), .B(n1775), .Y(n2845) );
  OAI21X1 U67 ( .A(n1773), .B(n1798), .C(n2844), .Y(n2318) );
  NAND2X1 U68 ( .A(\mem<31><3> ), .B(n1775), .Y(n2844) );
  OAI21X1 U69 ( .A(n1773), .B(n1796), .C(n2843), .Y(n2317) );
  NAND2X1 U70 ( .A(\mem<31><4> ), .B(n1775), .Y(n2843) );
  OAI21X1 U71 ( .A(n1773), .B(n1794), .C(n2842), .Y(n2316) );
  NAND2X1 U72 ( .A(\mem<31><5> ), .B(n1775), .Y(n2842) );
  OAI21X1 U73 ( .A(n1773), .B(n1792), .C(n2841), .Y(n2315) );
  NAND2X1 U74 ( .A(\mem<31><6> ), .B(n1775), .Y(n2841) );
  OAI21X1 U75 ( .A(n1773), .B(n1790), .C(n2840), .Y(n2314) );
  NAND2X1 U76 ( .A(\mem<31><7> ), .B(n1775), .Y(n2840) );
  OAI21X1 U77 ( .A(n1773), .B(n1789), .C(n2839), .Y(n2313) );
  NAND2X1 U78 ( .A(\mem<31><8> ), .B(n1774), .Y(n2839) );
  OAI21X1 U79 ( .A(n1773), .B(n1788), .C(n2838), .Y(n2312) );
  NAND2X1 U80 ( .A(\mem<31><9> ), .B(n1774), .Y(n2838) );
  OAI21X1 U81 ( .A(n1773), .B(n1786), .C(n2837), .Y(n2311) );
  NAND2X1 U82 ( .A(\mem<31><10> ), .B(n1774), .Y(n2837) );
  OAI21X1 U83 ( .A(n1773), .B(n1785), .C(n2836), .Y(n2310) );
  NAND2X1 U84 ( .A(\mem<31><11> ), .B(n1774), .Y(n2836) );
  OAI21X1 U85 ( .A(n1773), .B(n1784), .C(n2835), .Y(n2309) );
  NAND2X1 U86 ( .A(\mem<31><12> ), .B(n1774), .Y(n2835) );
  OAI21X1 U87 ( .A(n1773), .B(n1783), .C(n2834), .Y(n2308) );
  NAND2X1 U88 ( .A(\mem<31><13> ), .B(n1774), .Y(n2834) );
  OAI21X1 U89 ( .A(n1773), .B(n1781), .C(n2833), .Y(n2307) );
  NAND2X1 U90 ( .A(\mem<31><14> ), .B(n1774), .Y(n2833) );
  OAI21X1 U91 ( .A(n1773), .B(n1780), .C(n2832), .Y(n2306) );
  NAND2X1 U92 ( .A(\mem<31><15> ), .B(n1774), .Y(n2832) );
  OAI21X1 U95 ( .A(n1804), .B(n1770), .C(n2829), .Y(n2305) );
  NAND2X1 U96 ( .A(\mem<30><0> ), .B(n1772), .Y(n2829) );
  OAI21X1 U97 ( .A(n1802), .B(n1770), .C(n2828), .Y(n2304) );
  NAND2X1 U98 ( .A(\mem<30><1> ), .B(n1772), .Y(n2828) );
  OAI21X1 U99 ( .A(n1800), .B(n1770), .C(n2827), .Y(n2303) );
  NAND2X1 U100 ( .A(\mem<30><2> ), .B(n1772), .Y(n2827) );
  OAI21X1 U101 ( .A(n1798), .B(n1770), .C(n2826), .Y(n2302) );
  NAND2X1 U102 ( .A(\mem<30><3> ), .B(n1772), .Y(n2826) );
  OAI21X1 U103 ( .A(n1796), .B(n1770), .C(n2825), .Y(n2301) );
  NAND2X1 U104 ( .A(\mem<30><4> ), .B(n1772), .Y(n2825) );
  OAI21X1 U105 ( .A(n1794), .B(n1770), .C(n2824), .Y(n2300) );
  NAND2X1 U106 ( .A(\mem<30><5> ), .B(n1772), .Y(n2824) );
  OAI21X1 U107 ( .A(n1792), .B(n1770), .C(n2823), .Y(n2299) );
  NAND2X1 U108 ( .A(\mem<30><6> ), .B(n1772), .Y(n2823) );
  OAI21X1 U109 ( .A(n1790), .B(n1770), .C(n2822), .Y(n2298) );
  NAND2X1 U110 ( .A(\mem<30><7> ), .B(n1772), .Y(n2822) );
  OAI21X1 U111 ( .A(n1789), .B(n1770), .C(n2821), .Y(n2297) );
  NAND2X1 U112 ( .A(\mem<30><8> ), .B(n1771), .Y(n2821) );
  OAI21X1 U113 ( .A(n1788), .B(n1770), .C(n2820), .Y(n2296) );
  NAND2X1 U114 ( .A(\mem<30><9> ), .B(n1771), .Y(n2820) );
  OAI21X1 U115 ( .A(n1786), .B(n1770), .C(n2819), .Y(n2295) );
  NAND2X1 U116 ( .A(\mem<30><10> ), .B(n1771), .Y(n2819) );
  OAI21X1 U117 ( .A(n1785), .B(n1770), .C(n2818), .Y(n2294) );
  NAND2X1 U118 ( .A(\mem<30><11> ), .B(n1771), .Y(n2818) );
  OAI21X1 U119 ( .A(n1784), .B(n1770), .C(n2817), .Y(n2293) );
  NAND2X1 U120 ( .A(\mem<30><12> ), .B(n1771), .Y(n2817) );
  OAI21X1 U121 ( .A(n1783), .B(n1770), .C(n2816), .Y(n2292) );
  NAND2X1 U122 ( .A(\mem<30><13> ), .B(n1771), .Y(n2816) );
  OAI21X1 U123 ( .A(n1781), .B(n1770), .C(n2815), .Y(n2291) );
  NAND2X1 U124 ( .A(\mem<30><14> ), .B(n1771), .Y(n2815) );
  OAI21X1 U125 ( .A(n1780), .B(n1770), .C(n2814), .Y(n2290) );
  NAND2X1 U126 ( .A(\mem<30><15> ), .B(n1771), .Y(n2814) );
  OAI21X1 U129 ( .A(n1804), .B(n1767), .C(n2812), .Y(n2289) );
  NAND2X1 U130 ( .A(\mem<29><0> ), .B(n1769), .Y(n2812) );
  OAI21X1 U131 ( .A(n1802), .B(n1767), .C(n2811), .Y(n2288) );
  NAND2X1 U132 ( .A(\mem<29><1> ), .B(n1769), .Y(n2811) );
  OAI21X1 U133 ( .A(n1800), .B(n1767), .C(n2810), .Y(n2287) );
  NAND2X1 U134 ( .A(\mem<29><2> ), .B(n1769), .Y(n2810) );
  OAI21X1 U135 ( .A(n1798), .B(n1767), .C(n2809), .Y(n2286) );
  NAND2X1 U136 ( .A(\mem<29><3> ), .B(n1769), .Y(n2809) );
  OAI21X1 U137 ( .A(n1796), .B(n1767), .C(n2808), .Y(n2285) );
  NAND2X1 U138 ( .A(\mem<29><4> ), .B(n1769), .Y(n2808) );
  OAI21X1 U139 ( .A(n1794), .B(n1767), .C(n2807), .Y(n2284) );
  NAND2X1 U140 ( .A(\mem<29><5> ), .B(n1769), .Y(n2807) );
  OAI21X1 U141 ( .A(n1792), .B(n1767), .C(n2806), .Y(n2283) );
  NAND2X1 U142 ( .A(\mem<29><6> ), .B(n1769), .Y(n2806) );
  OAI21X1 U143 ( .A(n1790), .B(n1767), .C(n2805), .Y(n2282) );
  NAND2X1 U144 ( .A(\mem<29><7> ), .B(n1769), .Y(n2805) );
  OAI21X1 U145 ( .A(n1789), .B(n1767), .C(n2804), .Y(n2281) );
  NAND2X1 U146 ( .A(\mem<29><8> ), .B(n1768), .Y(n2804) );
  OAI21X1 U147 ( .A(n1788), .B(n1767), .C(n2803), .Y(n2280) );
  NAND2X1 U148 ( .A(\mem<29><9> ), .B(n1768), .Y(n2803) );
  OAI21X1 U149 ( .A(n1786), .B(n1767), .C(n2802), .Y(n2279) );
  NAND2X1 U150 ( .A(\mem<29><10> ), .B(n1768), .Y(n2802) );
  OAI21X1 U151 ( .A(n1785), .B(n1767), .C(n2801), .Y(n2278) );
  NAND2X1 U152 ( .A(\mem<29><11> ), .B(n1768), .Y(n2801) );
  OAI21X1 U153 ( .A(n1784), .B(n1767), .C(n2800), .Y(n2277) );
  NAND2X1 U154 ( .A(\mem<29><12> ), .B(n1768), .Y(n2800) );
  OAI21X1 U155 ( .A(n1783), .B(n1767), .C(n2799), .Y(n2276) );
  NAND2X1 U156 ( .A(\mem<29><13> ), .B(n1768), .Y(n2799) );
  OAI21X1 U157 ( .A(n1781), .B(n1767), .C(n2798), .Y(n2275) );
  NAND2X1 U158 ( .A(\mem<29><14> ), .B(n1768), .Y(n2798) );
  OAI21X1 U159 ( .A(n1780), .B(n1767), .C(n2797), .Y(n2274) );
  NAND2X1 U160 ( .A(\mem<29><15> ), .B(n1768), .Y(n2797) );
  OAI21X1 U163 ( .A(n1804), .B(n1764), .C(n2795), .Y(n2273) );
  NAND2X1 U164 ( .A(\mem<28><0> ), .B(n1766), .Y(n2795) );
  OAI21X1 U165 ( .A(n1802), .B(n1764), .C(n2794), .Y(n2272) );
  NAND2X1 U166 ( .A(\mem<28><1> ), .B(n1766), .Y(n2794) );
  OAI21X1 U167 ( .A(n1800), .B(n1764), .C(n2793), .Y(n2271) );
  NAND2X1 U168 ( .A(\mem<28><2> ), .B(n1766), .Y(n2793) );
  OAI21X1 U169 ( .A(n1798), .B(n1764), .C(n2792), .Y(n2270) );
  NAND2X1 U170 ( .A(\mem<28><3> ), .B(n1766), .Y(n2792) );
  OAI21X1 U171 ( .A(n1796), .B(n1764), .C(n2791), .Y(n2269) );
  NAND2X1 U172 ( .A(\mem<28><4> ), .B(n1766), .Y(n2791) );
  OAI21X1 U173 ( .A(n1794), .B(n1764), .C(n2790), .Y(n2268) );
  NAND2X1 U174 ( .A(\mem<28><5> ), .B(n1766), .Y(n2790) );
  OAI21X1 U175 ( .A(n1792), .B(n1764), .C(n2789), .Y(n2267) );
  NAND2X1 U176 ( .A(\mem<28><6> ), .B(n1766), .Y(n2789) );
  OAI21X1 U177 ( .A(n1790), .B(n1764), .C(n2788), .Y(n2266) );
  NAND2X1 U178 ( .A(\mem<28><7> ), .B(n1766), .Y(n2788) );
  OAI21X1 U179 ( .A(n1789), .B(n1764), .C(n2787), .Y(n2265) );
  NAND2X1 U180 ( .A(\mem<28><8> ), .B(n1765), .Y(n2787) );
  OAI21X1 U181 ( .A(n1788), .B(n1764), .C(n2786), .Y(n2264) );
  NAND2X1 U182 ( .A(\mem<28><9> ), .B(n1765), .Y(n2786) );
  OAI21X1 U183 ( .A(n1786), .B(n1764), .C(n2785), .Y(n2263) );
  NAND2X1 U184 ( .A(\mem<28><10> ), .B(n1765), .Y(n2785) );
  OAI21X1 U185 ( .A(n1785), .B(n1764), .C(n2784), .Y(n2262) );
  NAND2X1 U186 ( .A(\mem<28><11> ), .B(n1765), .Y(n2784) );
  OAI21X1 U187 ( .A(n1784), .B(n1764), .C(n2783), .Y(n2261) );
  NAND2X1 U188 ( .A(\mem<28><12> ), .B(n1765), .Y(n2783) );
  OAI21X1 U189 ( .A(n1783), .B(n1764), .C(n2782), .Y(n2260) );
  NAND2X1 U190 ( .A(\mem<28><13> ), .B(n1765), .Y(n2782) );
  OAI21X1 U191 ( .A(n1781), .B(n1764), .C(n2781), .Y(n2259) );
  NAND2X1 U192 ( .A(\mem<28><14> ), .B(n1765), .Y(n2781) );
  OAI21X1 U193 ( .A(n1780), .B(n1764), .C(n2780), .Y(n2258) );
  NAND2X1 U194 ( .A(\mem<28><15> ), .B(n1765), .Y(n2780) );
  OAI21X1 U197 ( .A(n1804), .B(n1761), .C(n2778), .Y(n2257) );
  NAND2X1 U198 ( .A(\mem<27><0> ), .B(n1763), .Y(n2778) );
  OAI21X1 U199 ( .A(n1802), .B(n1761), .C(n2777), .Y(n2256) );
  NAND2X1 U200 ( .A(\mem<27><1> ), .B(n1763), .Y(n2777) );
  OAI21X1 U201 ( .A(n1800), .B(n1761), .C(n2776), .Y(n2255) );
  NAND2X1 U202 ( .A(\mem<27><2> ), .B(n1763), .Y(n2776) );
  OAI21X1 U203 ( .A(n1798), .B(n1761), .C(n2775), .Y(n2254) );
  NAND2X1 U204 ( .A(\mem<27><3> ), .B(n1763), .Y(n2775) );
  OAI21X1 U205 ( .A(n1796), .B(n1761), .C(n2774), .Y(n2253) );
  NAND2X1 U206 ( .A(\mem<27><4> ), .B(n1763), .Y(n2774) );
  OAI21X1 U207 ( .A(n1794), .B(n1761), .C(n2773), .Y(n2252) );
  NAND2X1 U208 ( .A(\mem<27><5> ), .B(n1763), .Y(n2773) );
  OAI21X1 U209 ( .A(n1792), .B(n1761), .C(n2772), .Y(n2251) );
  NAND2X1 U210 ( .A(\mem<27><6> ), .B(n1763), .Y(n2772) );
  OAI21X1 U211 ( .A(n1790), .B(n1761), .C(n2771), .Y(n2250) );
  NAND2X1 U212 ( .A(\mem<27><7> ), .B(n1763), .Y(n2771) );
  OAI21X1 U213 ( .A(n1789), .B(n1761), .C(n2770), .Y(n2249) );
  NAND2X1 U214 ( .A(\mem<27><8> ), .B(n1762), .Y(n2770) );
  OAI21X1 U215 ( .A(n1788), .B(n1761), .C(n2769), .Y(n2248) );
  NAND2X1 U216 ( .A(\mem<27><9> ), .B(n1762), .Y(n2769) );
  OAI21X1 U217 ( .A(n1786), .B(n1761), .C(n2768), .Y(n2247) );
  NAND2X1 U218 ( .A(\mem<27><10> ), .B(n1762), .Y(n2768) );
  OAI21X1 U219 ( .A(n1785), .B(n1761), .C(n2767), .Y(n2246) );
  NAND2X1 U220 ( .A(\mem<27><11> ), .B(n1762), .Y(n2767) );
  OAI21X1 U221 ( .A(n1784), .B(n1761), .C(n2766), .Y(n2245) );
  NAND2X1 U222 ( .A(\mem<27><12> ), .B(n1762), .Y(n2766) );
  OAI21X1 U223 ( .A(n1783), .B(n1761), .C(n2765), .Y(n2244) );
  NAND2X1 U224 ( .A(\mem<27><13> ), .B(n1762), .Y(n2765) );
  OAI21X1 U225 ( .A(n1781), .B(n1761), .C(n2764), .Y(n2243) );
  NAND2X1 U226 ( .A(\mem<27><14> ), .B(n1762), .Y(n2764) );
  OAI21X1 U227 ( .A(n1780), .B(n1761), .C(n2763), .Y(n2242) );
  NAND2X1 U228 ( .A(\mem<27><15> ), .B(n1762), .Y(n2763) );
  OAI21X1 U231 ( .A(n1804), .B(n1758), .C(n2761), .Y(n2241) );
  NAND2X1 U232 ( .A(\mem<26><0> ), .B(n1760), .Y(n2761) );
  OAI21X1 U233 ( .A(n1802), .B(n1758), .C(n2760), .Y(n2240) );
  NAND2X1 U234 ( .A(\mem<26><1> ), .B(n1760), .Y(n2760) );
  OAI21X1 U235 ( .A(n1800), .B(n1758), .C(n2759), .Y(n2239) );
  NAND2X1 U236 ( .A(\mem<26><2> ), .B(n1760), .Y(n2759) );
  OAI21X1 U237 ( .A(n1798), .B(n1758), .C(n2758), .Y(n2238) );
  NAND2X1 U238 ( .A(\mem<26><3> ), .B(n1760), .Y(n2758) );
  OAI21X1 U239 ( .A(n1796), .B(n1758), .C(n2757), .Y(n2237) );
  NAND2X1 U240 ( .A(\mem<26><4> ), .B(n1760), .Y(n2757) );
  OAI21X1 U241 ( .A(n1794), .B(n1758), .C(n2756), .Y(n2236) );
  NAND2X1 U242 ( .A(\mem<26><5> ), .B(n1760), .Y(n2756) );
  OAI21X1 U243 ( .A(n1792), .B(n1758), .C(n2755), .Y(n2235) );
  NAND2X1 U244 ( .A(\mem<26><6> ), .B(n1760), .Y(n2755) );
  OAI21X1 U245 ( .A(n1790), .B(n1758), .C(n2754), .Y(n2234) );
  NAND2X1 U246 ( .A(\mem<26><7> ), .B(n1760), .Y(n2754) );
  OAI21X1 U247 ( .A(n1789), .B(n1758), .C(n2753), .Y(n2233) );
  NAND2X1 U248 ( .A(\mem<26><8> ), .B(n1759), .Y(n2753) );
  OAI21X1 U249 ( .A(n1788), .B(n1758), .C(n2752), .Y(n2232) );
  NAND2X1 U250 ( .A(\mem<26><9> ), .B(n1759), .Y(n2752) );
  OAI21X1 U251 ( .A(n1786), .B(n1758), .C(n2751), .Y(n2231) );
  NAND2X1 U252 ( .A(\mem<26><10> ), .B(n1759), .Y(n2751) );
  OAI21X1 U253 ( .A(n1785), .B(n1758), .C(n2750), .Y(n2230) );
  NAND2X1 U254 ( .A(\mem<26><11> ), .B(n1759), .Y(n2750) );
  OAI21X1 U255 ( .A(n1784), .B(n1758), .C(n2749), .Y(n2229) );
  NAND2X1 U256 ( .A(\mem<26><12> ), .B(n1759), .Y(n2749) );
  OAI21X1 U257 ( .A(n1783), .B(n1758), .C(n2748), .Y(n2228) );
  NAND2X1 U258 ( .A(\mem<26><13> ), .B(n1759), .Y(n2748) );
  OAI21X1 U259 ( .A(n1781), .B(n1758), .C(n2747), .Y(n2227) );
  NAND2X1 U260 ( .A(\mem<26><14> ), .B(n1759), .Y(n2747) );
  OAI21X1 U261 ( .A(n1780), .B(n1758), .C(n2746), .Y(n2226) );
  NAND2X1 U262 ( .A(\mem<26><15> ), .B(n1759), .Y(n2746) );
  OAI21X1 U265 ( .A(n1804), .B(n1755), .C(n2744), .Y(n2225) );
  NAND2X1 U266 ( .A(\mem<25><0> ), .B(n1757), .Y(n2744) );
  OAI21X1 U267 ( .A(n1802), .B(n1755), .C(n2743), .Y(n2224) );
  NAND2X1 U268 ( .A(\mem<25><1> ), .B(n1757), .Y(n2743) );
  OAI21X1 U269 ( .A(n1800), .B(n1755), .C(n2742), .Y(n2223) );
  NAND2X1 U270 ( .A(\mem<25><2> ), .B(n1757), .Y(n2742) );
  OAI21X1 U271 ( .A(n1798), .B(n1755), .C(n2741), .Y(n2222) );
  NAND2X1 U272 ( .A(\mem<25><3> ), .B(n1757), .Y(n2741) );
  OAI21X1 U273 ( .A(n1796), .B(n1755), .C(n2740), .Y(n2221) );
  NAND2X1 U274 ( .A(\mem<25><4> ), .B(n1757), .Y(n2740) );
  OAI21X1 U275 ( .A(n1794), .B(n1755), .C(n2739), .Y(n2220) );
  NAND2X1 U276 ( .A(\mem<25><5> ), .B(n1757), .Y(n2739) );
  OAI21X1 U277 ( .A(n1792), .B(n1755), .C(n2738), .Y(n2219) );
  NAND2X1 U278 ( .A(\mem<25><6> ), .B(n1757), .Y(n2738) );
  OAI21X1 U279 ( .A(n1790), .B(n1755), .C(n2737), .Y(n2218) );
  NAND2X1 U280 ( .A(\mem<25><7> ), .B(n1757), .Y(n2737) );
  OAI21X1 U281 ( .A(n1789), .B(n1755), .C(n2736), .Y(n2217) );
  NAND2X1 U282 ( .A(\mem<25><8> ), .B(n1756), .Y(n2736) );
  OAI21X1 U283 ( .A(n1788), .B(n1755), .C(n2735), .Y(n2216) );
  NAND2X1 U284 ( .A(\mem<25><9> ), .B(n1756), .Y(n2735) );
  OAI21X1 U285 ( .A(n1786), .B(n1755), .C(n2734), .Y(n2215) );
  NAND2X1 U286 ( .A(\mem<25><10> ), .B(n1756), .Y(n2734) );
  OAI21X1 U287 ( .A(n1785), .B(n1755), .C(n2733), .Y(n2214) );
  NAND2X1 U288 ( .A(\mem<25><11> ), .B(n1756), .Y(n2733) );
  OAI21X1 U289 ( .A(n1784), .B(n1755), .C(n2732), .Y(n2213) );
  NAND2X1 U290 ( .A(\mem<25><12> ), .B(n1756), .Y(n2732) );
  OAI21X1 U291 ( .A(n1783), .B(n1755), .C(n2731), .Y(n2212) );
  NAND2X1 U292 ( .A(\mem<25><13> ), .B(n1756), .Y(n2731) );
  OAI21X1 U293 ( .A(n1781), .B(n1755), .C(n2730), .Y(n2211) );
  NAND2X1 U294 ( .A(\mem<25><14> ), .B(n1756), .Y(n2730) );
  OAI21X1 U295 ( .A(n1780), .B(n1755), .C(n2729), .Y(n2210) );
  NAND2X1 U296 ( .A(\mem<25><15> ), .B(n1756), .Y(n2729) );
  OAI21X1 U299 ( .A(n1804), .B(n1752), .C(n2727), .Y(n2209) );
  NAND2X1 U300 ( .A(\mem<24><0> ), .B(n1754), .Y(n2727) );
  OAI21X1 U301 ( .A(n1802), .B(n1752), .C(n2726), .Y(n2208) );
  NAND2X1 U302 ( .A(\mem<24><1> ), .B(n1754), .Y(n2726) );
  OAI21X1 U303 ( .A(n1800), .B(n1752), .C(n2725), .Y(n2207) );
  NAND2X1 U304 ( .A(\mem<24><2> ), .B(n1754), .Y(n2725) );
  OAI21X1 U305 ( .A(n1798), .B(n1752), .C(n2724), .Y(n2206) );
  NAND2X1 U306 ( .A(\mem<24><3> ), .B(n1754), .Y(n2724) );
  OAI21X1 U307 ( .A(n1796), .B(n1752), .C(n2723), .Y(n2205) );
  NAND2X1 U308 ( .A(\mem<24><4> ), .B(n1754), .Y(n2723) );
  OAI21X1 U309 ( .A(n1794), .B(n1752), .C(n2722), .Y(n2204) );
  NAND2X1 U310 ( .A(\mem<24><5> ), .B(n1754), .Y(n2722) );
  OAI21X1 U311 ( .A(n1792), .B(n1752), .C(n2721), .Y(n2203) );
  NAND2X1 U312 ( .A(\mem<24><6> ), .B(n1754), .Y(n2721) );
  OAI21X1 U313 ( .A(n1790), .B(n1752), .C(n2720), .Y(n2202) );
  NAND2X1 U314 ( .A(\mem<24><7> ), .B(n1754), .Y(n2720) );
  OAI21X1 U315 ( .A(n1789), .B(n1752), .C(n2719), .Y(n2201) );
  NAND2X1 U316 ( .A(\mem<24><8> ), .B(n1753), .Y(n2719) );
  OAI21X1 U317 ( .A(n1788), .B(n1752), .C(n2718), .Y(n2200) );
  NAND2X1 U318 ( .A(\mem<24><9> ), .B(n1753), .Y(n2718) );
  OAI21X1 U319 ( .A(n1786), .B(n1752), .C(n2717), .Y(n2199) );
  NAND2X1 U320 ( .A(\mem<24><10> ), .B(n1753), .Y(n2717) );
  OAI21X1 U321 ( .A(n1785), .B(n1752), .C(n2716), .Y(n2198) );
  NAND2X1 U322 ( .A(\mem<24><11> ), .B(n1753), .Y(n2716) );
  OAI21X1 U323 ( .A(n1784), .B(n1752), .C(n2715), .Y(n2197) );
  NAND2X1 U324 ( .A(\mem<24><12> ), .B(n1753), .Y(n2715) );
  OAI21X1 U325 ( .A(n1783), .B(n1752), .C(n2714), .Y(n2196) );
  NAND2X1 U326 ( .A(\mem<24><13> ), .B(n1753), .Y(n2714) );
  OAI21X1 U327 ( .A(n1781), .B(n1752), .C(n2713), .Y(n2195) );
  NAND2X1 U328 ( .A(\mem<24><14> ), .B(n1753), .Y(n2713) );
  OAI21X1 U329 ( .A(n1780), .B(n1752), .C(n2712), .Y(n2194) );
  NAND2X1 U330 ( .A(\mem<24><15> ), .B(n1753), .Y(n2712) );
  NAND3X1 U333 ( .A(net59458), .B(n2709), .C(N14), .Y(n2710) );
  OAI21X1 U334 ( .A(n1804), .B(n1749), .C(n2708), .Y(n2193) );
  NAND2X1 U335 ( .A(\mem<23><0> ), .B(n1751), .Y(n2708) );
  OAI21X1 U336 ( .A(n1802), .B(n1749), .C(n2707), .Y(n2192) );
  NAND2X1 U337 ( .A(\mem<23><1> ), .B(n1751), .Y(n2707) );
  OAI21X1 U338 ( .A(n1800), .B(n1749), .C(n2706), .Y(n2191) );
  NAND2X1 U339 ( .A(\mem<23><2> ), .B(n1751), .Y(n2706) );
  OAI21X1 U340 ( .A(n1798), .B(n1749), .C(n2705), .Y(n2190) );
  NAND2X1 U341 ( .A(\mem<23><3> ), .B(n1751), .Y(n2705) );
  OAI21X1 U342 ( .A(n1796), .B(n1749), .C(n2704), .Y(n2189) );
  NAND2X1 U343 ( .A(\mem<23><4> ), .B(n1751), .Y(n2704) );
  OAI21X1 U344 ( .A(n1794), .B(n1749), .C(n2703), .Y(n2188) );
  NAND2X1 U345 ( .A(\mem<23><5> ), .B(n1751), .Y(n2703) );
  OAI21X1 U346 ( .A(n1792), .B(n1749), .C(n2702), .Y(n2187) );
  NAND2X1 U347 ( .A(\mem<23><6> ), .B(n1751), .Y(n2702) );
  OAI21X1 U348 ( .A(n1790), .B(n1749), .C(n2701), .Y(n2186) );
  NAND2X1 U349 ( .A(\mem<23><7> ), .B(n1751), .Y(n2701) );
  OAI21X1 U350 ( .A(n1789), .B(n1749), .C(n2700), .Y(n2185) );
  NAND2X1 U351 ( .A(\mem<23><8> ), .B(n1750), .Y(n2700) );
  OAI21X1 U352 ( .A(n1788), .B(n1749), .C(n2699), .Y(n2184) );
  NAND2X1 U353 ( .A(\mem<23><9> ), .B(n1750), .Y(n2699) );
  OAI21X1 U354 ( .A(n1786), .B(n1749), .C(n2698), .Y(n2183) );
  NAND2X1 U355 ( .A(\mem<23><10> ), .B(n1750), .Y(n2698) );
  OAI21X1 U356 ( .A(n1785), .B(n1749), .C(n2697), .Y(n2182) );
  NAND2X1 U357 ( .A(\mem<23><11> ), .B(n1750), .Y(n2697) );
  OAI21X1 U358 ( .A(n1784), .B(n1749), .C(n2696), .Y(n2181) );
  NAND2X1 U359 ( .A(\mem<23><12> ), .B(n1750), .Y(n2696) );
  OAI21X1 U360 ( .A(n1783), .B(n1749), .C(n2695), .Y(n2180) );
  NAND2X1 U361 ( .A(\mem<23><13> ), .B(n1750), .Y(n2695) );
  OAI21X1 U362 ( .A(n1781), .B(n1749), .C(n2694), .Y(n2179) );
  NAND2X1 U363 ( .A(\mem<23><14> ), .B(n1750), .Y(n2694) );
  OAI21X1 U364 ( .A(n1780), .B(n1749), .C(n2693), .Y(n2178) );
  NAND2X1 U365 ( .A(\mem<23><15> ), .B(n1750), .Y(n2693) );
  OAI21X1 U368 ( .A(n1804), .B(n1746), .C(n2692), .Y(n2177) );
  NAND2X1 U369 ( .A(\mem<22><0> ), .B(n1748), .Y(n2692) );
  OAI21X1 U370 ( .A(n1802), .B(n1746), .C(n2691), .Y(n2176) );
  NAND2X1 U371 ( .A(\mem<22><1> ), .B(n1748), .Y(n2691) );
  OAI21X1 U372 ( .A(n1800), .B(n1746), .C(n2690), .Y(n2175) );
  NAND2X1 U373 ( .A(\mem<22><2> ), .B(n1748), .Y(n2690) );
  OAI21X1 U374 ( .A(n1798), .B(n1746), .C(n2689), .Y(n2174) );
  NAND2X1 U375 ( .A(\mem<22><3> ), .B(n1748), .Y(n2689) );
  OAI21X1 U376 ( .A(n1796), .B(n1746), .C(n2688), .Y(n2173) );
  NAND2X1 U377 ( .A(\mem<22><4> ), .B(n1748), .Y(n2688) );
  OAI21X1 U378 ( .A(n1794), .B(n1746), .C(n2687), .Y(n2172) );
  NAND2X1 U379 ( .A(\mem<22><5> ), .B(n1748), .Y(n2687) );
  OAI21X1 U380 ( .A(n1792), .B(n1746), .C(n2686), .Y(n2171) );
  NAND2X1 U381 ( .A(\mem<22><6> ), .B(n1748), .Y(n2686) );
  OAI21X1 U382 ( .A(n1790), .B(n1746), .C(n2685), .Y(n2170) );
  NAND2X1 U383 ( .A(\mem<22><7> ), .B(n1748), .Y(n2685) );
  OAI21X1 U384 ( .A(n1789), .B(n1746), .C(n2684), .Y(n2169) );
  NAND2X1 U385 ( .A(\mem<22><8> ), .B(n1747), .Y(n2684) );
  OAI21X1 U386 ( .A(n1788), .B(n1746), .C(n2683), .Y(n2168) );
  NAND2X1 U387 ( .A(\mem<22><9> ), .B(n1747), .Y(n2683) );
  OAI21X1 U388 ( .A(n1786), .B(n1746), .C(n2682), .Y(n2167) );
  NAND2X1 U389 ( .A(\mem<22><10> ), .B(n1747), .Y(n2682) );
  OAI21X1 U390 ( .A(n1785), .B(n1746), .C(n2681), .Y(n2166) );
  NAND2X1 U391 ( .A(\mem<22><11> ), .B(n1747), .Y(n2681) );
  OAI21X1 U392 ( .A(n1784), .B(n1746), .C(n2680), .Y(n2165) );
  NAND2X1 U393 ( .A(\mem<22><12> ), .B(n1747), .Y(n2680) );
  OAI21X1 U394 ( .A(n1783), .B(n1746), .C(n2679), .Y(n2164) );
  NAND2X1 U395 ( .A(\mem<22><13> ), .B(n1747), .Y(n2679) );
  OAI21X1 U396 ( .A(n1781), .B(n1746), .C(n2678), .Y(n2163) );
  NAND2X1 U397 ( .A(\mem<22><14> ), .B(n1747), .Y(n2678) );
  OAI21X1 U398 ( .A(n1780), .B(n1746), .C(n2677), .Y(n2162) );
  NAND2X1 U399 ( .A(\mem<22><15> ), .B(n1747), .Y(n2677) );
  OAI21X1 U402 ( .A(n1804), .B(n1743), .C(n2676), .Y(n2161) );
  NAND2X1 U403 ( .A(\mem<21><0> ), .B(n1745), .Y(n2676) );
  OAI21X1 U404 ( .A(n1802), .B(n1743), .C(n2675), .Y(n2160) );
  NAND2X1 U405 ( .A(\mem<21><1> ), .B(n1745), .Y(n2675) );
  OAI21X1 U406 ( .A(n1800), .B(n1743), .C(n2674), .Y(n2159) );
  NAND2X1 U407 ( .A(\mem<21><2> ), .B(n1745), .Y(n2674) );
  OAI21X1 U408 ( .A(n1798), .B(n1743), .C(n2673), .Y(n2158) );
  NAND2X1 U409 ( .A(\mem<21><3> ), .B(n1745), .Y(n2673) );
  OAI21X1 U410 ( .A(n1796), .B(n1743), .C(n2672), .Y(n2157) );
  NAND2X1 U411 ( .A(\mem<21><4> ), .B(n1745), .Y(n2672) );
  OAI21X1 U412 ( .A(n1794), .B(n1743), .C(n2671), .Y(n2156) );
  NAND2X1 U413 ( .A(\mem<21><5> ), .B(n1745), .Y(n2671) );
  OAI21X1 U414 ( .A(n1792), .B(n1743), .C(n2670), .Y(n2155) );
  NAND2X1 U415 ( .A(\mem<21><6> ), .B(n1745), .Y(n2670) );
  OAI21X1 U416 ( .A(n1790), .B(n1743), .C(n2669), .Y(n2154) );
  NAND2X1 U417 ( .A(\mem<21><7> ), .B(n1745), .Y(n2669) );
  OAI21X1 U418 ( .A(n1789), .B(n1743), .C(n2668), .Y(n2153) );
  NAND2X1 U419 ( .A(\mem<21><8> ), .B(n1744), .Y(n2668) );
  OAI21X1 U420 ( .A(n1788), .B(n1743), .C(n2667), .Y(n2152) );
  NAND2X1 U421 ( .A(\mem<21><9> ), .B(n1744), .Y(n2667) );
  OAI21X1 U422 ( .A(n1786), .B(n1743), .C(n2666), .Y(n2151) );
  NAND2X1 U423 ( .A(\mem<21><10> ), .B(n1744), .Y(n2666) );
  OAI21X1 U424 ( .A(n1785), .B(n1743), .C(n2665), .Y(n2150) );
  NAND2X1 U425 ( .A(\mem<21><11> ), .B(n1744), .Y(n2665) );
  OAI21X1 U426 ( .A(n1784), .B(n1743), .C(n2664), .Y(n2149) );
  NAND2X1 U427 ( .A(\mem<21><12> ), .B(n1744), .Y(n2664) );
  OAI21X1 U428 ( .A(n1783), .B(n1743), .C(n2663), .Y(n2148) );
  NAND2X1 U429 ( .A(\mem<21><13> ), .B(n1744), .Y(n2663) );
  OAI21X1 U430 ( .A(n1781), .B(n1743), .C(n2662), .Y(n2147) );
  NAND2X1 U431 ( .A(\mem<21><14> ), .B(n1744), .Y(n2662) );
  OAI21X1 U432 ( .A(n1780), .B(n1743), .C(n2661), .Y(n2146) );
  NAND2X1 U433 ( .A(\mem<21><15> ), .B(n1744), .Y(n2661) );
  OAI21X1 U436 ( .A(n1804), .B(n1740), .C(n2660), .Y(n2145) );
  NAND2X1 U437 ( .A(\mem<20><0> ), .B(n1742), .Y(n2660) );
  OAI21X1 U438 ( .A(n1802), .B(n1740), .C(n2659), .Y(n2144) );
  NAND2X1 U439 ( .A(\mem<20><1> ), .B(n1742), .Y(n2659) );
  OAI21X1 U440 ( .A(n1800), .B(n1740), .C(n2658), .Y(n2143) );
  NAND2X1 U441 ( .A(\mem<20><2> ), .B(n1742), .Y(n2658) );
  OAI21X1 U442 ( .A(n1798), .B(n1740), .C(n2657), .Y(n2142) );
  NAND2X1 U443 ( .A(\mem<20><3> ), .B(n1742), .Y(n2657) );
  OAI21X1 U444 ( .A(n1796), .B(n1740), .C(n2656), .Y(n2141) );
  NAND2X1 U445 ( .A(\mem<20><4> ), .B(n1742), .Y(n2656) );
  OAI21X1 U446 ( .A(n1794), .B(n1740), .C(n2655), .Y(n2140) );
  NAND2X1 U447 ( .A(\mem<20><5> ), .B(n1742), .Y(n2655) );
  OAI21X1 U448 ( .A(n1792), .B(n1740), .C(n2654), .Y(n2139) );
  NAND2X1 U449 ( .A(\mem<20><6> ), .B(n1742), .Y(n2654) );
  OAI21X1 U450 ( .A(n1790), .B(n1740), .C(n2653), .Y(n2138) );
  NAND2X1 U451 ( .A(\mem<20><7> ), .B(n1742), .Y(n2653) );
  OAI21X1 U452 ( .A(n1789), .B(n1740), .C(n2652), .Y(n2137) );
  NAND2X1 U453 ( .A(\mem<20><8> ), .B(n1741), .Y(n2652) );
  OAI21X1 U454 ( .A(n1788), .B(n1740), .C(n2651), .Y(n2136) );
  NAND2X1 U455 ( .A(\mem<20><9> ), .B(n1741), .Y(n2651) );
  OAI21X1 U456 ( .A(n1786), .B(n1740), .C(n2650), .Y(n2135) );
  NAND2X1 U457 ( .A(\mem<20><10> ), .B(n1741), .Y(n2650) );
  OAI21X1 U458 ( .A(n1785), .B(n1740), .C(n2649), .Y(n2134) );
  NAND2X1 U459 ( .A(\mem<20><11> ), .B(n1741), .Y(n2649) );
  OAI21X1 U460 ( .A(n1784), .B(n1740), .C(n2648), .Y(n2133) );
  NAND2X1 U461 ( .A(\mem<20><12> ), .B(n1741), .Y(n2648) );
  OAI21X1 U462 ( .A(n1783), .B(n1740), .C(n2647), .Y(n2132) );
  NAND2X1 U463 ( .A(\mem<20><13> ), .B(n1741), .Y(n2647) );
  OAI21X1 U464 ( .A(n1781), .B(n1740), .C(n2646), .Y(n2131) );
  NAND2X1 U465 ( .A(\mem<20><14> ), .B(n1741), .Y(n2646) );
  OAI21X1 U466 ( .A(n1780), .B(n1740), .C(n2645), .Y(n2130) );
  NAND2X1 U467 ( .A(\mem<20><15> ), .B(n1741), .Y(n2645) );
  OAI21X1 U470 ( .A(n1804), .B(n1737), .C(n2644), .Y(n2129) );
  NAND2X1 U471 ( .A(\mem<19><0> ), .B(n1739), .Y(n2644) );
  OAI21X1 U472 ( .A(n1802), .B(n1737), .C(n2643), .Y(n2128) );
  NAND2X1 U473 ( .A(\mem<19><1> ), .B(n1739), .Y(n2643) );
  OAI21X1 U474 ( .A(n1800), .B(n1737), .C(n2642), .Y(n2127) );
  NAND2X1 U475 ( .A(\mem<19><2> ), .B(n1739), .Y(n2642) );
  OAI21X1 U476 ( .A(n1798), .B(n1737), .C(n2641), .Y(n2126) );
  NAND2X1 U477 ( .A(\mem<19><3> ), .B(n1739), .Y(n2641) );
  OAI21X1 U478 ( .A(n1796), .B(n1737), .C(n2640), .Y(n2125) );
  NAND2X1 U479 ( .A(\mem<19><4> ), .B(n1739), .Y(n2640) );
  OAI21X1 U480 ( .A(n1794), .B(n1737), .C(n2639), .Y(n2124) );
  NAND2X1 U481 ( .A(\mem<19><5> ), .B(n1739), .Y(n2639) );
  OAI21X1 U482 ( .A(n1792), .B(n1737), .C(n2638), .Y(n2123) );
  NAND2X1 U483 ( .A(\mem<19><6> ), .B(n1739), .Y(n2638) );
  OAI21X1 U484 ( .A(n1790), .B(n1737), .C(n2637), .Y(n2122) );
  NAND2X1 U485 ( .A(\mem<19><7> ), .B(n1739), .Y(n2637) );
  OAI21X1 U486 ( .A(n1789), .B(n1737), .C(n2636), .Y(n2121) );
  NAND2X1 U487 ( .A(\mem<19><8> ), .B(n1738), .Y(n2636) );
  OAI21X1 U488 ( .A(n1788), .B(n1737), .C(n2635), .Y(n2120) );
  NAND2X1 U489 ( .A(\mem<19><9> ), .B(n1738), .Y(n2635) );
  OAI21X1 U490 ( .A(n1786), .B(n1737), .C(n2634), .Y(n2119) );
  NAND2X1 U491 ( .A(\mem<19><10> ), .B(n1738), .Y(n2634) );
  OAI21X1 U492 ( .A(n1785), .B(n1737), .C(n2633), .Y(n2118) );
  NAND2X1 U493 ( .A(\mem<19><11> ), .B(n1738), .Y(n2633) );
  OAI21X1 U494 ( .A(n1784), .B(n1737), .C(n2632), .Y(n2117) );
  NAND2X1 U495 ( .A(\mem<19><12> ), .B(n1738), .Y(n2632) );
  OAI21X1 U496 ( .A(n1783), .B(n1737), .C(n2631), .Y(n2116) );
  NAND2X1 U497 ( .A(\mem<19><13> ), .B(n1738), .Y(n2631) );
  OAI21X1 U498 ( .A(n1781), .B(n1737), .C(n2630), .Y(n2115) );
  NAND2X1 U499 ( .A(\mem<19><14> ), .B(n1738), .Y(n2630) );
  OAI21X1 U500 ( .A(n1780), .B(n1737), .C(n2629), .Y(n2114) );
  NAND2X1 U501 ( .A(\mem<19><15> ), .B(n1738), .Y(n2629) );
  OAI21X1 U504 ( .A(n1805), .B(n1734), .C(n2628), .Y(n2113) );
  NAND2X1 U505 ( .A(\mem<18><0> ), .B(n1736), .Y(n2628) );
  OAI21X1 U506 ( .A(n1803), .B(n1734), .C(n2627), .Y(n2112) );
  NAND2X1 U507 ( .A(\mem<18><1> ), .B(n1736), .Y(n2627) );
  OAI21X1 U508 ( .A(n1801), .B(n1734), .C(n2626), .Y(n2111) );
  NAND2X1 U509 ( .A(\mem<18><2> ), .B(n1736), .Y(n2626) );
  OAI21X1 U510 ( .A(n1799), .B(n1734), .C(n2625), .Y(n2110) );
  NAND2X1 U511 ( .A(\mem<18><3> ), .B(n1736), .Y(n2625) );
  OAI21X1 U512 ( .A(n1797), .B(n1734), .C(n2624), .Y(n2109) );
  NAND2X1 U513 ( .A(\mem<18><4> ), .B(n1736), .Y(n2624) );
  OAI21X1 U514 ( .A(n1795), .B(n1734), .C(n2623), .Y(n2108) );
  NAND2X1 U515 ( .A(\mem<18><5> ), .B(n1736), .Y(n2623) );
  OAI21X1 U516 ( .A(n1793), .B(n1734), .C(n2622), .Y(n2107) );
  NAND2X1 U517 ( .A(\mem<18><6> ), .B(n1736), .Y(n2622) );
  OAI21X1 U518 ( .A(n1791), .B(n1734), .C(n2621), .Y(n2106) );
  NAND2X1 U519 ( .A(\mem<18><7> ), .B(n1736), .Y(n2621) );
  OAI21X1 U520 ( .A(n1789), .B(n1734), .C(n2620), .Y(n2105) );
  NAND2X1 U521 ( .A(\mem<18><8> ), .B(n1735), .Y(n2620) );
  OAI21X1 U522 ( .A(n1788), .B(n1734), .C(n2619), .Y(n2104) );
  NAND2X1 U523 ( .A(\mem<18><9> ), .B(n1735), .Y(n2619) );
  OAI21X1 U524 ( .A(n1787), .B(n1734), .C(n2618), .Y(n2103) );
  NAND2X1 U525 ( .A(\mem<18><10> ), .B(n1735), .Y(n2618) );
  OAI21X1 U526 ( .A(n1785), .B(n1734), .C(n2617), .Y(n2102) );
  NAND2X1 U527 ( .A(\mem<18><11> ), .B(n1735), .Y(n2617) );
  OAI21X1 U528 ( .A(n1784), .B(n1734), .C(n2616), .Y(n2101) );
  NAND2X1 U529 ( .A(\mem<18><12> ), .B(n1735), .Y(n2616) );
  OAI21X1 U530 ( .A(n1783), .B(n1734), .C(n2615), .Y(n2100) );
  NAND2X1 U531 ( .A(\mem<18><13> ), .B(n1735), .Y(n2615) );
  OAI21X1 U532 ( .A(n1782), .B(n1734), .C(n2614), .Y(n2099) );
  NAND2X1 U533 ( .A(\mem<18><14> ), .B(n1735), .Y(n2614) );
  OAI21X1 U534 ( .A(n1780), .B(n1734), .C(n2613), .Y(n2098) );
  NAND2X1 U535 ( .A(\mem<18><15> ), .B(n1735), .Y(n2613) );
  OAI21X1 U538 ( .A(n1805), .B(n1731), .C(n2612), .Y(n2097) );
  NAND2X1 U539 ( .A(\mem<17><0> ), .B(n1733), .Y(n2612) );
  OAI21X1 U540 ( .A(n1803), .B(n1731), .C(n2611), .Y(n2096) );
  NAND2X1 U541 ( .A(\mem<17><1> ), .B(n1733), .Y(n2611) );
  OAI21X1 U542 ( .A(n1801), .B(n1731), .C(n2610), .Y(n2095) );
  NAND2X1 U543 ( .A(\mem<17><2> ), .B(n1733), .Y(n2610) );
  OAI21X1 U544 ( .A(n1799), .B(n1731), .C(n2609), .Y(n2094) );
  NAND2X1 U545 ( .A(\mem<17><3> ), .B(n1733), .Y(n2609) );
  OAI21X1 U546 ( .A(n1797), .B(n1731), .C(n2608), .Y(n2093) );
  NAND2X1 U547 ( .A(\mem<17><4> ), .B(n1733), .Y(n2608) );
  OAI21X1 U548 ( .A(n1795), .B(n1731), .C(n2607), .Y(n2092) );
  NAND2X1 U549 ( .A(\mem<17><5> ), .B(n1733), .Y(n2607) );
  OAI21X1 U550 ( .A(n1793), .B(n1731), .C(n2606), .Y(n2091) );
  NAND2X1 U551 ( .A(\mem<17><6> ), .B(n1733), .Y(n2606) );
  OAI21X1 U552 ( .A(n1791), .B(n1731), .C(n2605), .Y(n2090) );
  NAND2X1 U553 ( .A(\mem<17><7> ), .B(n1733), .Y(n2605) );
  OAI21X1 U554 ( .A(n1789), .B(n1731), .C(n2604), .Y(n2089) );
  NAND2X1 U555 ( .A(\mem<17><8> ), .B(n1732), .Y(n2604) );
  OAI21X1 U556 ( .A(n1788), .B(n1731), .C(n2603), .Y(n2088) );
  NAND2X1 U557 ( .A(\mem<17><9> ), .B(n1732), .Y(n2603) );
  OAI21X1 U558 ( .A(n1787), .B(n1731), .C(n2602), .Y(n2087) );
  NAND2X1 U559 ( .A(\mem<17><10> ), .B(n1732), .Y(n2602) );
  OAI21X1 U560 ( .A(n1785), .B(n1731), .C(n2601), .Y(n2086) );
  NAND2X1 U561 ( .A(\mem<17><11> ), .B(n1732), .Y(n2601) );
  OAI21X1 U562 ( .A(n1784), .B(n1731), .C(n2600), .Y(n2085) );
  NAND2X1 U563 ( .A(\mem<17><12> ), .B(n1732), .Y(n2600) );
  OAI21X1 U564 ( .A(n1783), .B(n1731), .C(n2599), .Y(n2084) );
  NAND2X1 U565 ( .A(\mem<17><13> ), .B(n1732), .Y(n2599) );
  OAI21X1 U566 ( .A(n1782), .B(n1731), .C(n2598), .Y(n2083) );
  NAND2X1 U567 ( .A(\mem<17><14> ), .B(n1732), .Y(n2598) );
  OAI21X1 U568 ( .A(n1780), .B(n1731), .C(n2597), .Y(n2082) );
  NAND2X1 U569 ( .A(\mem<17><15> ), .B(n1732), .Y(n2597) );
  OAI21X1 U572 ( .A(n1805), .B(n1728), .C(n2596), .Y(n2081) );
  NAND2X1 U573 ( .A(\mem<16><0> ), .B(n1730), .Y(n2596) );
  OAI21X1 U574 ( .A(n1803), .B(n1728), .C(n2595), .Y(n2080) );
  NAND2X1 U575 ( .A(\mem<16><1> ), .B(n1730), .Y(n2595) );
  OAI21X1 U576 ( .A(n1801), .B(n1728), .C(n2594), .Y(n2079) );
  NAND2X1 U577 ( .A(\mem<16><2> ), .B(n1730), .Y(n2594) );
  OAI21X1 U578 ( .A(n1799), .B(n1728), .C(n2593), .Y(n2078) );
  NAND2X1 U579 ( .A(\mem<16><3> ), .B(n1730), .Y(n2593) );
  OAI21X1 U580 ( .A(n1797), .B(n1728), .C(n2592), .Y(n2077) );
  NAND2X1 U581 ( .A(\mem<16><4> ), .B(n1730), .Y(n2592) );
  OAI21X1 U582 ( .A(n1795), .B(n1728), .C(n2591), .Y(n2076) );
  NAND2X1 U583 ( .A(\mem<16><5> ), .B(n1730), .Y(n2591) );
  OAI21X1 U584 ( .A(n1793), .B(n1728), .C(n2590), .Y(n2075) );
  NAND2X1 U585 ( .A(\mem<16><6> ), .B(n1730), .Y(n2590) );
  OAI21X1 U586 ( .A(n1791), .B(n1728), .C(n2589), .Y(n2074) );
  NAND2X1 U587 ( .A(\mem<16><7> ), .B(n1730), .Y(n2589) );
  OAI21X1 U588 ( .A(n1789), .B(n1728), .C(n2588), .Y(n2073) );
  NAND2X1 U589 ( .A(\mem<16><8> ), .B(n1729), .Y(n2588) );
  OAI21X1 U590 ( .A(n1788), .B(n1728), .C(n2587), .Y(n2072) );
  NAND2X1 U591 ( .A(\mem<16><9> ), .B(n1729), .Y(n2587) );
  OAI21X1 U592 ( .A(n1787), .B(n1728), .C(n2586), .Y(n2071) );
  NAND2X1 U593 ( .A(\mem<16><10> ), .B(n1729), .Y(n2586) );
  OAI21X1 U594 ( .A(n1785), .B(n1728), .C(n2585), .Y(n2070) );
  NAND2X1 U595 ( .A(\mem<16><11> ), .B(n1729), .Y(n2585) );
  OAI21X1 U596 ( .A(n1784), .B(n1728), .C(n2584), .Y(n2069) );
  NAND2X1 U597 ( .A(\mem<16><12> ), .B(n1729), .Y(n2584) );
  OAI21X1 U598 ( .A(n1783), .B(n1728), .C(n2583), .Y(n2068) );
  NAND2X1 U599 ( .A(\mem<16><13> ), .B(n1729), .Y(n2583) );
  OAI21X1 U600 ( .A(n1782), .B(n1728), .C(n2582), .Y(n2067) );
  NAND2X1 U601 ( .A(\mem<16><14> ), .B(n1729), .Y(n2582) );
  OAI21X1 U602 ( .A(n1780), .B(n1728), .C(n2581), .Y(n2066) );
  NAND2X1 U603 ( .A(\mem<16><15> ), .B(n1729), .Y(n2581) );
  NAND3X1 U606 ( .A(n2709), .B(net59460), .C(N14), .Y(n2580) );
  OAI21X1 U607 ( .A(n1805), .B(n1725), .C(n2579), .Y(n2065) );
  NAND2X1 U608 ( .A(\mem<15><0> ), .B(n1727), .Y(n2579) );
  OAI21X1 U609 ( .A(n1803), .B(n1725), .C(n2578), .Y(n2064) );
  NAND2X1 U610 ( .A(\mem<15><1> ), .B(n1727), .Y(n2578) );
  OAI21X1 U611 ( .A(n1801), .B(n1725), .C(n2577), .Y(n2063) );
  NAND2X1 U612 ( .A(\mem<15><2> ), .B(n1727), .Y(n2577) );
  OAI21X1 U613 ( .A(n1799), .B(n1725), .C(n2576), .Y(n2062) );
  NAND2X1 U614 ( .A(\mem<15><3> ), .B(n1727), .Y(n2576) );
  OAI21X1 U615 ( .A(n1797), .B(n1725), .C(n2575), .Y(n2061) );
  NAND2X1 U616 ( .A(\mem<15><4> ), .B(n1727), .Y(n2575) );
  OAI21X1 U617 ( .A(n1795), .B(n1725), .C(n2574), .Y(n2060) );
  NAND2X1 U618 ( .A(\mem<15><5> ), .B(n1727), .Y(n2574) );
  OAI21X1 U619 ( .A(n1793), .B(n1725), .C(n2573), .Y(n2059) );
  NAND2X1 U620 ( .A(\mem<15><6> ), .B(n1727), .Y(n2573) );
  OAI21X1 U621 ( .A(n1791), .B(n1725), .C(n2572), .Y(n2058) );
  NAND2X1 U622 ( .A(\mem<15><7> ), .B(n1727), .Y(n2572) );
  OAI21X1 U623 ( .A(n1789), .B(n1725), .C(n2571), .Y(n2057) );
  NAND2X1 U624 ( .A(\mem<15><8> ), .B(n1726), .Y(n2571) );
  OAI21X1 U625 ( .A(n1788), .B(n1725), .C(n2570), .Y(n2056) );
  NAND2X1 U626 ( .A(\mem<15><9> ), .B(n1726), .Y(n2570) );
  OAI21X1 U627 ( .A(n1787), .B(n1725), .C(n2569), .Y(n2055) );
  NAND2X1 U628 ( .A(\mem<15><10> ), .B(n1726), .Y(n2569) );
  OAI21X1 U629 ( .A(n1785), .B(n1725), .C(n2568), .Y(n2054) );
  NAND2X1 U630 ( .A(\mem<15><11> ), .B(n1726), .Y(n2568) );
  OAI21X1 U631 ( .A(n1784), .B(n1725), .C(n2567), .Y(n2053) );
  NAND2X1 U632 ( .A(\mem<15><12> ), .B(n1726), .Y(n2567) );
  OAI21X1 U633 ( .A(n1783), .B(n1725), .C(n2566), .Y(n2052) );
  NAND2X1 U634 ( .A(\mem<15><13> ), .B(n1726), .Y(n2566) );
  OAI21X1 U635 ( .A(n1782), .B(n1725), .C(n2565), .Y(n2051) );
  NAND2X1 U636 ( .A(\mem<15><14> ), .B(n1726), .Y(n2565) );
  OAI21X1 U637 ( .A(n1780), .B(n1725), .C(n2564), .Y(n2050) );
  NAND2X1 U638 ( .A(\mem<15><15> ), .B(n1726), .Y(n2564) );
  OAI21X1 U641 ( .A(n1805), .B(n1722), .C(n2563), .Y(n2049) );
  NAND2X1 U642 ( .A(\mem<14><0> ), .B(n1724), .Y(n2563) );
  OAI21X1 U643 ( .A(n1803), .B(n1722), .C(n2562), .Y(n2048) );
  NAND2X1 U644 ( .A(\mem<14><1> ), .B(n1724), .Y(n2562) );
  OAI21X1 U645 ( .A(n1801), .B(n1722), .C(n2561), .Y(n2047) );
  NAND2X1 U646 ( .A(\mem<14><2> ), .B(n1724), .Y(n2561) );
  OAI21X1 U647 ( .A(n1799), .B(n1722), .C(n2560), .Y(n2046) );
  NAND2X1 U648 ( .A(\mem<14><3> ), .B(n1724), .Y(n2560) );
  OAI21X1 U649 ( .A(n1797), .B(n1722), .C(n2559), .Y(n2045) );
  NAND2X1 U650 ( .A(\mem<14><4> ), .B(n1724), .Y(n2559) );
  OAI21X1 U651 ( .A(n1795), .B(n1722), .C(n2558), .Y(n2044) );
  NAND2X1 U652 ( .A(\mem<14><5> ), .B(n1724), .Y(n2558) );
  OAI21X1 U653 ( .A(n1793), .B(n1722), .C(n2557), .Y(n2043) );
  NAND2X1 U654 ( .A(\mem<14><6> ), .B(n1724), .Y(n2557) );
  OAI21X1 U655 ( .A(n1791), .B(n1722), .C(n2556), .Y(n2042) );
  NAND2X1 U656 ( .A(\mem<14><7> ), .B(n1724), .Y(n2556) );
  OAI21X1 U657 ( .A(n1789), .B(n1722), .C(n2555), .Y(n2041) );
  NAND2X1 U658 ( .A(\mem<14><8> ), .B(n1723), .Y(n2555) );
  OAI21X1 U659 ( .A(n1788), .B(n1722), .C(n2554), .Y(n2040) );
  NAND2X1 U660 ( .A(\mem<14><9> ), .B(n1723), .Y(n2554) );
  OAI21X1 U661 ( .A(n1787), .B(n1722), .C(n2553), .Y(n2039) );
  NAND2X1 U662 ( .A(\mem<14><10> ), .B(n1723), .Y(n2553) );
  OAI21X1 U663 ( .A(n1785), .B(n1722), .C(n2552), .Y(n2038) );
  NAND2X1 U664 ( .A(\mem<14><11> ), .B(n1723), .Y(n2552) );
  OAI21X1 U665 ( .A(n1784), .B(n1722), .C(n2551), .Y(n2037) );
  NAND2X1 U666 ( .A(\mem<14><12> ), .B(n1723), .Y(n2551) );
  OAI21X1 U667 ( .A(n1783), .B(n1722), .C(n2550), .Y(n2036) );
  NAND2X1 U668 ( .A(\mem<14><13> ), .B(n1723), .Y(n2550) );
  OAI21X1 U669 ( .A(n1782), .B(n1722), .C(n2549), .Y(n2035) );
  NAND2X1 U670 ( .A(\mem<14><14> ), .B(n1723), .Y(n2549) );
  OAI21X1 U671 ( .A(n1780), .B(n1722), .C(n2548), .Y(n2034) );
  NAND2X1 U672 ( .A(\mem<14><15> ), .B(n1723), .Y(n2548) );
  OAI21X1 U675 ( .A(n1805), .B(n1719), .C(n2547), .Y(n2033) );
  NAND2X1 U676 ( .A(\mem<13><0> ), .B(n1721), .Y(n2547) );
  OAI21X1 U677 ( .A(n1803), .B(n1719), .C(n2546), .Y(n2032) );
  NAND2X1 U678 ( .A(\mem<13><1> ), .B(n1721), .Y(n2546) );
  OAI21X1 U679 ( .A(n1801), .B(n1719), .C(n2545), .Y(n2031) );
  NAND2X1 U680 ( .A(\mem<13><2> ), .B(n1721), .Y(n2545) );
  OAI21X1 U681 ( .A(n1799), .B(n1719), .C(n2544), .Y(n2030) );
  NAND2X1 U682 ( .A(\mem<13><3> ), .B(n1721), .Y(n2544) );
  OAI21X1 U683 ( .A(n1797), .B(n1719), .C(n2543), .Y(n2029) );
  NAND2X1 U684 ( .A(\mem<13><4> ), .B(n1721), .Y(n2543) );
  OAI21X1 U685 ( .A(n1795), .B(n1719), .C(n2542), .Y(n2028) );
  NAND2X1 U686 ( .A(\mem<13><5> ), .B(n1721), .Y(n2542) );
  OAI21X1 U687 ( .A(n1793), .B(n1719), .C(n2541), .Y(n2027) );
  NAND2X1 U688 ( .A(\mem<13><6> ), .B(n1721), .Y(n2541) );
  OAI21X1 U689 ( .A(n1791), .B(n1719), .C(n2540), .Y(n2026) );
  NAND2X1 U690 ( .A(\mem<13><7> ), .B(n1721), .Y(n2540) );
  OAI21X1 U691 ( .A(n1789), .B(n1719), .C(n2539), .Y(n2025) );
  NAND2X1 U692 ( .A(\mem<13><8> ), .B(n1720), .Y(n2539) );
  OAI21X1 U693 ( .A(n1788), .B(n1719), .C(n2538), .Y(n2024) );
  NAND2X1 U694 ( .A(\mem<13><9> ), .B(n1720), .Y(n2538) );
  OAI21X1 U695 ( .A(n1787), .B(n1719), .C(n2537), .Y(n2023) );
  NAND2X1 U696 ( .A(\mem<13><10> ), .B(n1720), .Y(n2537) );
  OAI21X1 U697 ( .A(n1785), .B(n1719), .C(n2536), .Y(n2022) );
  NAND2X1 U698 ( .A(\mem<13><11> ), .B(n1720), .Y(n2536) );
  OAI21X1 U699 ( .A(n1784), .B(n1719), .C(n2535), .Y(n2021) );
  NAND2X1 U700 ( .A(\mem<13><12> ), .B(n1720), .Y(n2535) );
  OAI21X1 U701 ( .A(n1783), .B(n1719), .C(n2534), .Y(n2020) );
  NAND2X1 U702 ( .A(\mem<13><13> ), .B(n1720), .Y(n2534) );
  OAI21X1 U703 ( .A(n1782), .B(n1719), .C(n2533), .Y(n2019) );
  NAND2X1 U704 ( .A(\mem<13><14> ), .B(n1720), .Y(n2533) );
  OAI21X1 U705 ( .A(n1780), .B(n1719), .C(n2532), .Y(n2018) );
  NAND2X1 U706 ( .A(\mem<13><15> ), .B(n1720), .Y(n2532) );
  OAI21X1 U709 ( .A(n1805), .B(n1716), .C(n2531), .Y(n2017) );
  NAND2X1 U710 ( .A(\mem<12><0> ), .B(n1718), .Y(n2531) );
  OAI21X1 U711 ( .A(n1803), .B(n1716), .C(n2530), .Y(n2016) );
  NAND2X1 U712 ( .A(\mem<12><1> ), .B(n1718), .Y(n2530) );
  OAI21X1 U713 ( .A(n1801), .B(n1716), .C(n2529), .Y(n2015) );
  NAND2X1 U714 ( .A(\mem<12><2> ), .B(n1718), .Y(n2529) );
  OAI21X1 U715 ( .A(n1799), .B(n1716), .C(n2528), .Y(n2014) );
  NAND2X1 U716 ( .A(\mem<12><3> ), .B(n1718), .Y(n2528) );
  OAI21X1 U717 ( .A(n1797), .B(n1716), .C(n2527), .Y(n2013) );
  NAND2X1 U718 ( .A(\mem<12><4> ), .B(n1718), .Y(n2527) );
  OAI21X1 U719 ( .A(n1795), .B(n1716), .C(n2526), .Y(n2012) );
  NAND2X1 U720 ( .A(\mem<12><5> ), .B(n1718), .Y(n2526) );
  OAI21X1 U721 ( .A(n1793), .B(n1716), .C(n2525), .Y(n2011) );
  NAND2X1 U722 ( .A(\mem<12><6> ), .B(n1718), .Y(n2525) );
  OAI21X1 U723 ( .A(n1791), .B(n1716), .C(n2524), .Y(n2010) );
  NAND2X1 U724 ( .A(\mem<12><7> ), .B(n1718), .Y(n2524) );
  OAI21X1 U725 ( .A(n1789), .B(n1716), .C(n2523), .Y(n2009) );
  NAND2X1 U726 ( .A(\mem<12><8> ), .B(n1717), .Y(n2523) );
  OAI21X1 U727 ( .A(n1788), .B(n1716), .C(n2522), .Y(n2008) );
  NAND2X1 U728 ( .A(\mem<12><9> ), .B(n1717), .Y(n2522) );
  OAI21X1 U729 ( .A(n1787), .B(n1716), .C(n2521), .Y(n2007) );
  NAND2X1 U730 ( .A(\mem<12><10> ), .B(n1717), .Y(n2521) );
  OAI21X1 U731 ( .A(n1785), .B(n1716), .C(n2520), .Y(n2006) );
  NAND2X1 U732 ( .A(\mem<12><11> ), .B(n1717), .Y(n2520) );
  OAI21X1 U733 ( .A(n1784), .B(n1716), .C(n2519), .Y(n2005) );
  NAND2X1 U734 ( .A(\mem<12><12> ), .B(n1717), .Y(n2519) );
  OAI21X1 U735 ( .A(n1783), .B(n1716), .C(n2518), .Y(n2004) );
  NAND2X1 U736 ( .A(\mem<12><13> ), .B(n1717), .Y(n2518) );
  OAI21X1 U737 ( .A(n1782), .B(n1716), .C(n2517), .Y(n2003) );
  NAND2X1 U738 ( .A(\mem<12><14> ), .B(n1717), .Y(n2517) );
  OAI21X1 U739 ( .A(n1780), .B(n1716), .C(n2516), .Y(n2002) );
  NAND2X1 U740 ( .A(\mem<12><15> ), .B(n1717), .Y(n2516) );
  OAI21X1 U743 ( .A(n1805), .B(n1713), .C(n2515), .Y(n2001) );
  NAND2X1 U744 ( .A(\mem<11><0> ), .B(n1715), .Y(n2515) );
  OAI21X1 U745 ( .A(n1803), .B(n1713), .C(n2514), .Y(n2000) );
  NAND2X1 U746 ( .A(\mem<11><1> ), .B(n1715), .Y(n2514) );
  OAI21X1 U747 ( .A(n1801), .B(n1713), .C(n2513), .Y(n1999) );
  NAND2X1 U748 ( .A(\mem<11><2> ), .B(n1715), .Y(n2513) );
  OAI21X1 U749 ( .A(n1799), .B(n1713), .C(n2512), .Y(n1998) );
  NAND2X1 U750 ( .A(\mem<11><3> ), .B(n1715), .Y(n2512) );
  OAI21X1 U751 ( .A(n1797), .B(n1713), .C(n2511), .Y(n1997) );
  NAND2X1 U752 ( .A(\mem<11><4> ), .B(n1715), .Y(n2511) );
  OAI21X1 U753 ( .A(n1795), .B(n1713), .C(n2510), .Y(n1996) );
  NAND2X1 U754 ( .A(\mem<11><5> ), .B(n1715), .Y(n2510) );
  OAI21X1 U755 ( .A(n1793), .B(n1713), .C(n2509), .Y(n1995) );
  NAND2X1 U756 ( .A(\mem<11><6> ), .B(n1715), .Y(n2509) );
  OAI21X1 U757 ( .A(n1791), .B(n1713), .C(n2508), .Y(n1994) );
  NAND2X1 U758 ( .A(\mem<11><7> ), .B(n1715), .Y(n2508) );
  OAI21X1 U759 ( .A(n1789), .B(n1713), .C(n2507), .Y(n1993) );
  NAND2X1 U760 ( .A(\mem<11><8> ), .B(n1714), .Y(n2507) );
  OAI21X1 U761 ( .A(n1788), .B(n1713), .C(n2506), .Y(n1992) );
  NAND2X1 U762 ( .A(\mem<11><9> ), .B(n1714), .Y(n2506) );
  OAI21X1 U763 ( .A(n1787), .B(n1713), .C(n2505), .Y(n1991) );
  NAND2X1 U764 ( .A(\mem<11><10> ), .B(n1714), .Y(n2505) );
  OAI21X1 U765 ( .A(n1785), .B(n1713), .C(n2504), .Y(n1990) );
  NAND2X1 U766 ( .A(\mem<11><11> ), .B(n1714), .Y(n2504) );
  OAI21X1 U767 ( .A(n1784), .B(n1713), .C(n2503), .Y(n1989) );
  NAND2X1 U768 ( .A(\mem<11><12> ), .B(n1714), .Y(n2503) );
  OAI21X1 U769 ( .A(n1783), .B(n1713), .C(n2502), .Y(n1988) );
  NAND2X1 U770 ( .A(\mem<11><13> ), .B(n1714), .Y(n2502) );
  OAI21X1 U771 ( .A(n1782), .B(n1713), .C(n2501), .Y(n1987) );
  NAND2X1 U772 ( .A(\mem<11><14> ), .B(n1714), .Y(n2501) );
  OAI21X1 U773 ( .A(n1780), .B(n1713), .C(n2500), .Y(n1986) );
  NAND2X1 U774 ( .A(\mem<11><15> ), .B(n1714), .Y(n2500) );
  OAI21X1 U777 ( .A(n1805), .B(n1710), .C(n2499), .Y(n1985) );
  NAND2X1 U778 ( .A(\mem<10><0> ), .B(n1712), .Y(n2499) );
  OAI21X1 U779 ( .A(n1803), .B(n1710), .C(n2498), .Y(n1984) );
  NAND2X1 U780 ( .A(\mem<10><1> ), .B(n1712), .Y(n2498) );
  OAI21X1 U781 ( .A(n1801), .B(n1710), .C(n2497), .Y(n1983) );
  NAND2X1 U782 ( .A(\mem<10><2> ), .B(n1712), .Y(n2497) );
  OAI21X1 U783 ( .A(n1799), .B(n1710), .C(n2496), .Y(n1982) );
  NAND2X1 U784 ( .A(\mem<10><3> ), .B(n1712), .Y(n2496) );
  OAI21X1 U785 ( .A(n1797), .B(n1710), .C(n2495), .Y(n1981) );
  NAND2X1 U786 ( .A(\mem<10><4> ), .B(n1712), .Y(n2495) );
  OAI21X1 U787 ( .A(n1795), .B(n1710), .C(n2494), .Y(n1980) );
  NAND2X1 U788 ( .A(\mem<10><5> ), .B(n1712), .Y(n2494) );
  OAI21X1 U789 ( .A(n1793), .B(n1710), .C(n2493), .Y(n1979) );
  NAND2X1 U790 ( .A(\mem<10><6> ), .B(n1712), .Y(n2493) );
  OAI21X1 U791 ( .A(n1791), .B(n1710), .C(n2492), .Y(n1978) );
  NAND2X1 U792 ( .A(\mem<10><7> ), .B(n1712), .Y(n2492) );
  OAI21X1 U793 ( .A(n1789), .B(n1710), .C(n2491), .Y(n1977) );
  NAND2X1 U794 ( .A(\mem<10><8> ), .B(n1711), .Y(n2491) );
  OAI21X1 U795 ( .A(n1788), .B(n1710), .C(n2490), .Y(n1976) );
  NAND2X1 U796 ( .A(\mem<10><9> ), .B(n1711), .Y(n2490) );
  OAI21X1 U797 ( .A(n1787), .B(n1710), .C(n2489), .Y(n1975) );
  NAND2X1 U798 ( .A(\mem<10><10> ), .B(n1711), .Y(n2489) );
  OAI21X1 U799 ( .A(n1785), .B(n1710), .C(n2488), .Y(n1974) );
  NAND2X1 U800 ( .A(\mem<10><11> ), .B(n1711), .Y(n2488) );
  OAI21X1 U801 ( .A(n1784), .B(n1710), .C(n2487), .Y(n1973) );
  NAND2X1 U802 ( .A(\mem<10><12> ), .B(n1711), .Y(n2487) );
  OAI21X1 U803 ( .A(n1783), .B(n1710), .C(n2486), .Y(n1972) );
  NAND2X1 U804 ( .A(\mem<10><13> ), .B(n1711), .Y(n2486) );
  OAI21X1 U805 ( .A(n1782), .B(n1710), .C(n2485), .Y(n1971) );
  NAND2X1 U806 ( .A(\mem<10><14> ), .B(n1711), .Y(n2485) );
  OAI21X1 U807 ( .A(n1780), .B(n1710), .C(n2484), .Y(n1970) );
  NAND2X1 U808 ( .A(\mem<10><15> ), .B(n1711), .Y(n2484) );
  OAI21X1 U811 ( .A(n1805), .B(n1707), .C(n2483), .Y(n1969) );
  NAND2X1 U812 ( .A(\mem<9><0> ), .B(n1709), .Y(n2483) );
  OAI21X1 U813 ( .A(n1803), .B(n1707), .C(n2482), .Y(n1968) );
  NAND2X1 U814 ( .A(\mem<9><1> ), .B(n1709), .Y(n2482) );
  OAI21X1 U815 ( .A(n1801), .B(n1707), .C(n2481), .Y(n1967) );
  NAND2X1 U816 ( .A(\mem<9><2> ), .B(n1709), .Y(n2481) );
  OAI21X1 U817 ( .A(n1799), .B(n1707), .C(n2480), .Y(n1966) );
  NAND2X1 U818 ( .A(\mem<9><3> ), .B(n1709), .Y(n2480) );
  OAI21X1 U819 ( .A(n1797), .B(n1707), .C(n2479), .Y(n1965) );
  NAND2X1 U820 ( .A(\mem<9><4> ), .B(n1709), .Y(n2479) );
  OAI21X1 U821 ( .A(n1795), .B(n1707), .C(n2478), .Y(n1964) );
  NAND2X1 U822 ( .A(\mem<9><5> ), .B(n1709), .Y(n2478) );
  OAI21X1 U823 ( .A(n1793), .B(n1707), .C(n2477), .Y(n1963) );
  NAND2X1 U824 ( .A(\mem<9><6> ), .B(n1709), .Y(n2477) );
  OAI21X1 U825 ( .A(n1791), .B(n1707), .C(n2476), .Y(n1962) );
  NAND2X1 U826 ( .A(\mem<9><7> ), .B(n1709), .Y(n2476) );
  OAI21X1 U827 ( .A(n1789), .B(n1707), .C(n2475), .Y(n1961) );
  NAND2X1 U828 ( .A(\mem<9><8> ), .B(n1708), .Y(n2475) );
  OAI21X1 U829 ( .A(n1788), .B(n1707), .C(n2474), .Y(n1960) );
  NAND2X1 U830 ( .A(\mem<9><9> ), .B(n1708), .Y(n2474) );
  OAI21X1 U831 ( .A(n1787), .B(n1707), .C(n2473), .Y(n1959) );
  NAND2X1 U832 ( .A(\mem<9><10> ), .B(n1708), .Y(n2473) );
  OAI21X1 U833 ( .A(n1785), .B(n1707), .C(n2472), .Y(n1958) );
  NAND2X1 U834 ( .A(\mem<9><11> ), .B(n1708), .Y(n2472) );
  OAI21X1 U835 ( .A(n1784), .B(n1707), .C(n2471), .Y(n1957) );
  NAND2X1 U836 ( .A(\mem<9><12> ), .B(n1708), .Y(n2471) );
  OAI21X1 U837 ( .A(n1783), .B(n1707), .C(n2470), .Y(n1956) );
  NAND2X1 U838 ( .A(\mem<9><13> ), .B(n1708), .Y(n2470) );
  OAI21X1 U839 ( .A(n1782), .B(n1707), .C(n2469), .Y(n1955) );
  NAND2X1 U840 ( .A(\mem<9><14> ), .B(n1708), .Y(n2469) );
  OAI21X1 U841 ( .A(n1780), .B(n1707), .C(n2468), .Y(n1954) );
  NAND2X1 U842 ( .A(\mem<9><15> ), .B(n1708), .Y(n2468) );
  OAI21X1 U845 ( .A(n1805), .B(n1704), .C(n2467), .Y(n1953) );
  NAND2X1 U846 ( .A(\mem<8><0> ), .B(n1706), .Y(n2467) );
  OAI21X1 U847 ( .A(n1803), .B(n1704), .C(n2466), .Y(n1952) );
  NAND2X1 U848 ( .A(\mem<8><1> ), .B(n1706), .Y(n2466) );
  OAI21X1 U849 ( .A(n1801), .B(n1704), .C(n2465), .Y(n1951) );
  NAND2X1 U850 ( .A(\mem<8><2> ), .B(n1706), .Y(n2465) );
  OAI21X1 U851 ( .A(n1799), .B(n1704), .C(n2464), .Y(n1950) );
  NAND2X1 U852 ( .A(\mem<8><3> ), .B(n1706), .Y(n2464) );
  OAI21X1 U853 ( .A(n1797), .B(n1704), .C(n2463), .Y(n1949) );
  NAND2X1 U854 ( .A(\mem<8><4> ), .B(n1706), .Y(n2463) );
  OAI21X1 U855 ( .A(n1795), .B(n1704), .C(n2462), .Y(n1948) );
  NAND2X1 U856 ( .A(\mem<8><5> ), .B(n1706), .Y(n2462) );
  OAI21X1 U857 ( .A(n1793), .B(n1704), .C(n2461), .Y(n1947) );
  NAND2X1 U858 ( .A(\mem<8><6> ), .B(n1706), .Y(n2461) );
  OAI21X1 U859 ( .A(n1791), .B(n1704), .C(n2460), .Y(n1946) );
  NAND2X1 U860 ( .A(\mem<8><7> ), .B(n1706), .Y(n2460) );
  OAI21X1 U861 ( .A(n1789), .B(n1704), .C(n2459), .Y(n1945) );
  NAND2X1 U862 ( .A(\mem<8><8> ), .B(n1705), .Y(n2459) );
  OAI21X1 U863 ( .A(n1788), .B(n1704), .C(n2458), .Y(n1944) );
  NAND2X1 U864 ( .A(\mem<8><9> ), .B(n1705), .Y(n2458) );
  OAI21X1 U865 ( .A(n1787), .B(n1704), .C(n2457), .Y(n1943) );
  NAND2X1 U866 ( .A(\mem<8><10> ), .B(n1705), .Y(n2457) );
  OAI21X1 U867 ( .A(n1785), .B(n1704), .C(n2456), .Y(n1942) );
  NAND2X1 U868 ( .A(\mem<8><11> ), .B(n1705), .Y(n2456) );
  OAI21X1 U869 ( .A(n1784), .B(n1704), .C(n2455), .Y(n1941) );
  NAND2X1 U870 ( .A(\mem<8><12> ), .B(n1705), .Y(n2455) );
  OAI21X1 U871 ( .A(n1783), .B(n1704), .C(n2454), .Y(n1940) );
  NAND2X1 U872 ( .A(\mem<8><13> ), .B(n1705), .Y(n2454) );
  OAI21X1 U873 ( .A(n1782), .B(n1704), .C(n2453), .Y(n1939) );
  NAND2X1 U874 ( .A(\mem<8><14> ), .B(n1705), .Y(n2453) );
  OAI21X1 U875 ( .A(n1780), .B(n1704), .C(n2452), .Y(n1938) );
  NAND2X1 U876 ( .A(\mem<8><15> ), .B(n1705), .Y(n2452) );
  NAND3X1 U879 ( .A(n2709), .B(net59340), .C(net59458), .Y(n2451) );
  OAI21X1 U880 ( .A(n1805), .B(n1701), .C(n2450), .Y(n1937) );
  NAND2X1 U881 ( .A(\mem<7><0> ), .B(n1703), .Y(n2450) );
  OAI21X1 U882 ( .A(n1803), .B(n1701), .C(n2449), .Y(n1936) );
  NAND2X1 U883 ( .A(\mem<7><1> ), .B(n1703), .Y(n2449) );
  OAI21X1 U884 ( .A(n1801), .B(n1701), .C(n2448), .Y(n1935) );
  NAND2X1 U885 ( .A(\mem<7><2> ), .B(n1703), .Y(n2448) );
  OAI21X1 U886 ( .A(n1799), .B(n1701), .C(n2447), .Y(n1934) );
  NAND2X1 U887 ( .A(\mem<7><3> ), .B(n1703), .Y(n2447) );
  OAI21X1 U888 ( .A(n1797), .B(n1701), .C(n2446), .Y(n1933) );
  NAND2X1 U889 ( .A(\mem<7><4> ), .B(n1703), .Y(n2446) );
  OAI21X1 U890 ( .A(n1795), .B(n1701), .C(n2445), .Y(n1932) );
  NAND2X1 U891 ( .A(\mem<7><5> ), .B(n1703), .Y(n2445) );
  OAI21X1 U892 ( .A(n1793), .B(n1701), .C(n2444), .Y(n1931) );
  NAND2X1 U893 ( .A(\mem<7><6> ), .B(n1703), .Y(n2444) );
  OAI21X1 U894 ( .A(n1791), .B(n1701), .C(n2443), .Y(n1930) );
  NAND2X1 U895 ( .A(\mem<7><7> ), .B(n1703), .Y(n2443) );
  OAI21X1 U896 ( .A(n1789), .B(n1701), .C(n2442), .Y(n1929) );
  NAND2X1 U897 ( .A(\mem<7><8> ), .B(n1702), .Y(n2442) );
  OAI21X1 U898 ( .A(n1788), .B(n1701), .C(n2441), .Y(n1928) );
  NAND2X1 U899 ( .A(\mem<7><9> ), .B(n1702), .Y(n2441) );
  OAI21X1 U900 ( .A(n1787), .B(n1701), .C(n2440), .Y(n1927) );
  NAND2X1 U901 ( .A(\mem<7><10> ), .B(n1702), .Y(n2440) );
  OAI21X1 U902 ( .A(n1785), .B(n1701), .C(n2439), .Y(n1926) );
  NAND2X1 U903 ( .A(\mem<7><11> ), .B(n1702), .Y(n2439) );
  OAI21X1 U904 ( .A(n1784), .B(n1701), .C(n2438), .Y(n1925) );
  NAND2X1 U905 ( .A(\mem<7><12> ), .B(n1702), .Y(n2438) );
  OAI21X1 U906 ( .A(n1783), .B(n1701), .C(n2437), .Y(n1924) );
  NAND2X1 U907 ( .A(\mem<7><13> ), .B(n1702), .Y(n2437) );
  OAI21X1 U908 ( .A(n1782), .B(n1701), .C(n2436), .Y(n1923) );
  NAND2X1 U909 ( .A(\mem<7><14> ), .B(n1702), .Y(n2436) );
  OAI21X1 U910 ( .A(n1780), .B(n1701), .C(n2435), .Y(n1922) );
  NAND2X1 U911 ( .A(\mem<7><15> ), .B(n1702), .Y(n2435) );
  NOR3X1 U914 ( .A(net60096), .B(net60828), .C(net59640), .Y(n2830) );
  OAI21X1 U915 ( .A(n1805), .B(n1698), .C(n2434), .Y(n1921) );
  NAND2X1 U916 ( .A(\mem<6><0> ), .B(n1700), .Y(n2434) );
  OAI21X1 U917 ( .A(n1803), .B(n1698), .C(n2433), .Y(n1920) );
  NAND2X1 U918 ( .A(\mem<6><1> ), .B(n1700), .Y(n2433) );
  OAI21X1 U919 ( .A(n1801), .B(n1698), .C(n2432), .Y(n1919) );
  NAND2X1 U920 ( .A(\mem<6><2> ), .B(n1700), .Y(n2432) );
  OAI21X1 U921 ( .A(n1799), .B(n1698), .C(n2431), .Y(n1918) );
  NAND2X1 U922 ( .A(\mem<6><3> ), .B(n1700), .Y(n2431) );
  OAI21X1 U923 ( .A(n1797), .B(n1698), .C(n2430), .Y(n1917) );
  NAND2X1 U924 ( .A(\mem<6><4> ), .B(n1700), .Y(n2430) );
  OAI21X1 U925 ( .A(n1795), .B(n1698), .C(n2429), .Y(n1916) );
  NAND2X1 U926 ( .A(\mem<6><5> ), .B(n1700), .Y(n2429) );
  OAI21X1 U927 ( .A(n1793), .B(n1698), .C(n2428), .Y(n1915) );
  NAND2X1 U928 ( .A(\mem<6><6> ), .B(n1700), .Y(n2428) );
  OAI21X1 U929 ( .A(n1791), .B(n1698), .C(n2427), .Y(n1914) );
  NAND2X1 U930 ( .A(\mem<6><7> ), .B(n1700), .Y(n2427) );
  OAI21X1 U931 ( .A(n1789), .B(n1698), .C(n2426), .Y(n1913) );
  NAND2X1 U932 ( .A(\mem<6><8> ), .B(n1699), .Y(n2426) );
  OAI21X1 U933 ( .A(n1788), .B(n1698), .C(n2425), .Y(n1912) );
  NAND2X1 U934 ( .A(\mem<6><9> ), .B(n1699), .Y(n2425) );
  OAI21X1 U935 ( .A(n1787), .B(n1698), .C(n2424), .Y(n1911) );
  NAND2X1 U936 ( .A(\mem<6><10> ), .B(n1699), .Y(n2424) );
  OAI21X1 U937 ( .A(n1785), .B(n1698), .C(n2423), .Y(n1910) );
  NAND2X1 U938 ( .A(\mem<6><11> ), .B(n1699), .Y(n2423) );
  OAI21X1 U939 ( .A(n1784), .B(n1698), .C(n2422), .Y(n1909) );
  NAND2X1 U940 ( .A(\mem<6><12> ), .B(n1699), .Y(n2422) );
  OAI21X1 U941 ( .A(n1783), .B(n1698), .C(n2421), .Y(n1908) );
  NAND2X1 U942 ( .A(\mem<6><13> ), .B(n1699), .Y(n2421) );
  OAI21X1 U943 ( .A(n1782), .B(n1698), .C(n2420), .Y(n1907) );
  NAND2X1 U944 ( .A(\mem<6><14> ), .B(n1699), .Y(n2420) );
  OAI21X1 U945 ( .A(n1780), .B(n1698), .C(n2419), .Y(n1906) );
  NAND2X1 U946 ( .A(\mem<6><15> ), .B(n1699), .Y(n2419) );
  NOR3X1 U949 ( .A(net60096), .B(net60826), .C(net59640), .Y(n2813) );
  OAI21X1 U950 ( .A(n1804), .B(n1695), .C(n2418), .Y(n1905) );
  NAND2X1 U951 ( .A(\mem<5><0> ), .B(n1697), .Y(n2418) );
  OAI21X1 U952 ( .A(n1802), .B(n1695), .C(n2417), .Y(n1904) );
  NAND2X1 U953 ( .A(\mem<5><1> ), .B(n1697), .Y(n2417) );
  OAI21X1 U954 ( .A(n1800), .B(n1695), .C(n2416), .Y(n1903) );
  NAND2X1 U955 ( .A(\mem<5><2> ), .B(n1697), .Y(n2416) );
  OAI21X1 U956 ( .A(n1798), .B(n1695), .C(n2415), .Y(n1902) );
  NAND2X1 U957 ( .A(\mem<5><3> ), .B(n1697), .Y(n2415) );
  OAI21X1 U958 ( .A(n1796), .B(n1695), .C(n2414), .Y(n1901) );
  NAND2X1 U959 ( .A(\mem<5><4> ), .B(n1697), .Y(n2414) );
  OAI21X1 U960 ( .A(n1794), .B(n1695), .C(n2413), .Y(n1900) );
  NAND2X1 U961 ( .A(\mem<5><5> ), .B(n1697), .Y(n2413) );
  OAI21X1 U962 ( .A(n1792), .B(n1695), .C(n2412), .Y(n1899) );
  NAND2X1 U963 ( .A(\mem<5><6> ), .B(n1697), .Y(n2412) );
  OAI21X1 U964 ( .A(n1790), .B(n1695), .C(n2411), .Y(n1898) );
  NAND2X1 U965 ( .A(\mem<5><7> ), .B(n1697), .Y(n2411) );
  OAI21X1 U966 ( .A(n1789), .B(n1695), .C(n2410), .Y(n1897) );
  NAND2X1 U967 ( .A(\mem<5><8> ), .B(n1696), .Y(n2410) );
  OAI21X1 U968 ( .A(n1788), .B(n1695), .C(n2409), .Y(n1896) );
  NAND2X1 U969 ( .A(\mem<5><9> ), .B(n1696), .Y(n2409) );
  OAI21X1 U970 ( .A(n1786), .B(n1695), .C(n2408), .Y(n1895) );
  NAND2X1 U971 ( .A(\mem<5><10> ), .B(n1696), .Y(n2408) );
  OAI21X1 U972 ( .A(n1785), .B(n1695), .C(n2407), .Y(n1894) );
  NAND2X1 U973 ( .A(\mem<5><11> ), .B(n1696), .Y(n2407) );
  OAI21X1 U974 ( .A(n1784), .B(n1695), .C(n2406), .Y(n1893) );
  NAND2X1 U975 ( .A(\mem<5><12> ), .B(n1696), .Y(n2406) );
  OAI21X1 U976 ( .A(n1783), .B(n1695), .C(n2405), .Y(n1892) );
  NAND2X1 U977 ( .A(\mem<5><13> ), .B(n1696), .Y(n2405) );
  OAI21X1 U978 ( .A(n1781), .B(n1695), .C(n2404), .Y(n1891) );
  NAND2X1 U979 ( .A(\mem<5><14> ), .B(n1696), .Y(n2404) );
  OAI21X1 U980 ( .A(n1780), .B(n1695), .C(n2403), .Y(n1890) );
  NAND2X1 U981 ( .A(\mem<5><15> ), .B(n1696), .Y(n2403) );
  NOR3X1 U984 ( .A(net60828), .B(net60094), .C(net59640), .Y(n2796) );
  OAI21X1 U985 ( .A(n1805), .B(n1692), .C(n2402), .Y(n1889) );
  NAND2X1 U986 ( .A(\mem<4><0> ), .B(n1694), .Y(n2402) );
  OAI21X1 U987 ( .A(n1803), .B(n1692), .C(n2401), .Y(n1888) );
  NAND2X1 U988 ( .A(\mem<4><1> ), .B(n1694), .Y(n2401) );
  OAI21X1 U989 ( .A(n1801), .B(n1692), .C(n2400), .Y(n1887) );
  NAND2X1 U990 ( .A(\mem<4><2> ), .B(n1694), .Y(n2400) );
  OAI21X1 U991 ( .A(n1799), .B(n1692), .C(n2399), .Y(n1886) );
  NAND2X1 U992 ( .A(\mem<4><3> ), .B(n1694), .Y(n2399) );
  OAI21X1 U993 ( .A(n1797), .B(n1692), .C(n2398), .Y(n1885) );
  NAND2X1 U994 ( .A(\mem<4><4> ), .B(n1694), .Y(n2398) );
  OAI21X1 U995 ( .A(n1795), .B(n1692), .C(n2397), .Y(n1884) );
  NAND2X1 U996 ( .A(\mem<4><5> ), .B(n1694), .Y(n2397) );
  OAI21X1 U997 ( .A(n1793), .B(n1692), .C(n2396), .Y(n1883) );
  NAND2X1 U998 ( .A(\mem<4><6> ), .B(n1694), .Y(n2396) );
  OAI21X1 U999 ( .A(n1791), .B(n1692), .C(n2395), .Y(n1882) );
  NAND2X1 U1000 ( .A(\mem<4><7> ), .B(n1694), .Y(n2395) );
  OAI21X1 U1001 ( .A(n1789), .B(n1692), .C(n2394), .Y(n1881) );
  NAND2X1 U1002 ( .A(\mem<4><8> ), .B(n1693), .Y(n2394) );
  OAI21X1 U1003 ( .A(n1788), .B(n1692), .C(n2393), .Y(n1880) );
  NAND2X1 U1004 ( .A(\mem<4><9> ), .B(n1693), .Y(n2393) );
  OAI21X1 U1005 ( .A(n1787), .B(n1692), .C(n2392), .Y(n1879) );
  NAND2X1 U1006 ( .A(\mem<4><10> ), .B(n1693), .Y(n2392) );
  OAI21X1 U1007 ( .A(n1785), .B(n1692), .C(n2391), .Y(n1878) );
  NAND2X1 U1008 ( .A(\mem<4><11> ), .B(n1693), .Y(n2391) );
  OAI21X1 U1009 ( .A(n1784), .B(n1692), .C(n2390), .Y(n1877) );
  NAND2X1 U1010 ( .A(\mem<4><12> ), .B(n1693), .Y(n2390) );
  OAI21X1 U1011 ( .A(n1783), .B(n1692), .C(n2389), .Y(n1876) );
  NAND2X1 U1012 ( .A(\mem<4><13> ), .B(n1693), .Y(n2389) );
  OAI21X1 U1013 ( .A(n1782), .B(n1692), .C(n2388), .Y(n1875) );
  NAND2X1 U1014 ( .A(\mem<4><14> ), .B(n1693), .Y(n2388) );
  OAI21X1 U1015 ( .A(n1780), .B(n1692), .C(n2387), .Y(n1874) );
  NAND2X1 U1016 ( .A(\mem<4><15> ), .B(n1693), .Y(n2387) );
  NOR3X1 U1019 ( .A(net60826), .B(net60094), .C(net59640), .Y(n2779) );
  OAI21X1 U1020 ( .A(n1804), .B(n1689), .C(n2386), .Y(n1873) );
  NAND2X1 U1021 ( .A(\mem<3><0> ), .B(n1691), .Y(n2386) );
  OAI21X1 U1022 ( .A(n1802), .B(n1689), .C(n2385), .Y(n1872) );
  NAND2X1 U1023 ( .A(\mem<3><1> ), .B(n1691), .Y(n2385) );
  OAI21X1 U1024 ( .A(n1800), .B(n1689), .C(n2384), .Y(n1871) );
  NAND2X1 U1025 ( .A(\mem<3><2> ), .B(n1691), .Y(n2384) );
  OAI21X1 U1026 ( .A(n1798), .B(n1689), .C(n2383), .Y(n1870) );
  NAND2X1 U1027 ( .A(\mem<3><3> ), .B(n1691), .Y(n2383) );
  OAI21X1 U1028 ( .A(n1796), .B(n1689), .C(n2382), .Y(n1869) );
  NAND2X1 U1029 ( .A(\mem<3><4> ), .B(n1691), .Y(n2382) );
  OAI21X1 U1030 ( .A(n1794), .B(n1689), .C(n2381), .Y(n1868) );
  NAND2X1 U1031 ( .A(\mem<3><5> ), .B(n1691), .Y(n2381) );
  OAI21X1 U1032 ( .A(n1792), .B(n1689), .C(n2380), .Y(n1867) );
  NAND2X1 U1033 ( .A(\mem<3><6> ), .B(n1691), .Y(n2380) );
  OAI21X1 U1034 ( .A(n1790), .B(n1689), .C(n2379), .Y(n1866) );
  NAND2X1 U1035 ( .A(\mem<3><7> ), .B(n1691), .Y(n2379) );
  OAI21X1 U1036 ( .A(n1789), .B(n1689), .C(n2378), .Y(n1865) );
  NAND2X1 U1037 ( .A(\mem<3><8> ), .B(n1690), .Y(n2378) );
  OAI21X1 U1038 ( .A(n1788), .B(n1689), .C(n2377), .Y(n1864) );
  NAND2X1 U1039 ( .A(\mem<3><9> ), .B(n1690), .Y(n2377) );
  OAI21X1 U1040 ( .A(n1786), .B(n1689), .C(n2376), .Y(n1863) );
  NAND2X1 U1041 ( .A(\mem<3><10> ), .B(n1690), .Y(n2376) );
  OAI21X1 U1042 ( .A(n1785), .B(n1689), .C(n2375), .Y(n1862) );
  NAND2X1 U1043 ( .A(\mem<3><11> ), .B(n1690), .Y(n2375) );
  OAI21X1 U1044 ( .A(n1784), .B(n1689), .C(n2374), .Y(n1861) );
  NAND2X1 U1045 ( .A(\mem<3><12> ), .B(n1690), .Y(n2374) );
  OAI21X1 U1046 ( .A(n1783), .B(n1689), .C(n2373), .Y(n1860) );
  NAND2X1 U1047 ( .A(\mem<3><13> ), .B(n1690), .Y(n2373) );
  OAI21X1 U1048 ( .A(n1781), .B(n1689), .C(n2372), .Y(n1859) );
  NAND2X1 U1049 ( .A(\mem<3><14> ), .B(n1690), .Y(n2372) );
  OAI21X1 U1050 ( .A(n1780), .B(n1689), .C(n2371), .Y(n1858) );
  NAND2X1 U1051 ( .A(\mem<3><15> ), .B(n1690), .Y(n2371) );
  NOR3X1 U1054 ( .A(net60828), .B(net59638), .C(net60096), .Y(n2762) );
  OAI21X1 U1055 ( .A(n1805), .B(n1686), .C(n2370), .Y(n1857) );
  NAND2X1 U1056 ( .A(\mem<2><0> ), .B(n1688), .Y(n2370) );
  OAI21X1 U1057 ( .A(n1803), .B(n1686), .C(n2369), .Y(n1856) );
  NAND2X1 U1058 ( .A(\mem<2><1> ), .B(n1688), .Y(n2369) );
  OAI21X1 U1059 ( .A(n1801), .B(n1686), .C(n2368), .Y(n1855) );
  NAND2X1 U1060 ( .A(\mem<2><2> ), .B(n1688), .Y(n2368) );
  OAI21X1 U1061 ( .A(n1799), .B(n1686), .C(n2367), .Y(n1854) );
  NAND2X1 U1062 ( .A(\mem<2><3> ), .B(n1688), .Y(n2367) );
  OAI21X1 U1063 ( .A(n1797), .B(n1686), .C(n2366), .Y(n1853) );
  NAND2X1 U1064 ( .A(\mem<2><4> ), .B(n1688), .Y(n2366) );
  OAI21X1 U1065 ( .A(n1795), .B(n1686), .C(n2365), .Y(n1852) );
  NAND2X1 U1066 ( .A(\mem<2><5> ), .B(n1688), .Y(n2365) );
  OAI21X1 U1067 ( .A(n1793), .B(n1686), .C(n2364), .Y(n1851) );
  NAND2X1 U1068 ( .A(\mem<2><6> ), .B(n1688), .Y(n2364) );
  OAI21X1 U1069 ( .A(n1791), .B(n1686), .C(n2363), .Y(n1850) );
  NAND2X1 U1070 ( .A(\mem<2><7> ), .B(n1688), .Y(n2363) );
  OAI21X1 U1071 ( .A(n1789), .B(n1686), .C(n2362), .Y(n1849) );
  NAND2X1 U1072 ( .A(\mem<2><8> ), .B(n1687), .Y(n2362) );
  OAI21X1 U1073 ( .A(n1788), .B(n1686), .C(n2361), .Y(n1848) );
  NAND2X1 U1074 ( .A(\mem<2><9> ), .B(n1687), .Y(n2361) );
  OAI21X1 U1075 ( .A(n1787), .B(n1686), .C(n2360), .Y(n1847) );
  NAND2X1 U1076 ( .A(\mem<2><10> ), .B(n1687), .Y(n2360) );
  OAI21X1 U1077 ( .A(n1785), .B(n1686), .C(n2359), .Y(n1846) );
  NAND2X1 U1078 ( .A(\mem<2><11> ), .B(n1687), .Y(n2359) );
  OAI21X1 U1079 ( .A(n1784), .B(n1686), .C(n2358), .Y(n1845) );
  NAND2X1 U1080 ( .A(\mem<2><12> ), .B(n1687), .Y(n2358) );
  OAI21X1 U1081 ( .A(n1783), .B(n1686), .C(n2357), .Y(n1844) );
  NAND2X1 U1082 ( .A(\mem<2><13> ), .B(n1687), .Y(n2357) );
  OAI21X1 U1083 ( .A(n1782), .B(n1686), .C(n2356), .Y(n1843) );
  NAND2X1 U1084 ( .A(\mem<2><14> ), .B(n1687), .Y(n2356) );
  OAI21X1 U1085 ( .A(n1780), .B(n1686), .C(n2355), .Y(n1842) );
  NAND2X1 U1086 ( .A(\mem<2><15> ), .B(n1687), .Y(n2355) );
  NOR3X1 U1089 ( .A(net60826), .B(net59638), .C(net60096), .Y(n2745) );
  OAI21X1 U1090 ( .A(n1804), .B(n1683), .C(n2354), .Y(n1841) );
  NAND2X1 U1091 ( .A(\mem<1><0> ), .B(n1685), .Y(n2354) );
  OAI21X1 U1092 ( .A(n1802), .B(n1683), .C(n2353), .Y(n1840) );
  NAND2X1 U1093 ( .A(\mem<1><1> ), .B(n1685), .Y(n2353) );
  OAI21X1 U1094 ( .A(n1800), .B(n1683), .C(n2352), .Y(n1839) );
  NAND2X1 U1095 ( .A(\mem<1><2> ), .B(n1685), .Y(n2352) );
  OAI21X1 U1096 ( .A(n1798), .B(n1683), .C(n2351), .Y(n1838) );
  NAND2X1 U1097 ( .A(\mem<1><3> ), .B(n1685), .Y(n2351) );
  OAI21X1 U1098 ( .A(n1796), .B(n1683), .C(n2350), .Y(n1837) );
  NAND2X1 U1099 ( .A(\mem<1><4> ), .B(n1685), .Y(n2350) );
  OAI21X1 U1100 ( .A(n1794), .B(n1683), .C(n2349), .Y(n1836) );
  NAND2X1 U1101 ( .A(\mem<1><5> ), .B(n1685), .Y(n2349) );
  OAI21X1 U1102 ( .A(n1792), .B(n1683), .C(n2348), .Y(n1835) );
  NAND2X1 U1103 ( .A(\mem<1><6> ), .B(n1685), .Y(n2348) );
  OAI21X1 U1104 ( .A(n1790), .B(n1683), .C(n2347), .Y(n1834) );
  NAND2X1 U1105 ( .A(\mem<1><7> ), .B(n1685), .Y(n2347) );
  OAI21X1 U1106 ( .A(n1789), .B(n1683), .C(n2346), .Y(n1833) );
  NAND2X1 U1107 ( .A(\mem<1><8> ), .B(n1684), .Y(n2346) );
  OAI21X1 U1108 ( .A(n1788), .B(n1683), .C(n2345), .Y(n1832) );
  NAND2X1 U1109 ( .A(\mem<1><9> ), .B(n1684), .Y(n2345) );
  OAI21X1 U1110 ( .A(n1786), .B(n1683), .C(n2344), .Y(n1831) );
  NAND2X1 U1111 ( .A(\mem<1><10> ), .B(n1684), .Y(n2344) );
  OAI21X1 U1112 ( .A(n1785), .B(n1683), .C(n2343), .Y(n1830) );
  NAND2X1 U1113 ( .A(\mem<1><11> ), .B(n1684), .Y(n2343) );
  OAI21X1 U1114 ( .A(n1784), .B(n1683), .C(n2342), .Y(n1829) );
  NAND2X1 U1115 ( .A(\mem<1><12> ), .B(n1684), .Y(n2342) );
  OAI21X1 U1116 ( .A(n1783), .B(n1683), .C(n2341), .Y(n1828) );
  NAND2X1 U1117 ( .A(\mem<1><13> ), .B(n1684), .Y(n2341) );
  OAI21X1 U1118 ( .A(n1781), .B(n1683), .C(n2340), .Y(n1827) );
  NAND2X1 U1119 ( .A(\mem<1><14> ), .B(n1684), .Y(n2340) );
  OAI21X1 U1120 ( .A(n1780), .B(n1683), .C(n2339), .Y(n1826) );
  NAND2X1 U1121 ( .A(\mem<1><15> ), .B(n1684), .Y(n2339) );
  NOR3X1 U1124 ( .A(net60094), .B(net59638), .C(net60828), .Y(n2728) );
  OAI21X1 U1125 ( .A(n1805), .B(n1680), .C(n2338), .Y(n1825) );
  NAND2X1 U1126 ( .A(\mem<0><0> ), .B(n1682), .Y(n2338) );
  OAI21X1 U1128 ( .A(n1803), .B(n1680), .C(n2337), .Y(n1824) );
  NAND2X1 U1129 ( .A(\mem<0><1> ), .B(n1682), .Y(n2337) );
  OAI21X1 U1131 ( .A(n1801), .B(n1680), .C(n2336), .Y(n1823) );
  NAND2X1 U1132 ( .A(\mem<0><2> ), .B(n1682), .Y(n2336) );
  OAI21X1 U1134 ( .A(n1799), .B(n1680), .C(n2335), .Y(n1822) );
  NAND2X1 U1135 ( .A(\mem<0><3> ), .B(n1682), .Y(n2335) );
  OAI21X1 U1137 ( .A(n1797), .B(n1680), .C(n2334), .Y(n1821) );
  NAND2X1 U1138 ( .A(\mem<0><4> ), .B(n1682), .Y(n2334) );
  OAI21X1 U1140 ( .A(n1795), .B(n1680), .C(n2333), .Y(n1820) );
  NAND2X1 U1141 ( .A(\mem<0><5> ), .B(n1682), .Y(n2333) );
  OAI21X1 U1143 ( .A(n1793), .B(n1680), .C(n2332), .Y(n1819) );
  NAND2X1 U1144 ( .A(\mem<0><6> ), .B(n1682), .Y(n2332) );
  OAI21X1 U1146 ( .A(n1791), .B(n1680), .C(n2331), .Y(n1818) );
  NAND2X1 U1147 ( .A(\mem<0><7> ), .B(n1682), .Y(n2331) );
  OAI21X1 U1149 ( .A(n1789), .B(n1680), .C(n2330), .Y(n1817) );
  NAND2X1 U1150 ( .A(\mem<0><8> ), .B(n1681), .Y(n2330) );
  OAI21X1 U1152 ( .A(n1788), .B(n1680), .C(n2329), .Y(n1816) );
  NAND2X1 U1153 ( .A(\mem<0><9> ), .B(n1681), .Y(n2329) );
  OAI21X1 U1155 ( .A(n1787), .B(n1680), .C(n2328), .Y(n1815) );
  NAND2X1 U1156 ( .A(\mem<0><10> ), .B(n1681), .Y(n2328) );
  OAI21X1 U1158 ( .A(n1785), .B(n1680), .C(n2327), .Y(n1814) );
  NAND2X1 U1159 ( .A(\mem<0><11> ), .B(n1681), .Y(n2327) );
  OAI21X1 U1161 ( .A(n1784), .B(n1680), .C(n2326), .Y(n1813) );
  NAND2X1 U1162 ( .A(\mem<0><12> ), .B(n1681), .Y(n2326) );
  OAI21X1 U1164 ( .A(n1783), .B(n1680), .C(n2325), .Y(n1812) );
  NAND2X1 U1165 ( .A(\mem<0><13> ), .B(n1681), .Y(n2325) );
  OAI21X1 U1167 ( .A(n1782), .B(n1680), .C(n2324), .Y(n1811) );
  NAND2X1 U1168 ( .A(\mem<0><14> ), .B(n1681), .Y(n2324) );
  OAI21X1 U1170 ( .A(n1780), .B(n1680), .C(n2323), .Y(n1810) );
  NAND2X1 U1171 ( .A(\mem<0><15> ), .B(n1681), .Y(n2323) );
  NOR3X1 U1174 ( .A(net60094), .B(net59638), .C(net60826), .Y(n2711) );
  NAND3X1 U1175 ( .A(net59460), .B(net59340), .C(n2709), .Y(n2322) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2709) );
  OR2X2 U3 ( .A(n2), .B(n1668), .Y(n40) );
  INVX1 U4 ( .A(net60826), .Y(\C2334/net60496 ) );
  INVX1 U5 ( .A(\C2334/net60504 ), .Y(\C2334/net60466 ) );
  INVX1 U6 ( .A(\C2334/net60506 ), .Y(\C2334/net60464 ) );
  INVX1 U7 ( .A(\C2334/net60506 ), .Y(\C2334/net60476 ) );
  INVX1 U8 ( .A(\C2334/net60506 ), .Y(\C2334/net60484 ) );
  INVX1 U9 ( .A(\C2334/net60504 ), .Y(\C2334/net60474 ) );
  INVX1 U10 ( .A(\C2334/net60506 ), .Y(\C2334/net60478 ) );
  INVX1 U11 ( .A(net100612), .Y(n1) );
  OR2X2 U12 ( .A(write), .B(rst), .Y(n2) );
  INVX1 U13 ( .A(net100612), .Y(net104441) );
  INVX1 U14 ( .A(n1666), .Y(n36) );
  INVX1 U15 ( .A(n1677), .Y(N19) );
  INVX1 U16 ( .A(net60828), .Y(\C2334/net60892 ) );
  INVX1 U17 ( .A(\C2334/net60160 ), .Y(\C2334/net59930 ) );
  INVX2 U18 ( .A(\C2334/net60504 ), .Y(\C2334/net60470 ) );
  INVX1 U19 ( .A(\C2334/net60892 ), .Y(\C2334/net60504 ) );
  INVX1 U20 ( .A(\C2334/net60892 ), .Y(\C2334/net60506 ) );
  INVX1 U21 ( .A(\C2334/net59930 ), .Y(\C2334/net59928 ) );
  INVX1 U22 ( .A(\C2334/net59930 ), .Y(\C2334/net59926 ) );
  INVX1 U23 ( .A(\C2334/net59930 ), .Y(\C2334/net59924 ) );
  INVX2 U24 ( .A(\C2334/net60496 ), .Y(n34) );
  INVX1 U25 ( .A(\C2334/net59930 ), .Y(\C2334/net59922 ) );
  INVX1 U26 ( .A(\C2334/net59930 ), .Y(\C2334/net59920 ) );
  INVX2 U27 ( .A(\C2334/net60496 ), .Y(\C2334/net60472 ) );
  INVX1 U28 ( .A(\C2334/net59930 ), .Y(\C2334/net59918 ) );
  INVX2 U29 ( .A(\C2334/net60504 ), .Y(\C2334/net60468 ) );
  INVX1 U30 ( .A(\C2334/net59934 ), .Y(\C2334/net59916 ) );
  INVX1 U31 ( .A(\C2334/net59934 ), .Y(\C2334/net59914 ) );
  INVX2 U32 ( .A(\C2334/net60506 ), .Y(\C2334/net60462 ) );
  INVX2 U33 ( .A(\C2334/net60506 ), .Y(\C2334/net60460 ) );
  INVX1 U34 ( .A(\C2334/net59934 ), .Y(\C2334/net59912 ) );
  INVX1 U35 ( .A(\C2334/net59934 ), .Y(\C2334/net59910 ) );
  INVX1 U36 ( .A(\C2334/net60506 ), .Y(\C2334/net60452 ) );
  INVX2 U37 ( .A(\C2334/net59934 ), .Y(\C2334/net59908 ) );
  INVX1 U38 ( .A(n1667), .Y(N31) );
  INVX1 U39 ( .A(net104441), .Y(n3) );
  OR2X2 U40 ( .A(n3), .B(\C2334/net11880 ), .Y(net100597) );
  OR2X2 U41 ( .A(write), .B(rst), .Y(net100612) );
  INVX1 U42 ( .A(n1), .Y(net101600) );
  OR2X2 U43 ( .A(n2), .B(\C2334/net11884 ), .Y(net100591) );
  INVX1 U44 ( .A(net100597), .Y(net100598) );
  MUX2X1 U45 ( .B(n31), .A(n16), .S(\C2334/net59380 ), .Y(\C2334/net11880 ) );
  MUX2X1 U46 ( .B(n32), .A(n33), .S(\C2334/net59512 ), .Y(n31) );
  MUX2X1 U47 ( .B(n28), .A(n25), .S(\C2334/net59712 ), .Y(n32) );
  MUX2X1 U48 ( .B(n29), .A(n30), .S(\C2334/net59922 ), .Y(n28) );
  MUX2X1 U49 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(\C2334/net60472 ), .Y(n29)
         );
  MUX2X1 U50 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(\C2334/net60460 ), .Y(n30)
         );
  MUX2X1 U51 ( .B(n26), .A(n27), .S(\C2334/net59922 ), .Y(n25) );
  MUX2X1 U52 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(\C2334/net60468 ), .Y(n26)
         );
  MUX2X1 U53 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(\C2334/net60470 ), .Y(n27)
         );
  INVX1 U54 ( .A(net59640), .Y(\C2334/net59712 ) );
  MUX2X1 U55 ( .B(n22), .A(n19), .S(\C2334/net59712 ), .Y(n33) );
  MUX2X1 U56 ( .B(n23), .A(n24), .S(\C2334/net59922 ), .Y(n22) );
  MUX2X1 U57 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n34), .Y(n23) );
  MUX2X1 U58 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n34), .Y(n24) );
  MUX2X1 U59 ( .B(n20), .A(n21), .S(\C2334/net59922 ), .Y(n19) );
  MUX2X1 U60 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n34), .Y(n20) );
  MUX2X1 U93 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n34), .Y(n21) );
  INVX1 U94 ( .A(net59460), .Y(\C2334/net59512 ) );
  MUX2X1 U127 ( .B(n17), .A(n18), .S(\C2334/net59512 ), .Y(n16) );
  MUX2X1 U128 ( .B(n13), .A(n10), .S(\C2334/net59712 ), .Y(n17) );
  MUX2X1 U161 ( .B(n14), .A(n15), .S(\C2334/net59922 ), .Y(n13) );
  MUX2X1 U162 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n34), .Y(n14) );
  MUX2X1 U195 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n34), .Y(n15) );
  MUX2X1 U196 ( .B(n11), .A(n12), .S(\C2334/net59922 ), .Y(n10) );
  MUX2X1 U229 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n34), .Y(n11) );
  MUX2X1 U230 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n34), .Y(n12) );
  MUX2X1 U263 ( .B(n7), .A(n4), .S(\C2334/net59712 ), .Y(n18) );
  MUX2X1 U264 ( .B(n8), .A(n9), .S(\C2334/net59922 ), .Y(n7) );
  MUX2X1 U297 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n34), .Y(n8) );
  MUX2X1 U298 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n34), .Y(n9) );
  MUX2X1 U331 ( .B(n5), .A(n6), .S(\C2334/net59922 ), .Y(n4) );
  MUX2X1 U332 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n34), .Y(n5) );
  MUX2X1 U366 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n34), .Y(n6) );
  INVX1 U367 ( .A(net59340), .Y(\C2334/net59380 ) );
  AND2X2 U400 ( .A(net101601), .B(n36), .Y(\data_out<0> ) );
  INVX1 U401 ( .A(net59640), .Y(\C2334/net59710 ) );
  INVX1 U434 ( .A(N13), .Y(net59460) );
  INVX1 U435 ( .A(net59460), .Y(\C2334/net59514 ) );
  INVX1 U468 ( .A(net60096), .Y(net60094) );
  INVX1 U469 ( .A(net60096), .Y(\C2334/net60160 ) );
  INVX1 U502 ( .A(net60828), .Y(net60826) );
  INVX1 U503 ( .A(N14), .Y(net59340) );
  INVX1 U536 ( .A(rst), .Y(net59006) );
  INVX1 U537 ( .A(net59640), .Y(net59638) );
  INVX2 U570 ( .A(N12), .Y(net59640) );
  INVX2 U571 ( .A(\C2334/net60496 ), .Y(\C2334/net60490 ) );
  INVX1 U604 ( .A(net59638), .Y(\C2334/net59722 ) );
  INVX1 U605 ( .A(\C2334/net59722 ), .Y(\C2334/net59716 ) );
  INVX1 U639 ( .A(\C2334/net59722 ), .Y(\C2334/net59718 ) );
  INVX1 U640 ( .A(\C2334/net60160 ), .Y(\C2334/net59934 ) );
  INVX1 U673 ( .A(n1203), .Y(n1737) );
  INVX1 U674 ( .A(n1204), .Y(n1740) );
  INVX1 U707 ( .A(n1205), .Y(n1743) );
  INVX1 U708 ( .A(n1206), .Y(n1746) );
  INVX1 U741 ( .A(n1207), .Y(n1749) );
  INVX1 U742 ( .A(n1208), .Y(n1752) );
  INVX1 U775 ( .A(n1209), .Y(n1755) );
  INVX1 U776 ( .A(n1210), .Y(n1758) );
  INVX1 U809 ( .A(n1211), .Y(n1761) );
  INVX1 U810 ( .A(n1212), .Y(n1764) );
  INVX1 U843 ( .A(n1213), .Y(n1767) );
  INVX1 U844 ( .A(n1214), .Y(n1770) );
  INVX1 U877 ( .A(n1215), .Y(n1773) );
  INVX1 U878 ( .A(n1184), .Y(n1680) );
  INVX1 U912 ( .A(n1185), .Y(n1683) );
  INVX1 U913 ( .A(n1186), .Y(n1686) );
  INVX1 U947 ( .A(n1187), .Y(n1689) );
  INVX1 U948 ( .A(n1188), .Y(n1692) );
  INVX1 U982 ( .A(n1189), .Y(n1695) );
  INVX1 U983 ( .A(n1190), .Y(n1698) );
  INVX1 U1017 ( .A(n1191), .Y(n1701) );
  INVX1 U1018 ( .A(n1192), .Y(n1704) );
  INVX1 U1052 ( .A(n1193), .Y(n1707) );
  INVX1 U1053 ( .A(n1194), .Y(n1710) );
  INVX1 U1087 ( .A(n1195), .Y(n1713) );
  INVX1 U1088 ( .A(n1196), .Y(n1716) );
  INVX1 U1122 ( .A(n1197), .Y(n1719) );
  INVX1 U1123 ( .A(n1198), .Y(n1722) );
  INVX1 U1127 ( .A(n1199), .Y(n1725) );
  INVX1 U1130 ( .A(n1200), .Y(n1728) );
  INVX1 U1133 ( .A(n1201), .Y(n1731) );
  INVX1 U1136 ( .A(n1202), .Y(n1734) );
  INVX4 U1139 ( .A(n2831), .Y(n1779) );
  OR2X2 U1142 ( .A(write), .B(rst), .Y(n37) );
  INVX1 U1145 ( .A(net104441), .Y(net104291) );
  AND2X2 U1148 ( .A(n1), .B(N31), .Y(\data_out<1> ) );
  INVX1 U1151 ( .A(net104291), .Y(net101601) );
  OR2X2 U1154 ( .A(n2), .B(n1674), .Y(n56) );
  AND2X2 U1157 ( .A(net101601), .B(N19), .Y(\data_out<13> ) );
  OR2X2 U1160 ( .A(net101600), .B(n1672), .Y(n48) );
  OR2X2 U1163 ( .A(n37), .B(n1671), .Y(n45) );
  OR2X2 U1166 ( .A(n37), .B(n1670), .Y(n43) );
  OR2X2 U1169 ( .A(n37), .B(n1669), .Y(n41) );
  OR2X2 U1172 ( .A(n2), .B(n1679), .Y(n64) );
  OR2X2 U1173 ( .A(n37), .B(n1676), .Y(n60) );
  OR2X2 U1177 ( .A(n37), .B(n1678), .Y(n62) );
  OR2X2 U1178 ( .A(n2), .B(n1675), .Y(n58) );
  OR2X2 U1179 ( .A(n2), .B(n1673), .Y(n52) );
  INVX1 U1180 ( .A(n41), .Y(\data_out<3> ) );
  INVX1 U1181 ( .A(n43), .Y(\data_out<5> ) );
  INVX1 U1182 ( .A(n45), .Y(\data_out<7> ) );
  INVX1 U1183 ( .A(n48), .Y(\data_out<8> ) );
  INVX1 U1184 ( .A(n52), .Y(\data_out<9> ) );
  AND2X2 U1185 ( .A(n1184), .B(n1778), .Y(n66) );
  INVX1 U1186 ( .A(n66), .Y(n68) );
  AND2X2 U1187 ( .A(\data_in<7> ), .B(n1777), .Y(n70) );
  AND2X2 U1188 ( .A(\data_in<6> ), .B(n1777), .Y(n72) );
  AND2X2 U1189 ( .A(\data_in<5> ), .B(n1777), .Y(n74) );
  AND2X2 U1190 ( .A(\data_in<4> ), .B(n1777), .Y(n76) );
  AND2X2 U1191 ( .A(\data_in<3> ), .B(n1777), .Y(n80) );
  AND2X2 U1192 ( .A(\data_in<2> ), .B(n1777), .Y(n82) );
  AND2X2 U1193 ( .A(\data_in<1> ), .B(n1777), .Y(n99) );
  AND2X2 U1194 ( .A(\data_in<0> ), .B(n1777), .Y(n101) );
  AND2X2 U1195 ( .A(n1185), .B(n1777), .Y(n118) );
  INVX1 U1196 ( .A(n118), .Y(n120) );
  AND2X2 U1197 ( .A(n1186), .B(n1777), .Y(n137) );
  INVX1 U1198 ( .A(n137), .Y(n139) );
  AND2X2 U1199 ( .A(n1187), .B(n1777), .Y(n156) );
  INVX1 U1200 ( .A(n156), .Y(n158) );
  AND2X2 U1201 ( .A(n1188), .B(n1777), .Y(n175) );
  INVX1 U1202 ( .A(n175), .Y(n177) );
  AND2X2 U1203 ( .A(n1189), .B(n1777), .Y(n194) );
  INVX1 U1204 ( .A(n194), .Y(n196) );
  AND2X2 U1205 ( .A(n1190), .B(n1776), .Y(n215) );
  INVX1 U1206 ( .A(n215), .Y(n217) );
  AND2X2 U1207 ( .A(n1191), .B(n1776), .Y(n233) );
  INVX1 U1208 ( .A(n233), .Y(n235) );
  AND2X2 U1209 ( .A(n1192), .B(n1776), .Y(n251) );
  INVX1 U1210 ( .A(n251), .Y(n253) );
  AND2X2 U1211 ( .A(n1193), .B(n1776), .Y(n269) );
  INVX1 U1212 ( .A(n269), .Y(n271) );
  AND2X2 U1213 ( .A(n1194), .B(n1776), .Y(n287) );
  INVX1 U1214 ( .A(n287), .Y(n289) );
  AND2X2 U1215 ( .A(n1195), .B(n1776), .Y(n305) );
  INVX1 U1216 ( .A(n305), .Y(n307) );
  AND2X2 U1217 ( .A(n1196), .B(n1776), .Y(n323) );
  INVX1 U1218 ( .A(n323), .Y(n325) );
  AND2X2 U1219 ( .A(n1197), .B(n1776), .Y(n341) );
  INVX1 U1220 ( .A(n341), .Y(n343) );
  AND2X2 U1221 ( .A(n1198), .B(n1776), .Y(n360) );
  INVX1 U1222 ( .A(n360), .Y(n362) );
  AND2X2 U1223 ( .A(n1199), .B(n1776), .Y(n378) );
  INVX1 U1224 ( .A(n378), .Y(n380) );
  AND2X2 U1225 ( .A(n1200), .B(n1776), .Y(n396) );
  INVX1 U1226 ( .A(n396), .Y(n398) );
  AND2X2 U1227 ( .A(n1201), .B(n1776), .Y(n414) );
  INVX1 U1228 ( .A(n414), .Y(n416) );
  AND2X2 U1229 ( .A(n1202), .B(n1776), .Y(n432) );
  INVX1 U1230 ( .A(n432), .Y(n434) );
  AND2X2 U1231 ( .A(n1203), .B(n1778), .Y(n450) );
  INVX1 U1232 ( .A(n450), .Y(n452) );
  AND2X2 U1233 ( .A(n1204), .B(n1778), .Y(n468) );
  INVX1 U1234 ( .A(n468), .Y(n470) );
  AND2X2 U1235 ( .A(n1205), .B(n1778), .Y(n486) );
  INVX1 U1236 ( .A(n486), .Y(n488) );
  AND2X2 U1237 ( .A(n1206), .B(n1777), .Y(n505) );
  INVX1 U1238 ( .A(n505), .Y(n507) );
  AND2X2 U1239 ( .A(n1207), .B(n1776), .Y(n523) );
  INVX1 U1240 ( .A(n523), .Y(n525) );
  AND2X2 U1241 ( .A(n1208), .B(n1778), .Y(n541) );
  INVX1 U1242 ( .A(n541), .Y(n543) );
  AND2X2 U1243 ( .A(n1209), .B(n1777), .Y(n559) );
  INVX1 U1244 ( .A(n559), .Y(n561) );
  AND2X2 U1245 ( .A(n1210), .B(n1776), .Y(n577) );
  INVX1 U1246 ( .A(n577), .Y(n579) );
  AND2X2 U1247 ( .A(n1211), .B(n1778), .Y(n595) );
  INVX1 U1248 ( .A(n595), .Y(n597) );
  AND2X2 U1249 ( .A(n1212), .B(n1777), .Y(n613) );
  INVX1 U1250 ( .A(n613), .Y(n615) );
  AND2X2 U1251 ( .A(n1213), .B(n1776), .Y(n631) );
  INVX1 U1252 ( .A(n631), .Y(n633) );
  AND2X2 U1253 ( .A(n1214), .B(n1778), .Y(n650) );
  INVX1 U1254 ( .A(n650), .Y(n1163) );
  AND2X2 U1255 ( .A(n1215), .B(n1778), .Y(n1164) );
  INVX1 U1256 ( .A(n1164), .Y(n1165) );
  BUFX2 U1257 ( .A(n68), .Y(n1681) );
  BUFX2 U1258 ( .A(n68), .Y(n1682) );
  BUFX2 U1259 ( .A(n120), .Y(n1684) );
  BUFX2 U1260 ( .A(n120), .Y(n1685) );
  BUFX2 U1261 ( .A(n139), .Y(n1687) );
  BUFX2 U1262 ( .A(n139), .Y(n1688) );
  BUFX2 U1263 ( .A(n158), .Y(n1690) );
  BUFX2 U1264 ( .A(n158), .Y(n1691) );
  BUFX2 U1265 ( .A(n177), .Y(n1693) );
  BUFX2 U1266 ( .A(n177), .Y(n1694) );
  BUFX2 U1267 ( .A(n196), .Y(n1696) );
  BUFX2 U1268 ( .A(n196), .Y(n1697) );
  BUFX2 U1269 ( .A(n217), .Y(n1699) );
  BUFX2 U1270 ( .A(n217), .Y(n1700) );
  BUFX2 U1271 ( .A(n235), .Y(n1702) );
  BUFX2 U1272 ( .A(n235), .Y(n1703) );
  BUFX2 U1273 ( .A(n253), .Y(n1705) );
  BUFX2 U1274 ( .A(n253), .Y(n1706) );
  BUFX2 U1275 ( .A(n271), .Y(n1708) );
  BUFX2 U1276 ( .A(n271), .Y(n1709) );
  BUFX2 U1277 ( .A(n289), .Y(n1711) );
  BUFX2 U1278 ( .A(n289), .Y(n1712) );
  BUFX2 U1279 ( .A(n307), .Y(n1714) );
  BUFX2 U1280 ( .A(n307), .Y(n1715) );
  BUFX2 U1281 ( .A(n325), .Y(n1717) );
  BUFX2 U1282 ( .A(n325), .Y(n1718) );
  BUFX2 U1283 ( .A(n343), .Y(n1720) );
  BUFX2 U1284 ( .A(n343), .Y(n1721) );
  BUFX2 U1285 ( .A(n362), .Y(n1723) );
  BUFX2 U1286 ( .A(n362), .Y(n1724) );
  BUFX2 U1287 ( .A(n380), .Y(n1726) );
  BUFX2 U1288 ( .A(n380), .Y(n1727) );
  BUFX2 U1289 ( .A(n398), .Y(n1729) );
  BUFX2 U1290 ( .A(n398), .Y(n1730) );
  BUFX2 U1291 ( .A(n416), .Y(n1732) );
  BUFX2 U1292 ( .A(n416), .Y(n1733) );
  BUFX2 U1293 ( .A(n434), .Y(n1735) );
  BUFX2 U1294 ( .A(n434), .Y(n1736) );
  BUFX2 U1295 ( .A(n452), .Y(n1738) );
  BUFX2 U1296 ( .A(n452), .Y(n1739) );
  BUFX2 U1297 ( .A(n470), .Y(n1741) );
  BUFX2 U1298 ( .A(n470), .Y(n1742) );
  BUFX2 U1299 ( .A(n488), .Y(n1744) );
  BUFX2 U1300 ( .A(n488), .Y(n1745) );
  BUFX2 U1301 ( .A(n507), .Y(n1747) );
  BUFX2 U1302 ( .A(n507), .Y(n1748) );
  BUFX2 U1303 ( .A(n525), .Y(n1750) );
  BUFX2 U1304 ( .A(n525), .Y(n1751) );
  BUFX2 U1305 ( .A(n543), .Y(n1753) );
  BUFX2 U1306 ( .A(n543), .Y(n1754) );
  BUFX2 U1307 ( .A(n561), .Y(n1756) );
  BUFX2 U1308 ( .A(n561), .Y(n1757) );
  BUFX2 U1309 ( .A(n579), .Y(n1759) );
  BUFX2 U1310 ( .A(n579), .Y(n1760) );
  BUFX2 U1311 ( .A(n597), .Y(n1762) );
  BUFX2 U1312 ( .A(n597), .Y(n1763) );
  BUFX2 U1313 ( .A(n615), .Y(n1765) );
  BUFX2 U1314 ( .A(n615), .Y(n1766) );
  BUFX2 U1315 ( .A(n633), .Y(n1768) );
  BUFX2 U1316 ( .A(n633), .Y(n1769) );
  BUFX2 U1317 ( .A(n1163), .Y(n1771) );
  BUFX2 U1318 ( .A(n1163), .Y(n1772) );
  BUFX2 U1319 ( .A(n1165), .Y(n1774) );
  BUFX2 U1320 ( .A(n1165), .Y(n1775) );
  INVX1 U1321 ( .A(net59460), .Y(net59458) );
  AND2X2 U1322 ( .A(\data_in<15> ), .B(n1778), .Y(n1166) );
  AND2X2 U1323 ( .A(\data_in<14> ), .B(n1778), .Y(n1167) );
  AND2X2 U1324 ( .A(\data_in<13> ), .B(n1778), .Y(n1168) );
  AND2X2 U1325 ( .A(\data_in<12> ), .B(n1778), .Y(n1169) );
  AND2X2 U1326 ( .A(\data_in<11> ), .B(n1778), .Y(n1170) );
  AND2X2 U1327 ( .A(\data_in<10> ), .B(n1778), .Y(n1171) );
  AND2X2 U1328 ( .A(\data_in<9> ), .B(n1778), .Y(n1172) );
  AND2X2 U1329 ( .A(\data_in<8> ), .B(n1778), .Y(n1173) );
  BUFX2 U1330 ( .A(n2322), .Y(n1174) );
  INVX1 U1331 ( .A(n1174), .Y(n1806) );
  BUFX2 U1332 ( .A(n2451), .Y(n1175) );
  INVX1 U1333 ( .A(n1175), .Y(n1809) );
  BUFX2 U1334 ( .A(n2580), .Y(n1176) );
  INVX1 U1335 ( .A(n1176), .Y(n1807) );
  BUFX2 U1336 ( .A(n2710), .Y(n1177) );
  INVX1 U1337 ( .A(n1177), .Y(n1808) );
  INVX1 U1338 ( .A(n40), .Y(\data_out<2> ) );
  INVX1 U1339 ( .A(net100591), .Y(net80056) );
  INVX1 U1340 ( .A(n56), .Y(\data_out<10> ) );
  INVX1 U1341 ( .A(n58), .Y(\data_out<11> ) );
  INVX1 U1342 ( .A(n60), .Y(\data_out<12> ) );
  INVX1 U1343 ( .A(n62), .Y(\data_out<14> ) );
  INVX1 U1344 ( .A(n64), .Y(\data_out<15> ) );
  AND2X1 U1345 ( .A(n1806), .B(n2711), .Y(n1184) );
  AND2X1 U1346 ( .A(n1806), .B(n2728), .Y(n1185) );
  AND2X1 U1347 ( .A(n1806), .B(n2745), .Y(n1186) );
  AND2X1 U1348 ( .A(n1806), .B(n2762), .Y(n1187) );
  AND2X1 U1349 ( .A(n1806), .B(n2779), .Y(n1188) );
  AND2X1 U1350 ( .A(n1806), .B(n2796), .Y(n1189) );
  AND2X1 U1351 ( .A(n1806), .B(n2813), .Y(n1190) );
  AND2X1 U1352 ( .A(n1806), .B(n2830), .Y(n1191) );
  AND2X1 U1353 ( .A(n1809), .B(n2711), .Y(n1192) );
  AND2X1 U1354 ( .A(n1809), .B(n2728), .Y(n1193) );
  AND2X1 U1355 ( .A(n1809), .B(n2745), .Y(n1194) );
  AND2X1 U1356 ( .A(n1809), .B(n2762), .Y(n1195) );
  AND2X1 U1357 ( .A(n1809), .B(n2779), .Y(n1196) );
  AND2X1 U1358 ( .A(n1809), .B(n2796), .Y(n1197) );
  AND2X1 U1359 ( .A(n1809), .B(n2813), .Y(n1198) );
  AND2X1 U1360 ( .A(n1809), .B(n2830), .Y(n1199) );
  AND2X1 U1361 ( .A(n1807), .B(n2711), .Y(n1200) );
  AND2X1 U1362 ( .A(n1807), .B(n2728), .Y(n1201) );
  AND2X1 U1363 ( .A(n1807), .B(n2745), .Y(n1202) );
  AND2X1 U1364 ( .A(n1807), .B(n2762), .Y(n1203) );
  AND2X1 U1365 ( .A(n1807), .B(n2779), .Y(n1204) );
  AND2X1 U1366 ( .A(n1807), .B(n2796), .Y(n1205) );
  AND2X1 U1367 ( .A(n1807), .B(n2813), .Y(n1206) );
  AND2X1 U1368 ( .A(n1807), .B(n2830), .Y(n1207) );
  AND2X1 U1369 ( .A(n2711), .B(n1808), .Y(n1208) );
  AND2X1 U1370 ( .A(n2728), .B(n1808), .Y(n1209) );
  AND2X1 U1371 ( .A(n2745), .B(n1808), .Y(n1210) );
  AND2X1 U1372 ( .A(n2762), .B(n1808), .Y(n1211) );
  AND2X1 U1373 ( .A(n2779), .B(n1808), .Y(n1212) );
  AND2X1 U1374 ( .A(n2796), .B(n1808), .Y(n1213) );
  AND2X1 U1375 ( .A(n2813), .B(n1808), .Y(n1214) );
  AND2X1 U1376 ( .A(n2830), .B(n1808), .Y(n1215) );
  MUX2X1 U1377 ( .B(n1217), .A(n1218), .S(\C2334/net59928 ), .Y(n1216) );
  MUX2X1 U1378 ( .B(n1220), .A(n1221), .S(\C2334/net59928 ), .Y(n1219) );
  MUX2X1 U1379 ( .B(n1223), .A(n1224), .S(\C2334/net59928 ), .Y(n1222) );
  MUX2X1 U1380 ( .B(n1226), .A(n1227), .S(\C2334/net59928 ), .Y(n1225) );
  MUX2X1 U1381 ( .B(n1229), .A(n1230), .S(\C2334/net59512 ), .Y(n1228) );
  MUX2X1 U1382 ( .B(n1232), .A(n1233), .S(\C2334/net59928 ), .Y(n1231) );
  MUX2X1 U1383 ( .B(n1235), .A(n1236), .S(\C2334/net59928 ), .Y(n1234) );
  MUX2X1 U1384 ( .B(n1238), .A(n1239), .S(\C2334/net59928 ), .Y(n1237) );
  MUX2X1 U1385 ( .B(n1241), .A(n1242), .S(\C2334/net59928 ), .Y(n1240) );
  MUX2X1 U1386 ( .B(n1244), .A(n1245), .S(\C2334/net59512 ), .Y(n1243) );
  MUX2X1 U1387 ( .B(n1247), .A(n1248), .S(\C2334/net59926 ), .Y(n1246) );
  MUX2X1 U1388 ( .B(n1250), .A(n1251), .S(\C2334/net59926 ), .Y(n1249) );
  MUX2X1 U1389 ( .B(n1253), .A(n1254), .S(\C2334/net59926 ), .Y(n1252) );
  MUX2X1 U1390 ( .B(n1256), .A(n1257), .S(\C2334/net59926 ), .Y(n1255) );
  MUX2X1 U1391 ( .B(n1259), .A(n1260), .S(\C2334/net59512 ), .Y(n1258) );
  MUX2X1 U1392 ( .B(n1262), .A(n1263), .S(\C2334/net59926 ), .Y(n1261) );
  MUX2X1 U1393 ( .B(n1265), .A(n1266), .S(\C2334/net59926 ), .Y(n1264) );
  MUX2X1 U1394 ( .B(n1268), .A(n1269), .S(\C2334/net59926 ), .Y(n1267) );
  MUX2X1 U1395 ( .B(n1271), .A(n1272), .S(\C2334/net59926 ), .Y(n1270) );
  MUX2X1 U1396 ( .B(n1274), .A(n1275), .S(\C2334/net59512 ), .Y(n1273) );
  MUX2X1 U1397 ( .B(n1277), .A(n1278), .S(\C2334/net59926 ), .Y(n1276) );
  MUX2X1 U1398 ( .B(n1280), .A(n1281), .S(\C2334/net59926 ), .Y(n1279) );
  MUX2X1 U1399 ( .B(n1283), .A(n1284), .S(\C2334/net59926 ), .Y(n1282) );
  MUX2X1 U1400 ( .B(n1286), .A(n1287), .S(\C2334/net59926 ), .Y(n1285) );
  MUX2X1 U1401 ( .B(n1289), .A(n1290), .S(\C2334/net59512 ), .Y(n1288) );
  MUX2X1 U1402 ( .B(n1292), .A(n1293), .S(\C2334/net59924 ), .Y(n1291) );
  MUX2X1 U1403 ( .B(n1295), .A(n1296), .S(\C2334/net59924 ), .Y(n1294) );
  MUX2X1 U1404 ( .B(n1298), .A(n1299), .S(\C2334/net59924 ), .Y(n1297) );
  MUX2X1 U1405 ( .B(n1301), .A(n1302), .S(\C2334/net59924 ), .Y(n1300) );
  MUX2X1 U1406 ( .B(n1304), .A(n1305), .S(\C2334/net59512 ), .Y(n1303) );
  MUX2X1 U1407 ( .B(n1307), .A(n1308), .S(\C2334/net59924 ), .Y(n1306) );
  MUX2X1 U1408 ( .B(n1310), .A(n1311), .S(\C2334/net59924 ), .Y(n1309) );
  MUX2X1 U1409 ( .B(n1313), .A(n1314), .S(\C2334/net59924 ), .Y(n1312) );
  MUX2X1 U1410 ( .B(n1316), .A(n1317), .S(\C2334/net59924 ), .Y(n1315) );
  MUX2X1 U1411 ( .B(n1319), .A(n1320), .S(\C2334/net59512 ), .Y(n1318) );
  MUX2X1 U1412 ( .B(n1322), .A(n1323), .S(\C2334/net59924 ), .Y(n1321) );
  MUX2X1 U1413 ( .B(n1325), .A(n1326), .S(\C2334/net59924 ), .Y(n1324) );
  MUX2X1 U1414 ( .B(n1328), .A(n1329), .S(\C2334/net59924 ), .Y(n1327) );
  MUX2X1 U1415 ( .B(n1331), .A(n1332), .S(\C2334/net59924 ), .Y(n1330) );
  MUX2X1 U1416 ( .B(n1334), .A(n1335), .S(\C2334/net59512 ), .Y(n1333) );
  MUX2X1 U1417 ( .B(n1337), .A(n1338), .S(\C2334/net59922 ), .Y(n1336) );
  MUX2X1 U1418 ( .B(n1340), .A(n1341), .S(\C2334/net59922 ), .Y(n1339) );
  MUX2X1 U1419 ( .B(n1343), .A(n1344), .S(\C2334/net59922 ), .Y(n1342) );
  MUX2X1 U1420 ( .B(n1346), .A(n1347), .S(\C2334/net59922 ), .Y(n1345) );
  MUX2X1 U1421 ( .B(n1349), .A(n1350), .S(\C2334/net59512 ), .Y(n1348) );
  MUX2X1 U1422 ( .B(n1352), .A(n1353), .S(\C2334/net59920 ), .Y(n1351) );
  MUX2X1 U1423 ( .B(n1355), .A(n1356), .S(\C2334/net59920 ), .Y(n1354) );
  MUX2X1 U1424 ( .B(n1358), .A(n1359), .S(\C2334/net59920 ), .Y(n1357) );
  MUX2X1 U1425 ( .B(n1361), .A(n1362), .S(\C2334/net59920 ), .Y(n1360) );
  MUX2X1 U1426 ( .B(n1364), .A(n1365), .S(\C2334/net59512 ), .Y(n1363) );
  MUX2X1 U1427 ( .B(n1367), .A(n1368), .S(\C2334/net59920 ), .Y(n1366) );
  MUX2X1 U1428 ( .B(n1370), .A(n1371), .S(\C2334/net59920 ), .Y(n1369) );
  MUX2X1 U1429 ( .B(n1373), .A(n1374), .S(\C2334/net59920 ), .Y(n1372) );
  MUX2X1 U1430 ( .B(n1376), .A(n1377), .S(\C2334/net59920 ), .Y(n1375) );
  MUX2X1 U1431 ( .B(n1379), .A(n1380), .S(\C2334/net59514 ), .Y(n1378) );
  MUX2X1 U1432 ( .B(n1382), .A(n1383), .S(\C2334/net59920 ), .Y(n1381) );
  MUX2X1 U1433 ( .B(n1385), .A(n1386), .S(\C2334/net59920 ), .Y(n1384) );
  MUX2X1 U1434 ( .B(n1388), .A(n1389), .S(\C2334/net59920 ), .Y(n1387) );
  MUX2X1 U1435 ( .B(n1391), .A(n1392), .S(\C2334/net59920 ), .Y(n1390) );
  MUX2X1 U1436 ( .B(n1394), .A(n1395), .S(\C2334/net59514 ), .Y(n1393) );
  MUX2X1 U1437 ( .B(n1397), .A(n1398), .S(\C2334/net59918 ), .Y(n1396) );
  MUX2X1 U1438 ( .B(n1400), .A(n1401), .S(\C2334/net59918 ), .Y(n1399) );
  MUX2X1 U1439 ( .B(n1403), .A(n1404), .S(\C2334/net59918 ), .Y(n1402) );
  MUX2X1 U1440 ( .B(n1406), .A(n1407), .S(\C2334/net59918 ), .Y(n1405) );
  MUX2X1 U1441 ( .B(n1409), .A(n1410), .S(\C2334/net59514 ), .Y(n1408) );
  MUX2X1 U1442 ( .B(n1412), .A(n1413), .S(\C2334/net59918 ), .Y(n1411) );
  MUX2X1 U1443 ( .B(n1415), .A(n1416), .S(\C2334/net59918 ), .Y(n1414) );
  MUX2X1 U1444 ( .B(n1418), .A(n1419), .S(\C2334/net59918 ), .Y(n1417) );
  MUX2X1 U1445 ( .B(n1421), .A(n1422), .S(\C2334/net59918 ), .Y(n1420) );
  MUX2X1 U1446 ( .B(n1424), .A(n1425), .S(\C2334/net59514 ), .Y(n1423) );
  MUX2X1 U1447 ( .B(n1427), .A(n1428), .S(\C2334/net59918 ), .Y(n1426) );
  MUX2X1 U1448 ( .B(n1430), .A(n1431), .S(\C2334/net59918 ), .Y(n1429) );
  MUX2X1 U1449 ( .B(n1433), .A(n1434), .S(\C2334/net59918 ), .Y(n1432) );
  MUX2X1 U1450 ( .B(n1436), .A(n1437), .S(\C2334/net59918 ), .Y(n1435) );
  MUX2X1 U1451 ( .B(n1439), .A(n1440), .S(\C2334/net59514 ), .Y(n1438) );
  MUX2X1 U1452 ( .B(n1442), .A(n1443), .S(\C2334/net59916 ), .Y(n1441) );
  MUX2X1 U1453 ( .B(n1445), .A(n1446), .S(\C2334/net59916 ), .Y(n1444) );
  MUX2X1 U1454 ( .B(n1448), .A(n1449), .S(\C2334/net59916 ), .Y(n1447) );
  MUX2X1 U1455 ( .B(n1451), .A(n1452), .S(\C2334/net59916 ), .Y(n1450) );
  MUX2X1 U1456 ( .B(n1454), .A(n1455), .S(\C2334/net59514 ), .Y(n1453) );
  MUX2X1 U1457 ( .B(n1457), .A(n1458), .S(\C2334/net59916 ), .Y(n1456) );
  MUX2X1 U1458 ( .B(n1460), .A(n1461), .S(\C2334/net59916 ), .Y(n1459) );
  MUX2X1 U1459 ( .B(n1463), .A(n1464), .S(\C2334/net59916 ), .Y(n1462) );
  MUX2X1 U1460 ( .B(n1466), .A(n1467), .S(\C2334/net59916 ), .Y(n1465) );
  MUX2X1 U1461 ( .B(n1469), .A(n1470), .S(\C2334/net59514 ), .Y(n1468) );
  MUX2X1 U1462 ( .B(n1472), .A(n1473), .S(\C2334/net59916 ), .Y(n1471) );
  MUX2X1 U1463 ( .B(n1475), .A(n1476), .S(\C2334/net59916 ), .Y(n1474) );
  MUX2X1 U1464 ( .B(n1478), .A(n1479), .S(\C2334/net59916 ), .Y(n1477) );
  MUX2X1 U1465 ( .B(n1481), .A(n1482), .S(\C2334/net59916 ), .Y(n1480) );
  MUX2X1 U1466 ( .B(n1484), .A(n1485), .S(\C2334/net59514 ), .Y(n1483) );
  MUX2X1 U1467 ( .B(n1487), .A(n1488), .S(\C2334/net59914 ), .Y(n1486) );
  MUX2X1 U1468 ( .B(n1490), .A(n1491), .S(\C2334/net59914 ), .Y(n1489) );
  MUX2X1 U1469 ( .B(n1493), .A(n1494), .S(\C2334/net59914 ), .Y(n1492) );
  MUX2X1 U1470 ( .B(n1496), .A(n1497), .S(\C2334/net59914 ), .Y(n1495) );
  MUX2X1 U1471 ( .B(n1499), .A(n1500), .S(\C2334/net59514 ), .Y(n1498) );
  MUX2X1 U1472 ( .B(n1502), .A(n1503), .S(\C2334/net59914 ), .Y(n1501) );
  MUX2X1 U1473 ( .B(n1505), .A(n1506), .S(\C2334/net59914 ), .Y(n1504) );
  MUX2X1 U1474 ( .B(n1508), .A(n1509), .S(\C2334/net59914 ), .Y(n1507) );
  MUX2X1 U1475 ( .B(n1511), .A(n1512), .S(\C2334/net59914 ), .Y(n1510) );
  MUX2X1 U1476 ( .B(n1514), .A(n1515), .S(\C2334/net59514 ), .Y(n1513) );
  MUX2X1 U1477 ( .B(n1517), .A(n1518), .S(\C2334/net59914 ), .Y(n1516) );
  MUX2X1 U1478 ( .B(n1520), .A(n1521), .S(\C2334/net59914 ), .Y(n1519) );
  MUX2X1 U1479 ( .B(n1523), .A(n1524), .S(\C2334/net59914 ), .Y(n1522) );
  MUX2X1 U1480 ( .B(n1526), .A(n1527), .S(\C2334/net59914 ), .Y(n1525) );
  MUX2X1 U1481 ( .B(n1529), .A(n1530), .S(\C2334/net59514 ), .Y(n1528) );
  MUX2X1 U1482 ( .B(n1532), .A(n1533), .S(\C2334/net59912 ), .Y(n1531) );
  MUX2X1 U1483 ( .B(n1535), .A(n1536), .S(\C2334/net59912 ), .Y(n1534) );
  MUX2X1 U1484 ( .B(n1538), .A(n1539), .S(\C2334/net59912 ), .Y(n1537) );
  MUX2X1 U1485 ( .B(n1541), .A(n1542), .S(\C2334/net59912 ), .Y(n1540) );
  MUX2X1 U1486 ( .B(n1544), .A(n1545), .S(\C2334/net59514 ), .Y(n1543) );
  MUX2X1 U1487 ( .B(n1547), .A(n1548), .S(\C2334/net59912 ), .Y(n1546) );
  MUX2X1 U1488 ( .B(n1550), .A(n1551), .S(\C2334/net59912 ), .Y(n1549) );
  MUX2X1 U1489 ( .B(n1553), .A(n1554), .S(\C2334/net59912 ), .Y(n1552) );
  MUX2X1 U1490 ( .B(n1556), .A(n1557), .S(\C2334/net59912 ), .Y(n1555) );
  MUX2X1 U1491 ( .B(n1559), .A(n1560), .S(\C2334/net59514 ), .Y(n1558) );
  MUX2X1 U1492 ( .B(n1562), .A(n1563), .S(\C2334/net59912 ), .Y(n1561) );
  MUX2X1 U1493 ( .B(n1565), .A(n1566), .S(\C2334/net59912 ), .Y(n1564) );
  MUX2X1 U1494 ( .B(n1568), .A(n1569), .S(\C2334/net59912 ), .Y(n1567) );
  MUX2X1 U1495 ( .B(n1571), .A(n1572), .S(\C2334/net59912 ), .Y(n1570) );
  MUX2X1 U1496 ( .B(n1574), .A(n1575), .S(\C2334/net59514 ), .Y(n1573) );
  MUX2X1 U1497 ( .B(n1577), .A(n1578), .S(\C2334/net59910 ), .Y(n1576) );
  MUX2X1 U1498 ( .B(n1580), .A(n1581), .S(\C2334/net59910 ), .Y(n1579) );
  MUX2X1 U1499 ( .B(n1583), .A(n1584), .S(\C2334/net59910 ), .Y(n1582) );
  MUX2X1 U1500 ( .B(n1586), .A(n1587), .S(\C2334/net59910 ), .Y(n1585) );
  MUX2X1 U1501 ( .B(n1589), .A(n1590), .S(\C2334/net59514 ), .Y(n1588) );
  MUX2X1 U1502 ( .B(n1592), .A(n1593), .S(\C2334/net59910 ), .Y(n1591) );
  MUX2X1 U1503 ( .B(n1595), .A(n1596), .S(\C2334/net59910 ), .Y(n1594) );
  MUX2X1 U1504 ( .B(n1598), .A(n1599), .S(\C2334/net59910 ), .Y(n1597) );
  MUX2X1 U1505 ( .B(n1601), .A(n1602), .S(\C2334/net59910 ), .Y(n1600) );
  MUX2X1 U1506 ( .B(n1604), .A(n1605), .S(\C2334/net59514 ), .Y(n1603) );
  MUX2X1 U1507 ( .B(n1607), .A(n1608), .S(\C2334/net59910 ), .Y(n1606) );
  MUX2X1 U1508 ( .B(n1610), .A(n1611), .S(\C2334/net59910 ), .Y(n1609) );
  MUX2X1 U1509 ( .B(n1613), .A(n1614), .S(\C2334/net59910 ), .Y(n1612) );
  MUX2X1 U1510 ( .B(n1616), .A(n1617), .S(\C2334/net59910 ), .Y(n1615) );
  MUX2X1 U1511 ( .B(n1619), .A(n1620), .S(\C2334/net59512 ), .Y(n1618) );
  MUX2X1 U1512 ( .B(n1622), .A(n1623), .S(\C2334/net59908 ), .Y(n1621) );
  MUX2X1 U1513 ( .B(n1625), .A(n1626), .S(\C2334/net59908 ), .Y(n1624) );
  MUX2X1 U1514 ( .B(n1628), .A(n1629), .S(\C2334/net59908 ), .Y(n1627) );
  MUX2X1 U1515 ( .B(n1631), .A(n1632), .S(\C2334/net59908 ), .Y(n1630) );
  MUX2X1 U1516 ( .B(n1634), .A(n1635), .S(\C2334/net59512 ), .Y(n1633) );
  MUX2X1 U1517 ( .B(n1637), .A(n1638), .S(\C2334/net59908 ), .Y(n1636) );
  MUX2X1 U1518 ( .B(n1640), .A(n1641), .S(\C2334/net59908 ), .Y(n1639) );
  MUX2X1 U1519 ( .B(n1643), .A(n1644), .S(\C2334/net59908 ), .Y(n1642) );
  MUX2X1 U1520 ( .B(n1646), .A(n1647), .S(\C2334/net59908 ), .Y(n1645) );
  MUX2X1 U1521 ( .B(n1649), .A(n1650), .S(\C2334/net59512 ), .Y(n1648) );
  MUX2X1 U1522 ( .B(n1652), .A(n1653), .S(\C2334/net59908 ), .Y(n1651) );
  MUX2X1 U1523 ( .B(n1655), .A(n1656), .S(\C2334/net59908 ), .Y(n1654) );
  MUX2X1 U1524 ( .B(n1658), .A(n1659), .S(\C2334/net59908 ), .Y(n1657) );
  MUX2X1 U1525 ( .B(n1661), .A(n1662), .S(\C2334/net59908 ), .Y(n1660) );
  MUX2X1 U1526 ( .B(n1664), .A(n1665), .S(\C2334/net59512 ), .Y(n1663) );
  MUX2X1 U1527 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(\C2334/net60490 ), .Y(
        n1218) );
  MUX2X1 U1528 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(\C2334/net60490 ), .Y(
        n1217) );
  MUX2X1 U1529 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(\C2334/net60490 ), .Y(
        n1221) );
  MUX2X1 U1530 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(\C2334/net60490 ), .Y(
        n1220) );
  MUX2X1 U1531 ( .B(n1219), .A(n1216), .S(\C2334/net59710 ), .Y(n1230) );
  MUX2X1 U1532 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(\C2334/net60460 ), .Y(
        n1224) );
  MUX2X1 U1533 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n34), .Y(n1223) );
  MUX2X1 U1534 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(\C2334/net60472 ), .Y(
        n1227) );
  MUX2X1 U1535 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(\C2334/net60462 ), .Y(
        n1226) );
  MUX2X1 U1536 ( .B(n1225), .A(n1222), .S(\C2334/net59710 ), .Y(n1229) );
  MUX2X1 U1537 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(\C2334/net60460 ), .Y(
        n1233) );
  MUX2X1 U1538 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(\C2334/net60490 ), .Y(
        n1232) );
  MUX2X1 U1539 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(\C2334/net60472 ), .Y(
        n1236) );
  MUX2X1 U1540 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(\C2334/net60462 ), .Y(
        n1235) );
  MUX2X1 U1541 ( .B(n1234), .A(n1231), .S(\C2334/net59710 ), .Y(n1245) );
  MUX2X1 U1542 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(\C2334/net60470 ), .Y(
        n1239) );
  MUX2X1 U1543 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(\C2334/net60468 ), .Y(
        n1238) );
  MUX2X1 U1544 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(\C2334/net60490 ), .Y(
        n1242) );
  MUX2X1 U1545 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(\C2334/net60468 ), .Y(
        n1241) );
  MUX2X1 U1546 ( .B(n1240), .A(n1237), .S(\C2334/net59710 ), .Y(n1244) );
  MUX2X1 U1547 ( .B(n1243), .A(n1228), .S(\C2334/net59380 ), .Y(n1666) );
  MUX2X1 U1548 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(\C2334/net60490 ), .Y(
        n1248) );
  MUX2X1 U1549 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(\C2334/net60490 ), .Y(
        n1247) );
  MUX2X1 U1550 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(\C2334/net60490 ), .Y(
        n1251) );
  MUX2X1 U1551 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(\C2334/net60490 ), .Y(
        n1250) );
  MUX2X1 U1552 ( .B(n1249), .A(n1246), .S(\C2334/net59710 ), .Y(n1260) );
  MUX2X1 U1553 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(\C2334/net60490 ), .Y(
        n1254) );
  MUX2X1 U1554 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(\C2334/net60490 ), .Y(
        n1253) );
  MUX2X1 U1555 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(\C2334/net60490 ), .Y(
        n1257) );
  MUX2X1 U1556 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(\C2334/net60490 ), .Y(
        n1256) );
  MUX2X1 U1557 ( .B(n1255), .A(n1252), .S(\C2334/net59710 ), .Y(n1259) );
  MUX2X1 U1558 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(\C2334/net60490 ), .Y(
        n1263) );
  MUX2X1 U1559 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(\C2334/net60490 ), .Y(
        n1262) );
  MUX2X1 U1560 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(\C2334/net60490 ), .Y(
        n1266) );
  MUX2X1 U1561 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(\C2334/net60490 ), .Y(
        n1265) );
  MUX2X1 U1562 ( .B(n1264), .A(n1261), .S(\C2334/net59710 ), .Y(n1275) );
  MUX2X1 U1563 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(\C2334/net60484 ), .Y(
        n1269) );
  MUX2X1 U1564 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n34), .Y(n1268) );
  MUX2X1 U1565 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(\C2334/net60478 ), .Y(
        n1272) );
  MUX2X1 U1566 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(\C2334/net60474 ), .Y(
        n1271) );
  MUX2X1 U1567 ( .B(n1270), .A(n1267), .S(\C2334/net59710 ), .Y(n1274) );
  MUX2X1 U1568 ( .B(n1273), .A(n1258), .S(\C2334/net59380 ), .Y(n1667) );
  MUX2X1 U1569 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(\C2334/net60460 ), .Y(
        n1278) );
  MUX2X1 U1570 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(\C2334/net60462 ), .Y(
        n1277) );
  MUX2X1 U1571 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(\C2334/net60484 ), .Y(
        n1281) );
  MUX2X1 U1572 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(\C2334/net60470 ), .Y(
        n1280) );
  MUX2X1 U1573 ( .B(n1279), .A(n1276), .S(\C2334/net59710 ), .Y(n1290) );
  MUX2X1 U1574 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(\C2334/net60468 ), .Y(
        n1284) );
  MUX2X1 U1575 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(\C2334/net60472 ), .Y(
        n1283) );
  MUX2X1 U1576 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(\C2334/net60466 ), .Y(
        n1287) );
  MUX2X1 U1577 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n34), .Y(n1286) );
  MUX2X1 U1578 ( .B(n1285), .A(n1282), .S(\C2334/net59710 ), .Y(n1289) );
  MUX2X1 U1579 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(\C2334/net60470 ), .Y(
        n1293) );
  MUX2X1 U1580 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(\C2334/net60468 ), .Y(
        n1292) );
  MUX2X1 U1581 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(\C2334/net60476 ), .Y(
        n1296) );
  MUX2X1 U1582 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(\C2334/net60468 ), .Y(
        n1295) );
  MUX2X1 U1583 ( .B(n1294), .A(n1291), .S(\C2334/net59710 ), .Y(n1305) );
  MUX2X1 U1584 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(\C2334/net60460 ), .Y(
        n1299) );
  MUX2X1 U1585 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(\C2334/net60476 ), .Y(
        n1298) );
  MUX2X1 U1586 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(\C2334/net60464 ), .Y(
        n1302) );
  MUX2X1 U1587 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(\C2334/net60472 ), .Y(
        n1301) );
  MUX2X1 U1588 ( .B(n1300), .A(n1297), .S(\C2334/net59710 ), .Y(n1304) );
  MUX2X1 U1589 ( .B(n1303), .A(n1288), .S(\C2334/net59380 ), .Y(n1668) );
  MUX2X1 U1590 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(\C2334/net60466 ), .Y(
        n1308) );
  MUX2X1 U1591 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(\C2334/net60466 ), .Y(
        n1307) );
  MUX2X1 U1592 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(\C2334/net60464 ), .Y(
        n1311) );
  MUX2X1 U1593 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(\C2334/net60462 ), .Y(
        n1310) );
  MUX2X1 U1594 ( .B(n1309), .A(n1306), .S(\C2334/net59712 ), .Y(n1320) );
  MUX2X1 U1595 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(\C2334/net60484 ), .Y(
        n1314) );
  MUX2X1 U1596 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(\C2334/net60484 ), .Y(
        n1313) );
  MUX2X1 U1597 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(\C2334/net60484 ), .Y(
        n1317) );
  MUX2X1 U1598 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(\C2334/net60484 ), .Y(
        n1316) );
  MUX2X1 U1599 ( .B(n1315), .A(n1312), .S(\C2334/net59712 ), .Y(n1319) );
  MUX2X1 U1600 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(\C2334/net60484 ), .Y(
        n1323) );
  MUX2X1 U1601 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(\C2334/net60484 ), .Y(
        n1322) );
  MUX2X1 U1602 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(\C2334/net60484 ), .Y(
        n1326) );
  MUX2X1 U1603 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(\C2334/net60484 ), .Y(
        n1325) );
  MUX2X1 U1604 ( .B(n1324), .A(n1321), .S(\C2334/net59712 ), .Y(n1335) );
  MUX2X1 U1605 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(\C2334/net60484 ), .Y(
        n1329) );
  MUX2X1 U1606 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(\C2334/net60484 ), .Y(
        n1328) );
  MUX2X1 U1607 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(\C2334/net60484 ), .Y(
        n1332) );
  MUX2X1 U1608 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(\C2334/net60484 ), .Y(
        n1331) );
  MUX2X1 U1609 ( .B(n1330), .A(n1327), .S(\C2334/net59712 ), .Y(n1334) );
  MUX2X1 U1610 ( .B(n1333), .A(n1318), .S(\C2334/net59380 ), .Y(n1669) );
  MUX2X1 U1611 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(\C2334/net60472 ), .Y(
        n1338) );
  MUX2X1 U1612 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(\C2334/net60462 ), .Y(
        n1337) );
  MUX2X1 U1613 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(\C2334/net60462 ), .Y(
        n1341) );
  MUX2X1 U1614 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(\C2334/net60468 ), .Y(
        n1340) );
  MUX2X1 U1615 ( .B(n1339), .A(n1336), .S(\C2334/net59712 ), .Y(n1350) );
  MUX2X1 U1616 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(\C2334/net60470 ), .Y(
        n1344) );
  MUX2X1 U1617 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(\C2334/net60470 ), .Y(
        n1343) );
  MUX2X1 U1618 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(\C2334/net60460 ), .Y(
        n1347) );
  MUX2X1 U1619 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(\C2334/net60472 ), .Y(
        n1346) );
  MUX2X1 U1620 ( .B(n1345), .A(n1342), .S(\C2334/net59712 ), .Y(n1349) );
  MUX2X1 U1621 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(\C2334/net60478 ), .Y(
        n1353) );
  MUX2X1 U1622 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(\C2334/net60478 ), .Y(
        n1352) );
  MUX2X1 U1623 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(\C2334/net60478 ), .Y(
        n1356) );
  MUX2X1 U1624 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(\C2334/net60478 ), .Y(
        n1355) );
  MUX2X1 U1625 ( .B(n1354), .A(n1351), .S(\C2334/net59712 ), .Y(n1365) );
  MUX2X1 U1626 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(\C2334/net60478 ), .Y(
        n1359) );
  MUX2X1 U1627 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(\C2334/net60478 ), .Y(
        n1358) );
  MUX2X1 U1628 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(\C2334/net60478 ), .Y(
        n1362) );
  MUX2X1 U1629 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(\C2334/net60478 ), .Y(
        n1361) );
  MUX2X1 U1630 ( .B(n1360), .A(n1357), .S(\C2334/net59712 ), .Y(n1364) );
  MUX2X1 U1631 ( .B(n1363), .A(n1348), .S(\C2334/net59380 ), .Y(n1670) );
  MUX2X1 U1632 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(\C2334/net60478 ), .Y(
        n1368) );
  MUX2X1 U1633 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(\C2334/net60478 ), .Y(
        n1367) );
  MUX2X1 U1634 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(\C2334/net60478 ), .Y(
        n1371) );
  MUX2X1 U1635 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(\C2334/net60478 ), .Y(
        n1370) );
  MUX2X1 U1636 ( .B(n1369), .A(n1366), .S(\C2334/net59712 ), .Y(n1380) );
  MUX2X1 U1637 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(\C2334/net60476 ), .Y(
        n1374) );
  MUX2X1 U1638 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(\C2334/net60476 ), .Y(
        n1373) );
  MUX2X1 U1639 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(\C2334/net60476 ), .Y(
        n1377) );
  MUX2X1 U1640 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(\C2334/net60476 ), .Y(
        n1376) );
  MUX2X1 U1641 ( .B(n1375), .A(n1372), .S(\C2334/net59712 ), .Y(n1379) );
  MUX2X1 U1642 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(\C2334/net60476 ), .Y(
        n1383) );
  MUX2X1 U1643 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(\C2334/net60476 ), .Y(
        n1382) );
  MUX2X1 U1644 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(\C2334/net60476 ), .Y(
        n1386) );
  MUX2X1 U1645 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(\C2334/net60476 ), .Y(
        n1385) );
  MUX2X1 U1646 ( .B(n1384), .A(n1381), .S(\C2334/net59710 ), .Y(n1395) );
  MUX2X1 U1647 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(\C2334/net60476 ), .Y(
        n1389) );
  MUX2X1 U1648 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(\C2334/net60476 ), .Y(
        n1388) );
  MUX2X1 U1649 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(\C2334/net60476 ), .Y(
        n1392) );
  MUX2X1 U1650 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(\C2334/net60476 ), .Y(
        n1391) );
  MUX2X1 U1651 ( .B(n1390), .A(n1387), .S(\C2334/net59712 ), .Y(n1394) );
  MUX2X1 U1652 ( .B(n1393), .A(n1378), .S(\C2334/net59380 ), .Y(
        \C2334/net11884 ) );
  MUX2X1 U1653 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(\C2334/net60474 ), .Y(
        n1398) );
  MUX2X1 U1654 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(\C2334/net60474 ), .Y(
        n1397) );
  MUX2X1 U1655 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(\C2334/net60474 ), .Y(
        n1401) );
  MUX2X1 U1656 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(\C2334/net60474 ), .Y(
        n1400) );
  MUX2X1 U1657 ( .B(n1399), .A(n1396), .S(\C2334/net59710 ), .Y(n1410) );
  MUX2X1 U1658 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(\C2334/net60474 ), .Y(
        n1404) );
  MUX2X1 U1659 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(\C2334/net60474 ), .Y(
        n1403) );
  MUX2X1 U1660 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(\C2334/net60474 ), .Y(
        n1407) );
  MUX2X1 U1661 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(\C2334/net60474 ), .Y(
        n1406) );
  MUX2X1 U1662 ( .B(n1405), .A(n1402), .S(\C2334/net59710 ), .Y(n1409) );
  MUX2X1 U1663 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(\C2334/net60474 ), .Y(
        n1413) );
  MUX2X1 U1664 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(\C2334/net60474 ), .Y(
        n1412) );
  MUX2X1 U1665 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(\C2334/net60474 ), .Y(
        n1416) );
  MUX2X1 U1666 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(\C2334/net60474 ), .Y(
        n1415) );
  MUX2X1 U1667 ( .B(n1414), .A(n1411), .S(\C2334/net59710 ), .Y(n1425) );
  MUX2X1 U1668 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(\C2334/net60472 ), .Y(
        n1419) );
  MUX2X1 U1669 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(\C2334/net60472 ), .Y(
        n1418) );
  MUX2X1 U1670 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(\C2334/net60472 ), .Y(
        n1422) );
  MUX2X1 U1671 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(\C2334/net60472 ), .Y(
        n1421) );
  MUX2X1 U1672 ( .B(n1420), .A(n1417), .S(\C2334/net59710 ), .Y(n1424) );
  MUX2X1 U1673 ( .B(n1423), .A(n1408), .S(\C2334/net59380 ), .Y(n1671) );
  MUX2X1 U1674 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(\C2334/net60472 ), .Y(
        n1428) );
  MUX2X1 U1675 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(\C2334/net60472 ), .Y(
        n1427) );
  MUX2X1 U1676 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(\C2334/net60472 ), .Y(
        n1431) );
  MUX2X1 U1677 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(\C2334/net60472 ), .Y(
        n1430) );
  MUX2X1 U1678 ( .B(n1429), .A(n1426), .S(\C2334/net59712 ), .Y(n1440) );
  MUX2X1 U1679 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(\C2334/net60472 ), .Y(
        n1434) );
  MUX2X1 U1680 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(\C2334/net60472 ), .Y(
        n1433) );
  MUX2X1 U1681 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(\C2334/net60472 ), .Y(
        n1437) );
  MUX2X1 U1682 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(\C2334/net60472 ), .Y(
        n1436) );
  MUX2X1 U1683 ( .B(n1435), .A(n1432), .S(\C2334/net59712 ), .Y(n1439) );
  MUX2X1 U1684 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(\C2334/net60470 ), .Y(
        n1443) );
  MUX2X1 U1685 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(\C2334/net60470 ), .Y(
        n1442) );
  MUX2X1 U1686 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(\C2334/net60470 ), .Y(
        n1446) );
  MUX2X1 U1687 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(\C2334/net60470 ), .Y(
        n1445) );
  MUX2X1 U1688 ( .B(n1444), .A(n1441), .S(\C2334/net59712 ), .Y(n1455) );
  MUX2X1 U1689 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(\C2334/net60470 ), .Y(
        n1449) );
  MUX2X1 U1690 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(\C2334/net60470 ), .Y(
        n1448) );
  MUX2X1 U1691 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(\C2334/net60470 ), .Y(
        n1452) );
  MUX2X1 U1692 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(\C2334/net60470 ), .Y(
        n1451) );
  MUX2X1 U1693 ( .B(n1450), .A(n1447), .S(\C2334/net59712 ), .Y(n1454) );
  MUX2X1 U1694 ( .B(n1453), .A(n1438), .S(\C2334/net59380 ), .Y(n1672) );
  MUX2X1 U1695 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(\C2334/net60470 ), .Y(
        n1458) );
  MUX2X1 U1696 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(\C2334/net60470 ), .Y(
        n1457) );
  MUX2X1 U1697 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(\C2334/net60470 ), .Y(
        n1461) );
  MUX2X1 U1698 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(\C2334/net60470 ), .Y(
        n1460) );
  MUX2X1 U1699 ( .B(n1459), .A(n1456), .S(\C2334/net59716 ), .Y(n1470) );
  MUX2X1 U1700 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(\C2334/net60468 ), .Y(
        n1464) );
  MUX2X1 U1701 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(\C2334/net60468 ), .Y(
        n1463) );
  MUX2X1 U1702 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(\C2334/net60468 ), .Y(
        n1467) );
  MUX2X1 U1703 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(\C2334/net60468 ), .Y(
        n1466) );
  MUX2X1 U1704 ( .B(n1465), .A(n1462), .S(\C2334/net59716 ), .Y(n1469) );
  MUX2X1 U1705 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(\C2334/net60468 ), .Y(
        n1473) );
  MUX2X1 U1706 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(\C2334/net60468 ), .Y(
        n1472) );
  MUX2X1 U1707 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(\C2334/net60468 ), .Y(
        n1476) );
  MUX2X1 U1708 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(\C2334/net60468 ), .Y(
        n1475) );
  MUX2X1 U1709 ( .B(n1474), .A(n1471), .S(\C2334/net59716 ), .Y(n1485) );
  MUX2X1 U1710 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(\C2334/net60468 ), .Y(
        n1479) );
  MUX2X1 U1711 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(\C2334/net60468 ), .Y(
        n1478) );
  MUX2X1 U1712 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(\C2334/net60468 ), .Y(
        n1482) );
  MUX2X1 U1713 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(\C2334/net60468 ), .Y(
        n1481) );
  MUX2X1 U1714 ( .B(n1480), .A(n1477), .S(\C2334/net59716 ), .Y(n1484) );
  MUX2X1 U1715 ( .B(n1483), .A(n1468), .S(\C2334/net59380 ), .Y(n1673) );
  MUX2X1 U1716 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(\C2334/net60466 ), 
        .Y(n1488) );
  MUX2X1 U1717 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(\C2334/net60466 ), 
        .Y(n1487) );
  MUX2X1 U1718 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(\C2334/net60466 ), 
        .Y(n1491) );
  MUX2X1 U1719 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(\C2334/net60466 ), 
        .Y(n1490) );
  MUX2X1 U1720 ( .B(n1489), .A(n1486), .S(\C2334/net59716 ), .Y(n1500) );
  MUX2X1 U1721 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(\C2334/net60466 ), 
        .Y(n1494) );
  MUX2X1 U1722 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(\C2334/net60466 ), 
        .Y(n1493) );
  MUX2X1 U1723 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(\C2334/net60466 ), 
        .Y(n1497) );
  MUX2X1 U1724 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(\C2334/net60466 ), 
        .Y(n1496) );
  MUX2X1 U1725 ( .B(n1495), .A(n1492), .S(\C2334/net59716 ), .Y(n1499) );
  MUX2X1 U1726 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(\C2334/net60466 ), 
        .Y(n1503) );
  MUX2X1 U1727 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(\C2334/net60466 ), 
        .Y(n1502) );
  MUX2X1 U1728 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(\C2334/net60466 ), 
        .Y(n1506) );
  MUX2X1 U1729 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(\C2334/net60466 ), .Y(
        n1505) );
  MUX2X1 U1730 ( .B(n1504), .A(n1501), .S(\C2334/net59716 ), .Y(n1515) );
  MUX2X1 U1731 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(\C2334/net60464 ), .Y(
        n1509) );
  MUX2X1 U1732 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(\C2334/net60464 ), .Y(
        n1508) );
  MUX2X1 U1733 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(\C2334/net60464 ), .Y(
        n1512) );
  MUX2X1 U1734 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(\C2334/net60464 ), .Y(
        n1511) );
  MUX2X1 U1735 ( .B(n1510), .A(n1507), .S(\C2334/net59716 ), .Y(n1514) );
  MUX2X1 U1736 ( .B(n1513), .A(n1498), .S(\C2334/net59380 ), .Y(n1674) );
  MUX2X1 U1737 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(\C2334/net60464 ), 
        .Y(n1518) );
  MUX2X1 U1738 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(\C2334/net60464 ), 
        .Y(n1517) );
  MUX2X1 U1739 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(\C2334/net60464 ), 
        .Y(n1521) );
  MUX2X1 U1740 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(\C2334/net60464 ), 
        .Y(n1520) );
  MUX2X1 U1741 ( .B(n1519), .A(n1516), .S(\C2334/net59716 ), .Y(n1530) );
  MUX2X1 U1742 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(\C2334/net60464 ), 
        .Y(n1524) );
  MUX2X1 U1743 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(\C2334/net60464 ), 
        .Y(n1523) );
  MUX2X1 U1744 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(\C2334/net60464 ), 
        .Y(n1527) );
  MUX2X1 U1745 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(\C2334/net60464 ), 
        .Y(n1526) );
  MUX2X1 U1746 ( .B(n1525), .A(n1522), .S(\C2334/net59716 ), .Y(n1529) );
  MUX2X1 U1747 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(\C2334/net60462 ), 
        .Y(n1533) );
  MUX2X1 U1748 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(\C2334/net60462 ), 
        .Y(n1532) );
  MUX2X1 U1749 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(\C2334/net60462 ), 
        .Y(n1536) );
  MUX2X1 U1750 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(\C2334/net60462 ), .Y(
        n1535) );
  MUX2X1 U1751 ( .B(n1534), .A(n1531), .S(\C2334/net59716 ), .Y(n1545) );
  MUX2X1 U1752 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(\C2334/net60462 ), .Y(
        n1539) );
  MUX2X1 U1753 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(\C2334/net60462 ), .Y(
        n1538) );
  MUX2X1 U1754 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(\C2334/net60462 ), .Y(
        n1542) );
  MUX2X1 U1755 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(\C2334/net60462 ), .Y(
        n1541) );
  MUX2X1 U1756 ( .B(n1540), .A(n1537), .S(\C2334/net59716 ), .Y(n1544) );
  MUX2X1 U1757 ( .B(n1543), .A(n1528), .S(\C2334/net59380 ), .Y(n1675) );
  MUX2X1 U1758 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(\C2334/net60462 ), 
        .Y(n1548) );
  MUX2X1 U1759 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(\C2334/net60462 ), 
        .Y(n1547) );
  MUX2X1 U1760 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(\C2334/net60462 ), 
        .Y(n1551) );
  MUX2X1 U1761 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(\C2334/net60462 ), 
        .Y(n1550) );
  MUX2X1 U1762 ( .B(n1549), .A(n1546), .S(\C2334/net59718 ), .Y(n1560) );
  MUX2X1 U1763 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(\C2334/net60460 ), 
        .Y(n1554) );
  MUX2X1 U1764 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(\C2334/net60460 ), 
        .Y(n1553) );
  MUX2X1 U1765 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(\C2334/net60460 ), 
        .Y(n1557) );
  MUX2X1 U1766 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(\C2334/net60460 ), 
        .Y(n1556) );
  MUX2X1 U1767 ( .B(n1555), .A(n1552), .S(\C2334/net59718 ), .Y(n1559) );
  MUX2X1 U1768 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(\C2334/net60460 ), 
        .Y(n1563) );
  MUX2X1 U1769 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(\C2334/net60460 ), 
        .Y(n1562) );
  MUX2X1 U1770 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(\C2334/net60460 ), 
        .Y(n1566) );
  MUX2X1 U1771 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(\C2334/net60460 ), .Y(
        n1565) );
  MUX2X1 U1772 ( .B(n1564), .A(n1561), .S(\C2334/net59718 ), .Y(n1575) );
  MUX2X1 U1773 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(\C2334/net60460 ), .Y(
        n1569) );
  MUX2X1 U1774 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(\C2334/net60460 ), .Y(
        n1568) );
  MUX2X1 U1775 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(\C2334/net60460 ), .Y(
        n1572) );
  MUX2X1 U1776 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(\C2334/net60460 ), .Y(
        n1571) );
  MUX2X1 U1777 ( .B(n1570), .A(n1567), .S(\C2334/net59718 ), .Y(n1574) );
  MUX2X1 U1778 ( .B(n1573), .A(n1558), .S(\C2334/net59380 ), .Y(n1676) );
  MUX2X1 U1779 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(\C2334/net60470 ), 
        .Y(n1578) );
  MUX2X1 U1780 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(\C2334/net60468 ), 
        .Y(n1577) );
  MUX2X1 U1781 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(\C2334/net60470 ), 
        .Y(n1581) );
  MUX2X1 U1782 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(\C2334/net60468 ), 
        .Y(n1580) );
  MUX2X1 U1783 ( .B(n1579), .A(n1576), .S(\C2334/net59718 ), .Y(n1590) );
  MUX2X1 U1784 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n34), .Y(n1584) );
  MUX2X1 U1785 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(\C2334/net60462 ), 
        .Y(n1583) );
  MUX2X1 U1786 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(\C2334/net60472 ), 
        .Y(n1587) );
  MUX2X1 U1787 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(\C2334/net60470 ), 
        .Y(n1586) );
  MUX2X1 U1788 ( .B(n1585), .A(n1582), .S(\C2334/net59718 ), .Y(n1589) );
  MUX2X1 U1789 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(\C2334/net60462 ), 
        .Y(n1593) );
  MUX2X1 U1790 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(\C2334/net60460 ), 
        .Y(n1592) );
  MUX2X1 U1791 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(\C2334/net60468 ), 
        .Y(n1596) );
  MUX2X1 U1792 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(\C2334/net60460 ), .Y(
        n1595) );
  MUX2X1 U1793 ( .B(n1594), .A(n1591), .S(\C2334/net59718 ), .Y(n1605) );
  MUX2X1 U1794 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(\C2334/net60470 ), .Y(
        n1599) );
  MUX2X1 U1795 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(\C2334/net60462 ), .Y(
        n1598) );
  MUX2X1 U1796 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(\C2334/net60468 ), .Y(
        n1602) );
  MUX2X1 U1797 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(\C2334/net60470 ), .Y(
        n1601) );
  MUX2X1 U1798 ( .B(n1600), .A(n1597), .S(\C2334/net59718 ), .Y(n1604) );
  MUX2X1 U1799 ( .B(n1603), .A(n1588), .S(\C2334/net59380 ), .Y(n1677) );
  MUX2X1 U1800 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(\C2334/net60462 ), 
        .Y(n1608) );
  MUX2X1 U1801 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(\C2334/net60468 ), 
        .Y(n1607) );
  MUX2X1 U1802 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(\C2334/net60460 ), 
        .Y(n1611) );
  MUX2X1 U1803 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(\C2334/net60462 ), 
        .Y(n1610) );
  MUX2X1 U1804 ( .B(n1609), .A(n1606), .S(\C2334/net59718 ), .Y(n1620) );
  MUX2X1 U1805 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(\C2334/net60460 ), 
        .Y(n1614) );
  MUX2X1 U1806 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n34), .Y(n1613) );
  MUX2X1 U1807 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(\C2334/net60470 ), 
        .Y(n1617) );
  MUX2X1 U1808 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(\C2334/net60460 ), 
        .Y(n1616) );
  MUX2X1 U1809 ( .B(n1615), .A(n1612), .S(\C2334/net59718 ), .Y(n1619) );
  MUX2X1 U1810 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(\C2334/net60470 ), 
        .Y(n1623) );
  MUX2X1 U1811 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(\C2334/net60462 ), 
        .Y(n1622) );
  MUX2X1 U1812 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n34), .Y(n1626) );
  MUX2X1 U1813 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n34), .Y(n1625) );
  MUX2X1 U1814 ( .B(n1624), .A(n1621), .S(\C2334/net59718 ), .Y(n1635) );
  MUX2X1 U1815 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(\C2334/net60468 ), .Y(
        n1629) );
  MUX2X1 U1816 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(\C2334/net60460 ), .Y(
        n1628) );
  MUX2X1 U1817 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(\C2334/net60490 ), .Y(
        n1632) );
  MUX2X1 U1818 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(\C2334/net60468 ), .Y(
        n1631) );
  MUX2X1 U1819 ( .B(n1630), .A(n1627), .S(\C2334/net59718 ), .Y(n1634) );
  MUX2X1 U1820 ( .B(n1633), .A(n1618), .S(\C2334/net59380 ), .Y(n1678) );
  MUX2X1 U1821 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(\C2334/net60490 ), 
        .Y(n1638) );
  MUX2X1 U1822 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(\C2334/net60490 ), 
        .Y(n1637) );
  MUX2X1 U1823 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n34), .Y(n1641) );
  MUX2X1 U1824 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(\C2334/net60460 ), 
        .Y(n1640) );
  MUX2X1 U1825 ( .B(n1639), .A(n1636), .S(\C2334/net59718 ), .Y(n1650) );
  MUX2X1 U1826 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(\C2334/net60452 ), 
        .Y(n1644) );
  MUX2X1 U1827 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(\C2334/net60452 ), 
        .Y(n1643) );
  MUX2X1 U1828 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(\C2334/net60452 ), 
        .Y(n1647) );
  MUX2X1 U1829 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(\C2334/net60452 ), 
        .Y(n1646) );
  MUX2X1 U1830 ( .B(n1645), .A(n1642), .S(\C2334/net59716 ), .Y(n1649) );
  MUX2X1 U1831 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(\C2334/net60452 ), 
        .Y(n1653) );
  MUX2X1 U1832 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(\C2334/net60452 ), 
        .Y(n1652) );
  MUX2X1 U1833 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(\C2334/net60452 ), 
        .Y(n1656) );
  MUX2X1 U1834 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(\C2334/net60452 ), .Y(
        n1655) );
  MUX2X1 U1835 ( .B(n1654), .A(n1651), .S(\C2334/net59716 ), .Y(n1665) );
  MUX2X1 U1836 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(\C2334/net60452 ), .Y(
        n1659) );
  MUX2X1 U1837 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(\C2334/net60452 ), .Y(
        n1658) );
  MUX2X1 U1838 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(\C2334/net60452 ), .Y(
        n1662) );
  MUX2X1 U1839 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(\C2334/net60452 ), .Y(
        n1661) );
  MUX2X1 U1840 ( .B(n1660), .A(n1657), .S(\C2334/net59716 ), .Y(n1664) );
  MUX2X1 U1841 ( .B(n1663), .A(n1648), .S(\C2334/net59380 ), .Y(n1679) );
  BUFX2 U1842 ( .A(write), .Y(net65995) );
  INVX1 U1843 ( .A(N11), .Y(net60096) );
  INVX1 U1844 ( .A(N10), .Y(net60828) );
  INVX8 U1845 ( .A(n1779), .Y(n1776) );
  INVX8 U1846 ( .A(n1779), .Y(n1777) );
  INVX8 U1847 ( .A(n1779), .Y(n1778) );
  INVX8 U1848 ( .A(n1166), .Y(n1780) );
  INVX8 U1849 ( .A(n1167), .Y(n1781) );
  INVX8 U1850 ( .A(n1167), .Y(n1782) );
  INVX8 U1851 ( .A(n1168), .Y(n1783) );
  INVX8 U1852 ( .A(n1169), .Y(n1784) );
  INVX8 U1853 ( .A(n1170), .Y(n1785) );
  INVX8 U1854 ( .A(n1171), .Y(n1786) );
  INVX8 U1855 ( .A(n1171), .Y(n1787) );
  INVX8 U1856 ( .A(n1172), .Y(n1788) );
  INVX8 U1857 ( .A(n1173), .Y(n1789) );
  INVX8 U1858 ( .A(n70), .Y(n1790) );
  INVX8 U1859 ( .A(n70), .Y(n1791) );
  INVX8 U1860 ( .A(n72), .Y(n1792) );
  INVX8 U1861 ( .A(n72), .Y(n1793) );
  INVX8 U1862 ( .A(n74), .Y(n1794) );
  INVX8 U1863 ( .A(n74), .Y(n1795) );
  INVX8 U1864 ( .A(n76), .Y(n1796) );
  INVX8 U1865 ( .A(n76), .Y(n1797) );
  INVX8 U1866 ( .A(n80), .Y(n1798) );
  INVX8 U1867 ( .A(n80), .Y(n1799) );
  INVX8 U1868 ( .A(n82), .Y(n1800) );
  INVX8 U1869 ( .A(n82), .Y(n1801) );
  INVX8 U1870 ( .A(n99), .Y(n1802) );
  INVX8 U1871 ( .A(n99), .Y(n1803) );
  INVX8 U1872 ( .A(n101), .Y(n1804) );
  INVX8 U1873 ( .A(n101), .Y(n1805) );
endmodule


module memc_Size16_5 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n15, n17, n19, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41,
         n43, n45, n47, n48, n50, n52, n54, n56, n58, n60, n62, n64, n66, n68,
         n70, n72, n74, n76, n80, n82, n99, n101, n118, n120, n137, n139, n156,
         n158, n175, n177, n194, n196, n215, n217, n233, n235, n251, n253,
         n269, n271, n287, n289, n305, n307, n323, n325, n341, n343, n360,
         n362, n378, n380, n396, n398, n414, n416, n432, n434, n450, n452,
         n468, n470, n486, n488, n505, n507, n523, n525, n541, n543, n559,
         n561, n577, n579, n595, n597, n613, n615, n631, n633, n650, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1878), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1879), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1880), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1881), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1882), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1883), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1884), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1885), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1886), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1887), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1888), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1889), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1890), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1891), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1892), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1893), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1894), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1895), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1896), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1897), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1898), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1899), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1900), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1901), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1902), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1903), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1904), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1905), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1906), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1907), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1908), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1909), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1910), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1911), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1912), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1913), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1914), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1915), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1916), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1917), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1918), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1919), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1920), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1921), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1922), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1923), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1924), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1925), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1926), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1927), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1928), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1929), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1930), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1931), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1932), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1933), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1934), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1935), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1936), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1937), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1938), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1939), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1940), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1941), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1942), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1943), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1944), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1945), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1946), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1947), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1948), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1949), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1950), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1951), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1952), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1953), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1954), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1955), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1956), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1957), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1958), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1959), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1960), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1961), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1962), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1963), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1964), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1965), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1966), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1967), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1968), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1969), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1970), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1971), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1972), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1973), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1974), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1975), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1976), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1977), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1978), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1979), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1980), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1981), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1982), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1983), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1984), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1985), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1986), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1987), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1988), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1989), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1990), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1991), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1992), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1993), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1994), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1995), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1996), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1997), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1998), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1999), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2000), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2001), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2002), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2003), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2004), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2005), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2006), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2007), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2008), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2009), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2010), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2011), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2012), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2013), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2014), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2015), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2016), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2017), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2018), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2019), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2020), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2021), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2022), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2023), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2024), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2025), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2026), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2027), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2028), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2029), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2030), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2031), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2032), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2033), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2034), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2035), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2036), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2037), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2038), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2039), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2040), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2041), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2042), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2043), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2044), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2045), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2046), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2047), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2048), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2049), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2050), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2051), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2052), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2053), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2054), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2055), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2056), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2057), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2058), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2059), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2060), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2061), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2062), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2063), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2064), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2065), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2066), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2067), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2068), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2069), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2070), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2071), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2072), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2073), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2074), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2075), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2076), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2077), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2078), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2079), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2080), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2081), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2082), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2083), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2084), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2085), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2086), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2087), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2088), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2089), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2090), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2091), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2092), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2093), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2094), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2095), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2096), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2097), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2098), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2099), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2100), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2101), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2102), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2103), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2104), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2105), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2106), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2107), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2108), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2109), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2110), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2111), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2112), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2113), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2114), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2115), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2116), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2117), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2118), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2119), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2120), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2121), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2122), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2123), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2124), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2125), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2126), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2127), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2128), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2129), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2130), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2131), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2132), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2133), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2134), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2135), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2136), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2137), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2138), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2139), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2140), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2141), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2142), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2143), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2144), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2145), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2146), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2147), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2148), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2149), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2150), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2151), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2152), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2153), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2154), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2155), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2156), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2157), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2158), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2159), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2160), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2161), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2162), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2163), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2164), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2165), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2166), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2167), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2168), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2169), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2170), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2171), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2172), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2173), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2174), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2175), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2176), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2177), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2178), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2179), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2180), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2181), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2182), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2183), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2184), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2185), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2186), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2187), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2188), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2189), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2190), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2191), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2192), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2193), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2194), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2195), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2196), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2197), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2198), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2199), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2200), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2201), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2202), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2203), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2204), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2205), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2214), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2215), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2216), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2217), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2218), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2219), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2220), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2221), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2222), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2223), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2224), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2225), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2226), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2227), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2228), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2229), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2230), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2231), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2232), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2233), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2234), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2235), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2236), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2237), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2238), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2239), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2240), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2241), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2242), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2243), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2244), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2245), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2246), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2247), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2248), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2249), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2250), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2251), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2252), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2253), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2254), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2255), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2256), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2257), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2258), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2259), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2260), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2261), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2262), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2263), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2264), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2265), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2266), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2267), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2268), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2269), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2270), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2271), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2272), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2273), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2274), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2275), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2276), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2277), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2278), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2279), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2280), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2281), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2282), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2283), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2284), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2285), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2286), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2287), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2288), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2289), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2290), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2291), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2292), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2293), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2294), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2295), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2296), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2297), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2298), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2299), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2300), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2301), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2302), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2303), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2304), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2305), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2306), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2307), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2308), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2309), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2310), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2311), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2312), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2313), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2314), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2315), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2316), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2317), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2318), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2319), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2320), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2321), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2322), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2323), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2324), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2325), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2326), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2327), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2328), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2329), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2330), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2331), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2332), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2333), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2334), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2335), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2336), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2337), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2338), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2339), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2340), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2341), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2342), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2343), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2344), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2345), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2346), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2347), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2348), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2349), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2350), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2351), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2352), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2353), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2354), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2355), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2356), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2357), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2358), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2359), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2360), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2361), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2362), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2363), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2364), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2365), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2366), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2367), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2368), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2369), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2370), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2371), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2372), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2373), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2374), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2375), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2376), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2377), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2378), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2379), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2380), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2381), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2382), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2383), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2384), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2385), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2386), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2387), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2388), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2389), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(write), .B(n1873), .Y(n2899) );
  OAI21X1 U61 ( .A(n1825), .B(n1861), .C(n2915), .Y(n2389) );
  NAND2X1 U62 ( .A(\mem<31><0> ), .B(n1827), .Y(n2915) );
  OAI21X1 U63 ( .A(n1825), .B(n1858), .C(n2914), .Y(n2388) );
  NAND2X1 U64 ( .A(\mem<31><1> ), .B(n1827), .Y(n2914) );
  OAI21X1 U65 ( .A(n1825), .B(n1855), .C(n2913), .Y(n2387) );
  NAND2X1 U66 ( .A(\mem<31><2> ), .B(n1827), .Y(n2913) );
  OAI21X1 U67 ( .A(n1825), .B(n1852), .C(n2912), .Y(n2386) );
  NAND2X1 U68 ( .A(\mem<31><3> ), .B(n1827), .Y(n2912) );
  OAI21X1 U69 ( .A(n1825), .B(n1849), .C(n2911), .Y(n2385) );
  NAND2X1 U70 ( .A(\mem<31><4> ), .B(n1827), .Y(n2911) );
  OAI21X1 U71 ( .A(n1825), .B(n1846), .C(n2910), .Y(n2384) );
  NAND2X1 U72 ( .A(\mem<31><5> ), .B(n1827), .Y(n2910) );
  OAI21X1 U73 ( .A(n1825), .B(n1843), .C(n2909), .Y(n2383) );
  NAND2X1 U74 ( .A(\mem<31><6> ), .B(n1827), .Y(n2909) );
  OAI21X1 U75 ( .A(n1825), .B(n1840), .C(n2908), .Y(n2382) );
  NAND2X1 U76 ( .A(\mem<31><7> ), .B(n1827), .Y(n2908) );
  OAI21X1 U77 ( .A(n1825), .B(n1839), .C(n2907), .Y(n2381) );
  NAND2X1 U78 ( .A(\mem<31><8> ), .B(n1826), .Y(n2907) );
  OAI21X1 U79 ( .A(n1825), .B(n1838), .C(n2906), .Y(n2380) );
  NAND2X1 U80 ( .A(\mem<31><9> ), .B(n1826), .Y(n2906) );
  OAI21X1 U81 ( .A(n1825), .B(n1837), .C(n2905), .Y(n2379) );
  NAND2X1 U82 ( .A(\mem<31><10> ), .B(n1826), .Y(n2905) );
  OAI21X1 U83 ( .A(n1825), .B(n1836), .C(n2904), .Y(n2378) );
  NAND2X1 U84 ( .A(\mem<31><11> ), .B(n1826), .Y(n2904) );
  OAI21X1 U85 ( .A(n1825), .B(n1835), .C(n2903), .Y(n2377) );
  NAND2X1 U86 ( .A(\mem<31><12> ), .B(n1826), .Y(n2903) );
  OAI21X1 U87 ( .A(n1825), .B(n1834), .C(n2902), .Y(n2376) );
  NAND2X1 U88 ( .A(\mem<31><13> ), .B(n1826), .Y(n2902) );
  OAI21X1 U89 ( .A(n1825), .B(n1833), .C(n2901), .Y(n2375) );
  NAND2X1 U90 ( .A(\mem<31><14> ), .B(n1826), .Y(n2901) );
  OAI21X1 U91 ( .A(n1825), .B(n1832), .C(n2900), .Y(n2374) );
  NAND2X1 U92 ( .A(\mem<31><15> ), .B(n1826), .Y(n2900) );
  OAI21X1 U95 ( .A(n1861), .B(n1822), .C(n2897), .Y(n2373) );
  NAND2X1 U96 ( .A(\mem<30><0> ), .B(n1824), .Y(n2897) );
  OAI21X1 U97 ( .A(n1858), .B(n1822), .C(n2896), .Y(n2372) );
  NAND2X1 U98 ( .A(\mem<30><1> ), .B(n1824), .Y(n2896) );
  OAI21X1 U99 ( .A(n1855), .B(n1822), .C(n2895), .Y(n2371) );
  NAND2X1 U100 ( .A(\mem<30><2> ), .B(n1824), .Y(n2895) );
  OAI21X1 U101 ( .A(n1852), .B(n1822), .C(n2894), .Y(n2370) );
  NAND2X1 U102 ( .A(\mem<30><3> ), .B(n1824), .Y(n2894) );
  OAI21X1 U103 ( .A(n1849), .B(n1822), .C(n2893), .Y(n2369) );
  NAND2X1 U104 ( .A(\mem<30><4> ), .B(n1824), .Y(n2893) );
  OAI21X1 U105 ( .A(n1846), .B(n1822), .C(n2892), .Y(n2368) );
  NAND2X1 U106 ( .A(\mem<30><5> ), .B(n1824), .Y(n2892) );
  OAI21X1 U107 ( .A(n1843), .B(n1822), .C(n2891), .Y(n2367) );
  NAND2X1 U108 ( .A(\mem<30><6> ), .B(n1824), .Y(n2891) );
  OAI21X1 U109 ( .A(n1840), .B(n1822), .C(n2890), .Y(n2366) );
  NAND2X1 U110 ( .A(\mem<30><7> ), .B(n1824), .Y(n2890) );
  OAI21X1 U111 ( .A(n1839), .B(n1822), .C(n2889), .Y(n2365) );
  NAND2X1 U112 ( .A(\mem<30><8> ), .B(n1823), .Y(n2889) );
  OAI21X1 U113 ( .A(n1838), .B(n1822), .C(n2888), .Y(n2364) );
  NAND2X1 U114 ( .A(\mem<30><9> ), .B(n1823), .Y(n2888) );
  OAI21X1 U115 ( .A(n1837), .B(n1822), .C(n2887), .Y(n2363) );
  NAND2X1 U116 ( .A(\mem<30><10> ), .B(n1823), .Y(n2887) );
  OAI21X1 U117 ( .A(n1836), .B(n1822), .C(n2886), .Y(n2362) );
  NAND2X1 U118 ( .A(\mem<30><11> ), .B(n1823), .Y(n2886) );
  OAI21X1 U119 ( .A(n1835), .B(n1822), .C(n2885), .Y(n2361) );
  NAND2X1 U120 ( .A(\mem<30><12> ), .B(n1823), .Y(n2885) );
  OAI21X1 U121 ( .A(n1834), .B(n1822), .C(n2884), .Y(n2360) );
  NAND2X1 U122 ( .A(\mem<30><13> ), .B(n1823), .Y(n2884) );
  OAI21X1 U123 ( .A(n1833), .B(n1822), .C(n2883), .Y(n2359) );
  NAND2X1 U124 ( .A(\mem<30><14> ), .B(n1823), .Y(n2883) );
  OAI21X1 U125 ( .A(n1832), .B(n1822), .C(n2882), .Y(n2358) );
  NAND2X1 U126 ( .A(\mem<30><15> ), .B(n1823), .Y(n2882) );
  OAI21X1 U129 ( .A(n1861), .B(n1819), .C(n2880), .Y(n2357) );
  NAND2X1 U130 ( .A(\mem<29><0> ), .B(n1821), .Y(n2880) );
  OAI21X1 U131 ( .A(n1858), .B(n1819), .C(n2879), .Y(n2356) );
  NAND2X1 U132 ( .A(\mem<29><1> ), .B(n1821), .Y(n2879) );
  OAI21X1 U133 ( .A(n1855), .B(n1819), .C(n2878), .Y(n2355) );
  NAND2X1 U134 ( .A(\mem<29><2> ), .B(n1821), .Y(n2878) );
  OAI21X1 U135 ( .A(n1852), .B(n1819), .C(n2877), .Y(n2354) );
  NAND2X1 U136 ( .A(\mem<29><3> ), .B(n1821), .Y(n2877) );
  OAI21X1 U137 ( .A(n1849), .B(n1819), .C(n2876), .Y(n2353) );
  NAND2X1 U138 ( .A(\mem<29><4> ), .B(n1821), .Y(n2876) );
  OAI21X1 U139 ( .A(n1846), .B(n1819), .C(n2875), .Y(n2352) );
  NAND2X1 U140 ( .A(\mem<29><5> ), .B(n1821), .Y(n2875) );
  OAI21X1 U141 ( .A(n1843), .B(n1819), .C(n2874), .Y(n2351) );
  NAND2X1 U142 ( .A(\mem<29><6> ), .B(n1821), .Y(n2874) );
  OAI21X1 U143 ( .A(n1840), .B(n1819), .C(n2873), .Y(n2350) );
  NAND2X1 U144 ( .A(\mem<29><7> ), .B(n1821), .Y(n2873) );
  OAI21X1 U145 ( .A(n1839), .B(n1819), .C(n2872), .Y(n2349) );
  NAND2X1 U146 ( .A(\mem<29><8> ), .B(n1820), .Y(n2872) );
  OAI21X1 U147 ( .A(n1838), .B(n1819), .C(n2871), .Y(n2348) );
  NAND2X1 U148 ( .A(\mem<29><9> ), .B(n1820), .Y(n2871) );
  OAI21X1 U149 ( .A(n1837), .B(n1819), .C(n2870), .Y(n2347) );
  NAND2X1 U150 ( .A(\mem<29><10> ), .B(n1820), .Y(n2870) );
  OAI21X1 U151 ( .A(n1836), .B(n1819), .C(n2869), .Y(n2346) );
  NAND2X1 U152 ( .A(\mem<29><11> ), .B(n1820), .Y(n2869) );
  OAI21X1 U153 ( .A(n1835), .B(n1819), .C(n2868), .Y(n2345) );
  NAND2X1 U154 ( .A(\mem<29><12> ), .B(n1820), .Y(n2868) );
  OAI21X1 U155 ( .A(n1834), .B(n1819), .C(n2867), .Y(n2344) );
  NAND2X1 U156 ( .A(\mem<29><13> ), .B(n1820), .Y(n2867) );
  OAI21X1 U157 ( .A(n1833), .B(n1819), .C(n2866), .Y(n2343) );
  NAND2X1 U158 ( .A(\mem<29><14> ), .B(n1820), .Y(n2866) );
  OAI21X1 U159 ( .A(n1832), .B(n1819), .C(n2865), .Y(n2342) );
  NAND2X1 U160 ( .A(\mem<29><15> ), .B(n1820), .Y(n2865) );
  OAI21X1 U163 ( .A(n1861), .B(n1816), .C(n2863), .Y(n2341) );
  NAND2X1 U164 ( .A(\mem<28><0> ), .B(n1818), .Y(n2863) );
  OAI21X1 U165 ( .A(n1858), .B(n1816), .C(n2862), .Y(n2340) );
  NAND2X1 U166 ( .A(\mem<28><1> ), .B(n1818), .Y(n2862) );
  OAI21X1 U167 ( .A(n1855), .B(n1816), .C(n2861), .Y(n2339) );
  NAND2X1 U168 ( .A(\mem<28><2> ), .B(n1818), .Y(n2861) );
  OAI21X1 U169 ( .A(n1852), .B(n1816), .C(n2860), .Y(n2338) );
  NAND2X1 U170 ( .A(\mem<28><3> ), .B(n1818), .Y(n2860) );
  OAI21X1 U171 ( .A(n1849), .B(n1816), .C(n2859), .Y(n2337) );
  NAND2X1 U172 ( .A(\mem<28><4> ), .B(n1818), .Y(n2859) );
  OAI21X1 U173 ( .A(n1846), .B(n1816), .C(n2858), .Y(n2336) );
  NAND2X1 U174 ( .A(\mem<28><5> ), .B(n1818), .Y(n2858) );
  OAI21X1 U175 ( .A(n1843), .B(n1816), .C(n2857), .Y(n2335) );
  NAND2X1 U176 ( .A(\mem<28><6> ), .B(n1818), .Y(n2857) );
  OAI21X1 U177 ( .A(n1840), .B(n1816), .C(n2856), .Y(n2334) );
  NAND2X1 U178 ( .A(\mem<28><7> ), .B(n1818), .Y(n2856) );
  OAI21X1 U179 ( .A(n1839), .B(n1816), .C(n2855), .Y(n2333) );
  NAND2X1 U180 ( .A(\mem<28><8> ), .B(n1817), .Y(n2855) );
  OAI21X1 U181 ( .A(n1838), .B(n1816), .C(n2854), .Y(n2332) );
  NAND2X1 U182 ( .A(\mem<28><9> ), .B(n1817), .Y(n2854) );
  OAI21X1 U183 ( .A(n1837), .B(n1816), .C(n2853), .Y(n2331) );
  NAND2X1 U184 ( .A(\mem<28><10> ), .B(n1817), .Y(n2853) );
  OAI21X1 U185 ( .A(n1836), .B(n1816), .C(n2852), .Y(n2330) );
  NAND2X1 U186 ( .A(\mem<28><11> ), .B(n1817), .Y(n2852) );
  OAI21X1 U187 ( .A(n1835), .B(n1816), .C(n2851), .Y(n2329) );
  NAND2X1 U188 ( .A(\mem<28><12> ), .B(n1817), .Y(n2851) );
  OAI21X1 U189 ( .A(n1834), .B(n1816), .C(n2850), .Y(n2328) );
  NAND2X1 U190 ( .A(\mem<28><13> ), .B(n1817), .Y(n2850) );
  OAI21X1 U191 ( .A(n1833), .B(n1816), .C(n2849), .Y(n2327) );
  NAND2X1 U192 ( .A(\mem<28><14> ), .B(n1817), .Y(n2849) );
  OAI21X1 U193 ( .A(n1832), .B(n1816), .C(n2848), .Y(n2326) );
  NAND2X1 U194 ( .A(\mem<28><15> ), .B(n1817), .Y(n2848) );
  OAI21X1 U197 ( .A(n1861), .B(n1813), .C(n2846), .Y(n2325) );
  NAND2X1 U198 ( .A(\mem<27><0> ), .B(n1815), .Y(n2846) );
  OAI21X1 U199 ( .A(n1858), .B(n1813), .C(n2845), .Y(n2324) );
  NAND2X1 U200 ( .A(\mem<27><1> ), .B(n1815), .Y(n2845) );
  OAI21X1 U201 ( .A(n1855), .B(n1813), .C(n2844), .Y(n2323) );
  NAND2X1 U202 ( .A(\mem<27><2> ), .B(n1815), .Y(n2844) );
  OAI21X1 U203 ( .A(n1852), .B(n1813), .C(n2843), .Y(n2322) );
  NAND2X1 U204 ( .A(\mem<27><3> ), .B(n1815), .Y(n2843) );
  OAI21X1 U205 ( .A(n1849), .B(n1813), .C(n2842), .Y(n2321) );
  NAND2X1 U206 ( .A(\mem<27><4> ), .B(n1815), .Y(n2842) );
  OAI21X1 U207 ( .A(n1846), .B(n1813), .C(n2841), .Y(n2320) );
  NAND2X1 U208 ( .A(\mem<27><5> ), .B(n1815), .Y(n2841) );
  OAI21X1 U209 ( .A(n1843), .B(n1813), .C(n2840), .Y(n2319) );
  NAND2X1 U210 ( .A(\mem<27><6> ), .B(n1815), .Y(n2840) );
  OAI21X1 U211 ( .A(n1840), .B(n1813), .C(n2839), .Y(n2318) );
  NAND2X1 U212 ( .A(\mem<27><7> ), .B(n1815), .Y(n2839) );
  OAI21X1 U213 ( .A(n1839), .B(n1813), .C(n2838), .Y(n2317) );
  NAND2X1 U214 ( .A(\mem<27><8> ), .B(n1814), .Y(n2838) );
  OAI21X1 U215 ( .A(n1838), .B(n1813), .C(n2837), .Y(n2316) );
  NAND2X1 U216 ( .A(\mem<27><9> ), .B(n1814), .Y(n2837) );
  OAI21X1 U217 ( .A(n1837), .B(n1813), .C(n2836), .Y(n2315) );
  NAND2X1 U218 ( .A(\mem<27><10> ), .B(n1814), .Y(n2836) );
  OAI21X1 U219 ( .A(n1836), .B(n1813), .C(n2835), .Y(n2314) );
  NAND2X1 U220 ( .A(\mem<27><11> ), .B(n1814), .Y(n2835) );
  OAI21X1 U221 ( .A(n1835), .B(n1813), .C(n2834), .Y(n2313) );
  NAND2X1 U222 ( .A(\mem<27><12> ), .B(n1814), .Y(n2834) );
  OAI21X1 U223 ( .A(n1834), .B(n1813), .C(n2833), .Y(n2312) );
  NAND2X1 U224 ( .A(\mem<27><13> ), .B(n1814), .Y(n2833) );
  OAI21X1 U225 ( .A(n1833), .B(n1813), .C(n2832), .Y(n2311) );
  NAND2X1 U226 ( .A(\mem<27><14> ), .B(n1814), .Y(n2832) );
  OAI21X1 U227 ( .A(n1832), .B(n1813), .C(n2831), .Y(n2310) );
  NAND2X1 U228 ( .A(\mem<27><15> ), .B(n1814), .Y(n2831) );
  OAI21X1 U231 ( .A(n1861), .B(n1810), .C(n2829), .Y(n2309) );
  NAND2X1 U232 ( .A(\mem<26><0> ), .B(n1812), .Y(n2829) );
  OAI21X1 U233 ( .A(n1858), .B(n1810), .C(n2828), .Y(n2308) );
  NAND2X1 U234 ( .A(\mem<26><1> ), .B(n1812), .Y(n2828) );
  OAI21X1 U235 ( .A(n1855), .B(n1810), .C(n2827), .Y(n2307) );
  NAND2X1 U236 ( .A(\mem<26><2> ), .B(n1812), .Y(n2827) );
  OAI21X1 U237 ( .A(n1852), .B(n1810), .C(n2826), .Y(n2306) );
  NAND2X1 U238 ( .A(\mem<26><3> ), .B(n1812), .Y(n2826) );
  OAI21X1 U239 ( .A(n1849), .B(n1810), .C(n2825), .Y(n2305) );
  NAND2X1 U240 ( .A(\mem<26><4> ), .B(n1812), .Y(n2825) );
  OAI21X1 U241 ( .A(n1846), .B(n1810), .C(n2824), .Y(n2304) );
  NAND2X1 U242 ( .A(\mem<26><5> ), .B(n1812), .Y(n2824) );
  OAI21X1 U243 ( .A(n1843), .B(n1810), .C(n2823), .Y(n2303) );
  NAND2X1 U244 ( .A(\mem<26><6> ), .B(n1812), .Y(n2823) );
  OAI21X1 U245 ( .A(n1840), .B(n1810), .C(n2822), .Y(n2302) );
  NAND2X1 U246 ( .A(\mem<26><7> ), .B(n1812), .Y(n2822) );
  OAI21X1 U247 ( .A(n1839), .B(n1810), .C(n2821), .Y(n2301) );
  NAND2X1 U248 ( .A(\mem<26><8> ), .B(n1811), .Y(n2821) );
  OAI21X1 U249 ( .A(n1838), .B(n1810), .C(n2820), .Y(n2300) );
  NAND2X1 U250 ( .A(\mem<26><9> ), .B(n1811), .Y(n2820) );
  OAI21X1 U251 ( .A(n1837), .B(n1810), .C(n2819), .Y(n2299) );
  NAND2X1 U252 ( .A(\mem<26><10> ), .B(n1811), .Y(n2819) );
  OAI21X1 U253 ( .A(n1836), .B(n1810), .C(n2818), .Y(n2298) );
  NAND2X1 U254 ( .A(\mem<26><11> ), .B(n1811), .Y(n2818) );
  OAI21X1 U255 ( .A(n1835), .B(n1810), .C(n2817), .Y(n2297) );
  NAND2X1 U256 ( .A(\mem<26><12> ), .B(n1811), .Y(n2817) );
  OAI21X1 U257 ( .A(n1834), .B(n1810), .C(n2816), .Y(n2296) );
  NAND2X1 U258 ( .A(\mem<26><13> ), .B(n1811), .Y(n2816) );
  OAI21X1 U259 ( .A(n1833), .B(n1810), .C(n2815), .Y(n2295) );
  NAND2X1 U260 ( .A(\mem<26><14> ), .B(n1811), .Y(n2815) );
  OAI21X1 U261 ( .A(n1832), .B(n1810), .C(n2814), .Y(n2294) );
  NAND2X1 U262 ( .A(\mem<26><15> ), .B(n1811), .Y(n2814) );
  OAI21X1 U265 ( .A(n1861), .B(n1807), .C(n2812), .Y(n2293) );
  NAND2X1 U266 ( .A(\mem<25><0> ), .B(n1809), .Y(n2812) );
  OAI21X1 U267 ( .A(n1858), .B(n1807), .C(n2811), .Y(n2292) );
  NAND2X1 U268 ( .A(\mem<25><1> ), .B(n1809), .Y(n2811) );
  OAI21X1 U269 ( .A(n1855), .B(n1807), .C(n2810), .Y(n2291) );
  NAND2X1 U270 ( .A(\mem<25><2> ), .B(n1809), .Y(n2810) );
  OAI21X1 U271 ( .A(n1852), .B(n1807), .C(n2809), .Y(n2290) );
  NAND2X1 U272 ( .A(\mem<25><3> ), .B(n1809), .Y(n2809) );
  OAI21X1 U273 ( .A(n1849), .B(n1807), .C(n2808), .Y(n2289) );
  NAND2X1 U274 ( .A(\mem<25><4> ), .B(n1809), .Y(n2808) );
  OAI21X1 U275 ( .A(n1846), .B(n1807), .C(n2807), .Y(n2288) );
  NAND2X1 U276 ( .A(\mem<25><5> ), .B(n1809), .Y(n2807) );
  OAI21X1 U277 ( .A(n1843), .B(n1807), .C(n2806), .Y(n2287) );
  NAND2X1 U278 ( .A(\mem<25><6> ), .B(n1809), .Y(n2806) );
  OAI21X1 U279 ( .A(n1840), .B(n1807), .C(n2805), .Y(n2286) );
  NAND2X1 U280 ( .A(\mem<25><7> ), .B(n1809), .Y(n2805) );
  OAI21X1 U281 ( .A(n1839), .B(n1807), .C(n2804), .Y(n2285) );
  NAND2X1 U282 ( .A(\mem<25><8> ), .B(n1808), .Y(n2804) );
  OAI21X1 U283 ( .A(n1838), .B(n1807), .C(n2803), .Y(n2284) );
  NAND2X1 U284 ( .A(\mem<25><9> ), .B(n1808), .Y(n2803) );
  OAI21X1 U285 ( .A(n1837), .B(n1807), .C(n2802), .Y(n2283) );
  NAND2X1 U286 ( .A(\mem<25><10> ), .B(n1808), .Y(n2802) );
  OAI21X1 U287 ( .A(n1836), .B(n1807), .C(n2801), .Y(n2282) );
  NAND2X1 U288 ( .A(\mem<25><11> ), .B(n1808), .Y(n2801) );
  OAI21X1 U289 ( .A(n1835), .B(n1807), .C(n2800), .Y(n2281) );
  NAND2X1 U290 ( .A(\mem<25><12> ), .B(n1808), .Y(n2800) );
  OAI21X1 U291 ( .A(n1834), .B(n1807), .C(n2799), .Y(n2280) );
  NAND2X1 U292 ( .A(\mem<25><13> ), .B(n1808), .Y(n2799) );
  OAI21X1 U293 ( .A(n1833), .B(n1807), .C(n2798), .Y(n2279) );
  NAND2X1 U294 ( .A(\mem<25><14> ), .B(n1808), .Y(n2798) );
  OAI21X1 U295 ( .A(n1832), .B(n1807), .C(n2797), .Y(n2278) );
  NAND2X1 U296 ( .A(\mem<25><15> ), .B(n1808), .Y(n2797) );
  OAI21X1 U299 ( .A(n1861), .B(n1804), .C(n2795), .Y(n2277) );
  NAND2X1 U300 ( .A(\mem<24><0> ), .B(n1806), .Y(n2795) );
  OAI21X1 U301 ( .A(n1858), .B(n1804), .C(n2794), .Y(n2276) );
  NAND2X1 U302 ( .A(\mem<24><1> ), .B(n1806), .Y(n2794) );
  OAI21X1 U303 ( .A(n1855), .B(n1804), .C(n2793), .Y(n2275) );
  NAND2X1 U304 ( .A(\mem<24><2> ), .B(n1806), .Y(n2793) );
  OAI21X1 U305 ( .A(n1852), .B(n1804), .C(n2792), .Y(n2274) );
  NAND2X1 U306 ( .A(\mem<24><3> ), .B(n1806), .Y(n2792) );
  OAI21X1 U307 ( .A(n1849), .B(n1804), .C(n2791), .Y(n2273) );
  NAND2X1 U308 ( .A(\mem<24><4> ), .B(n1806), .Y(n2791) );
  OAI21X1 U309 ( .A(n1846), .B(n1804), .C(n2790), .Y(n2272) );
  NAND2X1 U310 ( .A(\mem<24><5> ), .B(n1806), .Y(n2790) );
  OAI21X1 U311 ( .A(n1843), .B(n1804), .C(n2789), .Y(n2271) );
  NAND2X1 U312 ( .A(\mem<24><6> ), .B(n1806), .Y(n2789) );
  OAI21X1 U313 ( .A(n1840), .B(n1804), .C(n2788), .Y(n2270) );
  NAND2X1 U314 ( .A(\mem<24><7> ), .B(n1806), .Y(n2788) );
  OAI21X1 U315 ( .A(n1839), .B(n1804), .C(n2787), .Y(n2269) );
  NAND2X1 U316 ( .A(\mem<24><8> ), .B(n1805), .Y(n2787) );
  OAI21X1 U317 ( .A(n1838), .B(n1804), .C(n2786), .Y(n2268) );
  NAND2X1 U318 ( .A(\mem<24><9> ), .B(n1805), .Y(n2786) );
  OAI21X1 U319 ( .A(n1837), .B(n1804), .C(n2785), .Y(n2267) );
  NAND2X1 U320 ( .A(\mem<24><10> ), .B(n1805), .Y(n2785) );
  OAI21X1 U321 ( .A(n1836), .B(n1804), .C(n2784), .Y(n2266) );
  NAND2X1 U322 ( .A(\mem<24><11> ), .B(n1805), .Y(n2784) );
  OAI21X1 U323 ( .A(n1835), .B(n1804), .C(n2783), .Y(n2265) );
  NAND2X1 U324 ( .A(\mem<24><12> ), .B(n1805), .Y(n2783) );
  OAI21X1 U325 ( .A(n1834), .B(n1804), .C(n2782), .Y(n2264) );
  NAND2X1 U326 ( .A(\mem<24><13> ), .B(n1805), .Y(n2782) );
  OAI21X1 U327 ( .A(n1833), .B(n1804), .C(n2781), .Y(n2263) );
  NAND2X1 U328 ( .A(\mem<24><14> ), .B(n1805), .Y(n2781) );
  OAI21X1 U329 ( .A(n1832), .B(n1804), .C(n2780), .Y(n2262) );
  NAND2X1 U330 ( .A(\mem<24><15> ), .B(n1805), .Y(n2780) );
  NAND3X1 U333 ( .A(n1870), .B(n2777), .C(N14), .Y(n2778) );
  OAI21X1 U334 ( .A(n1861), .B(n1801), .C(n2776), .Y(n2261) );
  NAND2X1 U335 ( .A(\mem<23><0> ), .B(n1803), .Y(n2776) );
  OAI21X1 U336 ( .A(n1858), .B(n1801), .C(n2775), .Y(n2260) );
  NAND2X1 U337 ( .A(\mem<23><1> ), .B(n1803), .Y(n2775) );
  OAI21X1 U338 ( .A(n1855), .B(n1801), .C(n2774), .Y(n2259) );
  NAND2X1 U339 ( .A(\mem<23><2> ), .B(n1803), .Y(n2774) );
  OAI21X1 U340 ( .A(n1852), .B(n1801), .C(n2773), .Y(n2258) );
  NAND2X1 U341 ( .A(\mem<23><3> ), .B(n1803), .Y(n2773) );
  OAI21X1 U342 ( .A(n1849), .B(n1801), .C(n2772), .Y(n2257) );
  NAND2X1 U343 ( .A(\mem<23><4> ), .B(n1803), .Y(n2772) );
  OAI21X1 U344 ( .A(n1846), .B(n1801), .C(n2771), .Y(n2256) );
  NAND2X1 U345 ( .A(\mem<23><5> ), .B(n1803), .Y(n2771) );
  OAI21X1 U346 ( .A(n1843), .B(n1801), .C(n2770), .Y(n2255) );
  NAND2X1 U347 ( .A(\mem<23><6> ), .B(n1803), .Y(n2770) );
  OAI21X1 U348 ( .A(n1840), .B(n1801), .C(n2769), .Y(n2254) );
  NAND2X1 U349 ( .A(\mem<23><7> ), .B(n1803), .Y(n2769) );
  OAI21X1 U350 ( .A(n1839), .B(n1801), .C(n2768), .Y(n2253) );
  NAND2X1 U351 ( .A(\mem<23><8> ), .B(n1802), .Y(n2768) );
  OAI21X1 U352 ( .A(n1838), .B(n1801), .C(n2767), .Y(n2252) );
  NAND2X1 U353 ( .A(\mem<23><9> ), .B(n1802), .Y(n2767) );
  OAI21X1 U354 ( .A(n1837), .B(n1801), .C(n2766), .Y(n2251) );
  NAND2X1 U355 ( .A(\mem<23><10> ), .B(n1802), .Y(n2766) );
  OAI21X1 U356 ( .A(n1836), .B(n1801), .C(n2765), .Y(n2250) );
  NAND2X1 U357 ( .A(\mem<23><11> ), .B(n1802), .Y(n2765) );
  OAI21X1 U358 ( .A(n1835), .B(n1801), .C(n2764), .Y(n2249) );
  NAND2X1 U359 ( .A(\mem<23><12> ), .B(n1802), .Y(n2764) );
  OAI21X1 U360 ( .A(n1834), .B(n1801), .C(n2763), .Y(n2248) );
  NAND2X1 U361 ( .A(\mem<23><13> ), .B(n1802), .Y(n2763) );
  OAI21X1 U362 ( .A(n1833), .B(n1801), .C(n2762), .Y(n2247) );
  NAND2X1 U363 ( .A(\mem<23><14> ), .B(n1802), .Y(n2762) );
  OAI21X1 U364 ( .A(n1832), .B(n1801), .C(n2761), .Y(n2246) );
  NAND2X1 U365 ( .A(\mem<23><15> ), .B(n1802), .Y(n2761) );
  OAI21X1 U368 ( .A(n1861), .B(n1798), .C(n2760), .Y(n2245) );
  NAND2X1 U369 ( .A(\mem<22><0> ), .B(n1800), .Y(n2760) );
  OAI21X1 U370 ( .A(n1858), .B(n1798), .C(n2759), .Y(n2244) );
  NAND2X1 U371 ( .A(\mem<22><1> ), .B(n1800), .Y(n2759) );
  OAI21X1 U372 ( .A(n1855), .B(n1798), .C(n2758), .Y(n2243) );
  NAND2X1 U373 ( .A(\mem<22><2> ), .B(n1800), .Y(n2758) );
  OAI21X1 U374 ( .A(n1852), .B(n1798), .C(n2757), .Y(n2242) );
  NAND2X1 U375 ( .A(\mem<22><3> ), .B(n1800), .Y(n2757) );
  OAI21X1 U376 ( .A(n1849), .B(n1798), .C(n2756), .Y(n2241) );
  NAND2X1 U377 ( .A(\mem<22><4> ), .B(n1800), .Y(n2756) );
  OAI21X1 U378 ( .A(n1846), .B(n1798), .C(n2755), .Y(n2240) );
  NAND2X1 U379 ( .A(\mem<22><5> ), .B(n1800), .Y(n2755) );
  OAI21X1 U380 ( .A(n1843), .B(n1798), .C(n2754), .Y(n2239) );
  NAND2X1 U381 ( .A(\mem<22><6> ), .B(n1800), .Y(n2754) );
  OAI21X1 U382 ( .A(n1840), .B(n1798), .C(n2753), .Y(n2238) );
  NAND2X1 U383 ( .A(\mem<22><7> ), .B(n1800), .Y(n2753) );
  OAI21X1 U384 ( .A(n1839), .B(n1798), .C(n2752), .Y(n2237) );
  NAND2X1 U385 ( .A(\mem<22><8> ), .B(n1799), .Y(n2752) );
  OAI21X1 U386 ( .A(n1838), .B(n1798), .C(n2751), .Y(n2236) );
  NAND2X1 U387 ( .A(\mem<22><9> ), .B(n1799), .Y(n2751) );
  OAI21X1 U388 ( .A(n1837), .B(n1798), .C(n2750), .Y(n2235) );
  NAND2X1 U389 ( .A(\mem<22><10> ), .B(n1799), .Y(n2750) );
  OAI21X1 U390 ( .A(n1836), .B(n1798), .C(n2749), .Y(n2234) );
  NAND2X1 U391 ( .A(\mem<22><11> ), .B(n1799), .Y(n2749) );
  OAI21X1 U392 ( .A(n1835), .B(n1798), .C(n2748), .Y(n2233) );
  NAND2X1 U393 ( .A(\mem<22><12> ), .B(n1799), .Y(n2748) );
  OAI21X1 U394 ( .A(n1834), .B(n1798), .C(n2747), .Y(n2232) );
  NAND2X1 U395 ( .A(\mem<22><13> ), .B(n1799), .Y(n2747) );
  OAI21X1 U396 ( .A(n1833), .B(n1798), .C(n2746), .Y(n2231) );
  NAND2X1 U397 ( .A(\mem<22><14> ), .B(n1799), .Y(n2746) );
  OAI21X1 U398 ( .A(n1832), .B(n1798), .C(n2745), .Y(n2230) );
  NAND2X1 U399 ( .A(\mem<22><15> ), .B(n1799), .Y(n2745) );
  OAI21X1 U402 ( .A(n1861), .B(n1795), .C(n2744), .Y(n2229) );
  NAND2X1 U403 ( .A(\mem<21><0> ), .B(n1797), .Y(n2744) );
  OAI21X1 U404 ( .A(n1858), .B(n1795), .C(n2743), .Y(n2228) );
  NAND2X1 U405 ( .A(\mem<21><1> ), .B(n1797), .Y(n2743) );
  OAI21X1 U406 ( .A(n1855), .B(n1795), .C(n2742), .Y(n2227) );
  NAND2X1 U407 ( .A(\mem<21><2> ), .B(n1797), .Y(n2742) );
  OAI21X1 U408 ( .A(n1852), .B(n1795), .C(n2741), .Y(n2226) );
  NAND2X1 U409 ( .A(\mem<21><3> ), .B(n1797), .Y(n2741) );
  OAI21X1 U410 ( .A(n1849), .B(n1795), .C(n2740), .Y(n2225) );
  NAND2X1 U411 ( .A(\mem<21><4> ), .B(n1797), .Y(n2740) );
  OAI21X1 U412 ( .A(n1846), .B(n1795), .C(n2739), .Y(n2224) );
  NAND2X1 U413 ( .A(\mem<21><5> ), .B(n1797), .Y(n2739) );
  OAI21X1 U414 ( .A(n1843), .B(n1795), .C(n2738), .Y(n2223) );
  NAND2X1 U415 ( .A(\mem<21><6> ), .B(n1797), .Y(n2738) );
  OAI21X1 U416 ( .A(n1840), .B(n1795), .C(n2737), .Y(n2222) );
  NAND2X1 U417 ( .A(\mem<21><7> ), .B(n1797), .Y(n2737) );
  OAI21X1 U418 ( .A(n1839), .B(n1795), .C(n2736), .Y(n2221) );
  NAND2X1 U419 ( .A(\mem<21><8> ), .B(n1796), .Y(n2736) );
  OAI21X1 U420 ( .A(n1838), .B(n1795), .C(n2735), .Y(n2220) );
  NAND2X1 U421 ( .A(\mem<21><9> ), .B(n1796), .Y(n2735) );
  OAI21X1 U422 ( .A(n1837), .B(n1795), .C(n2734), .Y(n2219) );
  NAND2X1 U423 ( .A(\mem<21><10> ), .B(n1796), .Y(n2734) );
  OAI21X1 U424 ( .A(n1836), .B(n1795), .C(n2733), .Y(n2218) );
  NAND2X1 U425 ( .A(\mem<21><11> ), .B(n1796), .Y(n2733) );
  OAI21X1 U426 ( .A(n1835), .B(n1795), .C(n2732), .Y(n2217) );
  NAND2X1 U427 ( .A(\mem<21><12> ), .B(n1796), .Y(n2732) );
  OAI21X1 U428 ( .A(n1834), .B(n1795), .C(n2731), .Y(n2216) );
  NAND2X1 U429 ( .A(\mem<21><13> ), .B(n1796), .Y(n2731) );
  OAI21X1 U430 ( .A(n1833), .B(n1795), .C(n2730), .Y(n2215) );
  NAND2X1 U431 ( .A(\mem<21><14> ), .B(n1796), .Y(n2730) );
  OAI21X1 U432 ( .A(n1832), .B(n1795), .C(n2729), .Y(n2214) );
  NAND2X1 U433 ( .A(\mem<21><15> ), .B(n1796), .Y(n2729) );
  OAI21X1 U436 ( .A(n1861), .B(n1792), .C(n2728), .Y(n2213) );
  NAND2X1 U437 ( .A(\mem<20><0> ), .B(n1794), .Y(n2728) );
  OAI21X1 U438 ( .A(n1858), .B(n1792), .C(n2727), .Y(n2212) );
  NAND2X1 U439 ( .A(\mem<20><1> ), .B(n1794), .Y(n2727) );
  OAI21X1 U440 ( .A(n1855), .B(n1792), .C(n2726), .Y(n2211) );
  NAND2X1 U441 ( .A(\mem<20><2> ), .B(n1794), .Y(n2726) );
  OAI21X1 U442 ( .A(n1852), .B(n1792), .C(n2725), .Y(n2210) );
  NAND2X1 U443 ( .A(\mem<20><3> ), .B(n1794), .Y(n2725) );
  OAI21X1 U444 ( .A(n1849), .B(n1792), .C(n2724), .Y(n2209) );
  NAND2X1 U445 ( .A(\mem<20><4> ), .B(n1794), .Y(n2724) );
  OAI21X1 U446 ( .A(n1846), .B(n1792), .C(n2723), .Y(n2208) );
  NAND2X1 U447 ( .A(\mem<20><5> ), .B(n1794), .Y(n2723) );
  OAI21X1 U448 ( .A(n1843), .B(n1792), .C(n2722), .Y(n2207) );
  NAND2X1 U449 ( .A(\mem<20><6> ), .B(n1794), .Y(n2722) );
  OAI21X1 U450 ( .A(n1840), .B(n1792), .C(n2721), .Y(n2206) );
  NAND2X1 U451 ( .A(\mem<20><7> ), .B(n1794), .Y(n2721) );
  OAI21X1 U452 ( .A(n1839), .B(n1792), .C(n2720), .Y(n2205) );
  NAND2X1 U453 ( .A(\mem<20><8> ), .B(n1793), .Y(n2720) );
  OAI21X1 U454 ( .A(n1838), .B(n1792), .C(n2719), .Y(n2204) );
  NAND2X1 U455 ( .A(\mem<20><9> ), .B(n1793), .Y(n2719) );
  OAI21X1 U456 ( .A(n1837), .B(n1792), .C(n2718), .Y(n2203) );
  NAND2X1 U457 ( .A(\mem<20><10> ), .B(n1793), .Y(n2718) );
  OAI21X1 U458 ( .A(n1836), .B(n1792), .C(n2717), .Y(n2202) );
  NAND2X1 U459 ( .A(\mem<20><11> ), .B(n1793), .Y(n2717) );
  OAI21X1 U460 ( .A(n1835), .B(n1792), .C(n2716), .Y(n2201) );
  NAND2X1 U461 ( .A(\mem<20><12> ), .B(n1793), .Y(n2716) );
  OAI21X1 U462 ( .A(n1834), .B(n1792), .C(n2715), .Y(n2200) );
  NAND2X1 U463 ( .A(\mem<20><13> ), .B(n1793), .Y(n2715) );
  OAI21X1 U464 ( .A(n1833), .B(n1792), .C(n2714), .Y(n2199) );
  NAND2X1 U465 ( .A(\mem<20><14> ), .B(n1793), .Y(n2714) );
  OAI21X1 U466 ( .A(n1832), .B(n1792), .C(n2713), .Y(n2198) );
  NAND2X1 U467 ( .A(\mem<20><15> ), .B(n1793), .Y(n2713) );
  OAI21X1 U470 ( .A(n1861), .B(n1789), .C(n2712), .Y(n2197) );
  NAND2X1 U471 ( .A(\mem<19><0> ), .B(n1791), .Y(n2712) );
  OAI21X1 U472 ( .A(n1858), .B(n1789), .C(n2711), .Y(n2196) );
  NAND2X1 U473 ( .A(\mem<19><1> ), .B(n1791), .Y(n2711) );
  OAI21X1 U474 ( .A(n1855), .B(n1789), .C(n2710), .Y(n2195) );
  NAND2X1 U475 ( .A(\mem<19><2> ), .B(n1791), .Y(n2710) );
  OAI21X1 U476 ( .A(n1852), .B(n1789), .C(n2709), .Y(n2194) );
  NAND2X1 U477 ( .A(\mem<19><3> ), .B(n1791), .Y(n2709) );
  OAI21X1 U478 ( .A(n1849), .B(n1789), .C(n2708), .Y(n2193) );
  NAND2X1 U479 ( .A(\mem<19><4> ), .B(n1791), .Y(n2708) );
  OAI21X1 U480 ( .A(n1846), .B(n1789), .C(n2707), .Y(n2192) );
  NAND2X1 U481 ( .A(\mem<19><5> ), .B(n1791), .Y(n2707) );
  OAI21X1 U482 ( .A(n1843), .B(n1789), .C(n2706), .Y(n2191) );
  NAND2X1 U483 ( .A(\mem<19><6> ), .B(n1791), .Y(n2706) );
  OAI21X1 U484 ( .A(n1840), .B(n1789), .C(n2705), .Y(n2190) );
  NAND2X1 U485 ( .A(\mem<19><7> ), .B(n1791), .Y(n2705) );
  OAI21X1 U486 ( .A(n1839), .B(n1789), .C(n2704), .Y(n2189) );
  NAND2X1 U487 ( .A(\mem<19><8> ), .B(n1790), .Y(n2704) );
  OAI21X1 U488 ( .A(n1838), .B(n1789), .C(n2703), .Y(n2188) );
  NAND2X1 U489 ( .A(\mem<19><9> ), .B(n1790), .Y(n2703) );
  OAI21X1 U490 ( .A(n1837), .B(n1789), .C(n2702), .Y(n2187) );
  NAND2X1 U491 ( .A(\mem<19><10> ), .B(n1790), .Y(n2702) );
  OAI21X1 U492 ( .A(n1836), .B(n1789), .C(n2701), .Y(n2186) );
  NAND2X1 U493 ( .A(\mem<19><11> ), .B(n1790), .Y(n2701) );
  OAI21X1 U494 ( .A(n1835), .B(n1789), .C(n2700), .Y(n2185) );
  NAND2X1 U495 ( .A(\mem<19><12> ), .B(n1790), .Y(n2700) );
  OAI21X1 U496 ( .A(n1834), .B(n1789), .C(n2699), .Y(n2184) );
  NAND2X1 U497 ( .A(\mem<19><13> ), .B(n1790), .Y(n2699) );
  OAI21X1 U498 ( .A(n1833), .B(n1789), .C(n2698), .Y(n2183) );
  NAND2X1 U499 ( .A(\mem<19><14> ), .B(n1790), .Y(n2698) );
  OAI21X1 U500 ( .A(n1832), .B(n1789), .C(n2697), .Y(n2182) );
  NAND2X1 U501 ( .A(\mem<19><15> ), .B(n1790), .Y(n2697) );
  OAI21X1 U504 ( .A(n1862), .B(n1786), .C(n2696), .Y(n2181) );
  NAND2X1 U505 ( .A(\mem<18><0> ), .B(n1788), .Y(n2696) );
  OAI21X1 U506 ( .A(n1859), .B(n1786), .C(n2695), .Y(n2180) );
  NAND2X1 U507 ( .A(\mem<18><1> ), .B(n1788), .Y(n2695) );
  OAI21X1 U508 ( .A(n1856), .B(n1786), .C(n2694), .Y(n2179) );
  NAND2X1 U509 ( .A(\mem<18><2> ), .B(n1788), .Y(n2694) );
  OAI21X1 U510 ( .A(n1853), .B(n1786), .C(n2693), .Y(n2178) );
  NAND2X1 U511 ( .A(\mem<18><3> ), .B(n1788), .Y(n2693) );
  OAI21X1 U512 ( .A(n1850), .B(n1786), .C(n2692), .Y(n2177) );
  NAND2X1 U513 ( .A(\mem<18><4> ), .B(n1788), .Y(n2692) );
  OAI21X1 U514 ( .A(n1847), .B(n1786), .C(n2691), .Y(n2176) );
  NAND2X1 U515 ( .A(\mem<18><5> ), .B(n1788), .Y(n2691) );
  OAI21X1 U516 ( .A(n1844), .B(n1786), .C(n2690), .Y(n2175) );
  NAND2X1 U517 ( .A(\mem<18><6> ), .B(n1788), .Y(n2690) );
  OAI21X1 U518 ( .A(n1841), .B(n1786), .C(n2689), .Y(n2174) );
  NAND2X1 U519 ( .A(\mem<18><7> ), .B(n1788), .Y(n2689) );
  OAI21X1 U520 ( .A(n1839), .B(n1786), .C(n2688), .Y(n2173) );
  NAND2X1 U521 ( .A(\mem<18><8> ), .B(n1787), .Y(n2688) );
  OAI21X1 U522 ( .A(n1838), .B(n1786), .C(n2687), .Y(n2172) );
  NAND2X1 U523 ( .A(\mem<18><9> ), .B(n1787), .Y(n2687) );
  OAI21X1 U524 ( .A(n1837), .B(n1786), .C(n2686), .Y(n2171) );
  NAND2X1 U525 ( .A(\mem<18><10> ), .B(n1787), .Y(n2686) );
  OAI21X1 U526 ( .A(n1836), .B(n1786), .C(n2685), .Y(n2170) );
  NAND2X1 U527 ( .A(\mem<18><11> ), .B(n1787), .Y(n2685) );
  OAI21X1 U528 ( .A(n1835), .B(n1786), .C(n2684), .Y(n2169) );
  NAND2X1 U529 ( .A(\mem<18><12> ), .B(n1787), .Y(n2684) );
  OAI21X1 U530 ( .A(n1834), .B(n1786), .C(n2683), .Y(n2168) );
  NAND2X1 U531 ( .A(\mem<18><13> ), .B(n1787), .Y(n2683) );
  OAI21X1 U532 ( .A(n1833), .B(n1786), .C(n2682), .Y(n2167) );
  NAND2X1 U533 ( .A(\mem<18><14> ), .B(n1787), .Y(n2682) );
  OAI21X1 U534 ( .A(n1832), .B(n1786), .C(n2681), .Y(n2166) );
  NAND2X1 U535 ( .A(\mem<18><15> ), .B(n1787), .Y(n2681) );
  OAI21X1 U538 ( .A(n1862), .B(n1783), .C(n2680), .Y(n2165) );
  NAND2X1 U539 ( .A(\mem<17><0> ), .B(n1785), .Y(n2680) );
  OAI21X1 U540 ( .A(n1859), .B(n1783), .C(n2679), .Y(n2164) );
  NAND2X1 U541 ( .A(\mem<17><1> ), .B(n1785), .Y(n2679) );
  OAI21X1 U542 ( .A(n1856), .B(n1783), .C(n2678), .Y(n2163) );
  NAND2X1 U543 ( .A(\mem<17><2> ), .B(n1785), .Y(n2678) );
  OAI21X1 U544 ( .A(n1853), .B(n1783), .C(n2677), .Y(n2162) );
  NAND2X1 U545 ( .A(\mem<17><3> ), .B(n1785), .Y(n2677) );
  OAI21X1 U546 ( .A(n1850), .B(n1783), .C(n2676), .Y(n2161) );
  NAND2X1 U547 ( .A(\mem<17><4> ), .B(n1785), .Y(n2676) );
  OAI21X1 U548 ( .A(n1847), .B(n1783), .C(n2675), .Y(n2160) );
  NAND2X1 U549 ( .A(\mem<17><5> ), .B(n1785), .Y(n2675) );
  OAI21X1 U550 ( .A(n1844), .B(n1783), .C(n2674), .Y(n2159) );
  NAND2X1 U551 ( .A(\mem<17><6> ), .B(n1785), .Y(n2674) );
  OAI21X1 U552 ( .A(n1841), .B(n1783), .C(n2673), .Y(n2158) );
  NAND2X1 U553 ( .A(\mem<17><7> ), .B(n1785), .Y(n2673) );
  OAI21X1 U554 ( .A(n1839), .B(n1783), .C(n2672), .Y(n2157) );
  NAND2X1 U555 ( .A(\mem<17><8> ), .B(n1784), .Y(n2672) );
  OAI21X1 U556 ( .A(n1838), .B(n1783), .C(n2671), .Y(n2156) );
  NAND2X1 U557 ( .A(\mem<17><9> ), .B(n1784), .Y(n2671) );
  OAI21X1 U558 ( .A(n1837), .B(n1783), .C(n2670), .Y(n2155) );
  NAND2X1 U559 ( .A(\mem<17><10> ), .B(n1784), .Y(n2670) );
  OAI21X1 U560 ( .A(n1836), .B(n1783), .C(n2669), .Y(n2154) );
  NAND2X1 U561 ( .A(\mem<17><11> ), .B(n1784), .Y(n2669) );
  OAI21X1 U562 ( .A(n1835), .B(n1783), .C(n2668), .Y(n2153) );
  NAND2X1 U563 ( .A(\mem<17><12> ), .B(n1784), .Y(n2668) );
  OAI21X1 U564 ( .A(n1834), .B(n1783), .C(n2667), .Y(n2152) );
  NAND2X1 U565 ( .A(\mem<17><13> ), .B(n1784), .Y(n2667) );
  OAI21X1 U566 ( .A(n1833), .B(n1783), .C(n2666), .Y(n2151) );
  NAND2X1 U567 ( .A(\mem<17><14> ), .B(n1784), .Y(n2666) );
  OAI21X1 U568 ( .A(n1832), .B(n1783), .C(n2665), .Y(n2150) );
  NAND2X1 U569 ( .A(\mem<17><15> ), .B(n1784), .Y(n2665) );
  OAI21X1 U572 ( .A(n1862), .B(n1780), .C(n2664), .Y(n2149) );
  NAND2X1 U573 ( .A(\mem<16><0> ), .B(n1782), .Y(n2664) );
  OAI21X1 U574 ( .A(n1859), .B(n1780), .C(n2663), .Y(n2148) );
  NAND2X1 U575 ( .A(\mem<16><1> ), .B(n1782), .Y(n2663) );
  OAI21X1 U576 ( .A(n1856), .B(n1780), .C(n2662), .Y(n2147) );
  NAND2X1 U577 ( .A(\mem<16><2> ), .B(n1782), .Y(n2662) );
  OAI21X1 U578 ( .A(n1853), .B(n1780), .C(n2661), .Y(n2146) );
  NAND2X1 U579 ( .A(\mem<16><3> ), .B(n1782), .Y(n2661) );
  OAI21X1 U580 ( .A(n1850), .B(n1780), .C(n2660), .Y(n2145) );
  NAND2X1 U581 ( .A(\mem<16><4> ), .B(n1782), .Y(n2660) );
  OAI21X1 U582 ( .A(n1847), .B(n1780), .C(n2659), .Y(n2144) );
  NAND2X1 U583 ( .A(\mem<16><5> ), .B(n1782), .Y(n2659) );
  OAI21X1 U584 ( .A(n1844), .B(n1780), .C(n2658), .Y(n2143) );
  NAND2X1 U585 ( .A(\mem<16><6> ), .B(n1782), .Y(n2658) );
  OAI21X1 U586 ( .A(n1841), .B(n1780), .C(n2657), .Y(n2142) );
  NAND2X1 U587 ( .A(\mem<16><7> ), .B(n1782), .Y(n2657) );
  OAI21X1 U588 ( .A(n1839), .B(n1780), .C(n2656), .Y(n2141) );
  NAND2X1 U589 ( .A(\mem<16><8> ), .B(n1781), .Y(n2656) );
  OAI21X1 U590 ( .A(n1838), .B(n1780), .C(n2655), .Y(n2140) );
  NAND2X1 U591 ( .A(\mem<16><9> ), .B(n1781), .Y(n2655) );
  OAI21X1 U592 ( .A(n1837), .B(n1780), .C(n2654), .Y(n2139) );
  NAND2X1 U593 ( .A(\mem<16><10> ), .B(n1781), .Y(n2654) );
  OAI21X1 U594 ( .A(n1836), .B(n1780), .C(n2653), .Y(n2138) );
  NAND2X1 U595 ( .A(\mem<16><11> ), .B(n1781), .Y(n2653) );
  OAI21X1 U596 ( .A(n1835), .B(n1780), .C(n2652), .Y(n2137) );
  NAND2X1 U597 ( .A(\mem<16><12> ), .B(n1781), .Y(n2652) );
  OAI21X1 U598 ( .A(n1834), .B(n1780), .C(n2651), .Y(n2136) );
  NAND2X1 U599 ( .A(\mem<16><13> ), .B(n1781), .Y(n2651) );
  OAI21X1 U600 ( .A(n1833), .B(n1780), .C(n2650), .Y(n2135) );
  NAND2X1 U601 ( .A(\mem<16><14> ), .B(n1781), .Y(n2650) );
  OAI21X1 U602 ( .A(n1832), .B(n1780), .C(n2649), .Y(n2134) );
  NAND2X1 U603 ( .A(\mem<16><15> ), .B(n1781), .Y(n2649) );
  NAND3X1 U606 ( .A(n2777), .B(n1871), .C(N14), .Y(n2648) );
  OAI21X1 U607 ( .A(n1862), .B(n1777), .C(n2647), .Y(n2133) );
  NAND2X1 U608 ( .A(\mem<15><0> ), .B(n1779), .Y(n2647) );
  OAI21X1 U609 ( .A(n1859), .B(n1777), .C(n2646), .Y(n2132) );
  NAND2X1 U610 ( .A(\mem<15><1> ), .B(n1779), .Y(n2646) );
  OAI21X1 U611 ( .A(n1856), .B(n1777), .C(n2645), .Y(n2131) );
  NAND2X1 U612 ( .A(\mem<15><2> ), .B(n1779), .Y(n2645) );
  OAI21X1 U613 ( .A(n1853), .B(n1777), .C(n2644), .Y(n2130) );
  NAND2X1 U614 ( .A(\mem<15><3> ), .B(n1779), .Y(n2644) );
  OAI21X1 U615 ( .A(n1850), .B(n1777), .C(n2643), .Y(n2129) );
  NAND2X1 U616 ( .A(\mem<15><4> ), .B(n1779), .Y(n2643) );
  OAI21X1 U617 ( .A(n1847), .B(n1777), .C(n2642), .Y(n2128) );
  NAND2X1 U618 ( .A(\mem<15><5> ), .B(n1779), .Y(n2642) );
  OAI21X1 U619 ( .A(n1844), .B(n1777), .C(n2641), .Y(n2127) );
  NAND2X1 U620 ( .A(\mem<15><6> ), .B(n1779), .Y(n2641) );
  OAI21X1 U621 ( .A(n1841), .B(n1777), .C(n2640), .Y(n2126) );
  NAND2X1 U622 ( .A(\mem<15><7> ), .B(n1779), .Y(n2640) );
  OAI21X1 U623 ( .A(n1839), .B(n1777), .C(n2639), .Y(n2125) );
  NAND2X1 U624 ( .A(\mem<15><8> ), .B(n1778), .Y(n2639) );
  OAI21X1 U625 ( .A(n1838), .B(n1777), .C(n2638), .Y(n2124) );
  NAND2X1 U626 ( .A(\mem<15><9> ), .B(n1778), .Y(n2638) );
  OAI21X1 U627 ( .A(n1837), .B(n1777), .C(n2637), .Y(n2123) );
  NAND2X1 U628 ( .A(\mem<15><10> ), .B(n1778), .Y(n2637) );
  OAI21X1 U629 ( .A(n1836), .B(n1777), .C(n2636), .Y(n2122) );
  NAND2X1 U630 ( .A(\mem<15><11> ), .B(n1778), .Y(n2636) );
  OAI21X1 U631 ( .A(n1835), .B(n1777), .C(n2635), .Y(n2121) );
  NAND2X1 U632 ( .A(\mem<15><12> ), .B(n1778), .Y(n2635) );
  OAI21X1 U633 ( .A(n1834), .B(n1777), .C(n2634), .Y(n2120) );
  NAND2X1 U634 ( .A(\mem<15><13> ), .B(n1778), .Y(n2634) );
  OAI21X1 U635 ( .A(n1833), .B(n1777), .C(n2633), .Y(n2119) );
  NAND2X1 U636 ( .A(\mem<15><14> ), .B(n1778), .Y(n2633) );
  OAI21X1 U637 ( .A(n1832), .B(n1777), .C(n2632), .Y(n2118) );
  NAND2X1 U638 ( .A(\mem<15><15> ), .B(n1778), .Y(n2632) );
  OAI21X1 U641 ( .A(n1862), .B(n1774), .C(n2631), .Y(n2117) );
  NAND2X1 U642 ( .A(\mem<14><0> ), .B(n1776), .Y(n2631) );
  OAI21X1 U643 ( .A(n1859), .B(n1774), .C(n2630), .Y(n2116) );
  NAND2X1 U644 ( .A(\mem<14><1> ), .B(n1776), .Y(n2630) );
  OAI21X1 U645 ( .A(n1856), .B(n1774), .C(n2629), .Y(n2115) );
  NAND2X1 U646 ( .A(\mem<14><2> ), .B(n1776), .Y(n2629) );
  OAI21X1 U647 ( .A(n1853), .B(n1774), .C(n2628), .Y(n2114) );
  NAND2X1 U648 ( .A(\mem<14><3> ), .B(n1776), .Y(n2628) );
  OAI21X1 U649 ( .A(n1850), .B(n1774), .C(n2627), .Y(n2113) );
  NAND2X1 U650 ( .A(\mem<14><4> ), .B(n1776), .Y(n2627) );
  OAI21X1 U651 ( .A(n1847), .B(n1774), .C(n2626), .Y(n2112) );
  NAND2X1 U652 ( .A(\mem<14><5> ), .B(n1776), .Y(n2626) );
  OAI21X1 U653 ( .A(n1844), .B(n1774), .C(n2625), .Y(n2111) );
  NAND2X1 U654 ( .A(\mem<14><6> ), .B(n1776), .Y(n2625) );
  OAI21X1 U655 ( .A(n1841), .B(n1774), .C(n2624), .Y(n2110) );
  NAND2X1 U656 ( .A(\mem<14><7> ), .B(n1776), .Y(n2624) );
  OAI21X1 U657 ( .A(n1839), .B(n1774), .C(n2623), .Y(n2109) );
  NAND2X1 U658 ( .A(\mem<14><8> ), .B(n1775), .Y(n2623) );
  OAI21X1 U659 ( .A(n1838), .B(n1774), .C(n2622), .Y(n2108) );
  NAND2X1 U660 ( .A(\mem<14><9> ), .B(n1775), .Y(n2622) );
  OAI21X1 U661 ( .A(n1837), .B(n1774), .C(n2621), .Y(n2107) );
  NAND2X1 U662 ( .A(\mem<14><10> ), .B(n1775), .Y(n2621) );
  OAI21X1 U663 ( .A(n1836), .B(n1774), .C(n2620), .Y(n2106) );
  NAND2X1 U664 ( .A(\mem<14><11> ), .B(n1775), .Y(n2620) );
  OAI21X1 U665 ( .A(n1835), .B(n1774), .C(n2619), .Y(n2105) );
  NAND2X1 U666 ( .A(\mem<14><12> ), .B(n1775), .Y(n2619) );
  OAI21X1 U667 ( .A(n1834), .B(n1774), .C(n2618), .Y(n2104) );
  NAND2X1 U668 ( .A(\mem<14><13> ), .B(n1775), .Y(n2618) );
  OAI21X1 U669 ( .A(n1833), .B(n1774), .C(n2617), .Y(n2103) );
  NAND2X1 U670 ( .A(\mem<14><14> ), .B(n1775), .Y(n2617) );
  OAI21X1 U671 ( .A(n1832), .B(n1774), .C(n2616), .Y(n2102) );
  NAND2X1 U672 ( .A(\mem<14><15> ), .B(n1775), .Y(n2616) );
  OAI21X1 U675 ( .A(n1862), .B(n1771), .C(n2615), .Y(n2101) );
  NAND2X1 U676 ( .A(\mem<13><0> ), .B(n1773), .Y(n2615) );
  OAI21X1 U677 ( .A(n1859), .B(n1771), .C(n2614), .Y(n2100) );
  NAND2X1 U678 ( .A(\mem<13><1> ), .B(n1773), .Y(n2614) );
  OAI21X1 U679 ( .A(n1856), .B(n1771), .C(n2613), .Y(n2099) );
  NAND2X1 U680 ( .A(\mem<13><2> ), .B(n1773), .Y(n2613) );
  OAI21X1 U681 ( .A(n1853), .B(n1771), .C(n2612), .Y(n2098) );
  NAND2X1 U682 ( .A(\mem<13><3> ), .B(n1773), .Y(n2612) );
  OAI21X1 U683 ( .A(n1850), .B(n1771), .C(n2611), .Y(n2097) );
  NAND2X1 U684 ( .A(\mem<13><4> ), .B(n1773), .Y(n2611) );
  OAI21X1 U685 ( .A(n1847), .B(n1771), .C(n2610), .Y(n2096) );
  NAND2X1 U686 ( .A(\mem<13><5> ), .B(n1773), .Y(n2610) );
  OAI21X1 U687 ( .A(n1844), .B(n1771), .C(n2609), .Y(n2095) );
  NAND2X1 U688 ( .A(\mem<13><6> ), .B(n1773), .Y(n2609) );
  OAI21X1 U689 ( .A(n1841), .B(n1771), .C(n2608), .Y(n2094) );
  NAND2X1 U690 ( .A(\mem<13><7> ), .B(n1773), .Y(n2608) );
  OAI21X1 U691 ( .A(n1839), .B(n1771), .C(n2607), .Y(n2093) );
  NAND2X1 U692 ( .A(\mem<13><8> ), .B(n1772), .Y(n2607) );
  OAI21X1 U693 ( .A(n1838), .B(n1771), .C(n2606), .Y(n2092) );
  NAND2X1 U694 ( .A(\mem<13><9> ), .B(n1772), .Y(n2606) );
  OAI21X1 U695 ( .A(n1837), .B(n1771), .C(n2605), .Y(n2091) );
  NAND2X1 U696 ( .A(\mem<13><10> ), .B(n1772), .Y(n2605) );
  OAI21X1 U697 ( .A(n1836), .B(n1771), .C(n2604), .Y(n2090) );
  NAND2X1 U698 ( .A(\mem<13><11> ), .B(n1772), .Y(n2604) );
  OAI21X1 U699 ( .A(n1835), .B(n1771), .C(n2603), .Y(n2089) );
  NAND2X1 U700 ( .A(\mem<13><12> ), .B(n1772), .Y(n2603) );
  OAI21X1 U701 ( .A(n1834), .B(n1771), .C(n2602), .Y(n2088) );
  NAND2X1 U702 ( .A(\mem<13><13> ), .B(n1772), .Y(n2602) );
  OAI21X1 U703 ( .A(n1833), .B(n1771), .C(n2601), .Y(n2087) );
  NAND2X1 U704 ( .A(\mem<13><14> ), .B(n1772), .Y(n2601) );
  OAI21X1 U705 ( .A(n1832), .B(n1771), .C(n2600), .Y(n2086) );
  NAND2X1 U706 ( .A(\mem<13><15> ), .B(n1772), .Y(n2600) );
  OAI21X1 U709 ( .A(n1862), .B(n1768), .C(n2599), .Y(n2085) );
  NAND2X1 U710 ( .A(\mem<12><0> ), .B(n1770), .Y(n2599) );
  OAI21X1 U711 ( .A(n1859), .B(n1768), .C(n2598), .Y(n2084) );
  NAND2X1 U712 ( .A(\mem<12><1> ), .B(n1770), .Y(n2598) );
  OAI21X1 U713 ( .A(n1856), .B(n1768), .C(n2597), .Y(n2083) );
  NAND2X1 U714 ( .A(\mem<12><2> ), .B(n1770), .Y(n2597) );
  OAI21X1 U715 ( .A(n1853), .B(n1768), .C(n2596), .Y(n2082) );
  NAND2X1 U716 ( .A(\mem<12><3> ), .B(n1770), .Y(n2596) );
  OAI21X1 U717 ( .A(n1850), .B(n1768), .C(n2595), .Y(n2081) );
  NAND2X1 U718 ( .A(\mem<12><4> ), .B(n1770), .Y(n2595) );
  OAI21X1 U719 ( .A(n1847), .B(n1768), .C(n2594), .Y(n2080) );
  NAND2X1 U720 ( .A(\mem<12><5> ), .B(n1770), .Y(n2594) );
  OAI21X1 U721 ( .A(n1844), .B(n1768), .C(n2593), .Y(n2079) );
  NAND2X1 U722 ( .A(\mem<12><6> ), .B(n1770), .Y(n2593) );
  OAI21X1 U723 ( .A(n1841), .B(n1768), .C(n2592), .Y(n2078) );
  NAND2X1 U724 ( .A(\mem<12><7> ), .B(n1770), .Y(n2592) );
  OAI21X1 U725 ( .A(n1839), .B(n1768), .C(n2591), .Y(n2077) );
  NAND2X1 U726 ( .A(\mem<12><8> ), .B(n1769), .Y(n2591) );
  OAI21X1 U727 ( .A(n1838), .B(n1768), .C(n2590), .Y(n2076) );
  NAND2X1 U728 ( .A(\mem<12><9> ), .B(n1769), .Y(n2590) );
  OAI21X1 U729 ( .A(n1837), .B(n1768), .C(n2589), .Y(n2075) );
  NAND2X1 U730 ( .A(\mem<12><10> ), .B(n1769), .Y(n2589) );
  OAI21X1 U731 ( .A(n1836), .B(n1768), .C(n2588), .Y(n2074) );
  NAND2X1 U732 ( .A(\mem<12><11> ), .B(n1769), .Y(n2588) );
  OAI21X1 U733 ( .A(n1835), .B(n1768), .C(n2587), .Y(n2073) );
  NAND2X1 U734 ( .A(\mem<12><12> ), .B(n1769), .Y(n2587) );
  OAI21X1 U735 ( .A(n1834), .B(n1768), .C(n2586), .Y(n2072) );
  NAND2X1 U736 ( .A(\mem<12><13> ), .B(n1769), .Y(n2586) );
  OAI21X1 U737 ( .A(n1833), .B(n1768), .C(n2585), .Y(n2071) );
  NAND2X1 U738 ( .A(\mem<12><14> ), .B(n1769), .Y(n2585) );
  OAI21X1 U739 ( .A(n1832), .B(n1768), .C(n2584), .Y(n2070) );
  NAND2X1 U740 ( .A(\mem<12><15> ), .B(n1769), .Y(n2584) );
  OAI21X1 U743 ( .A(n1862), .B(n1765), .C(n2583), .Y(n2069) );
  NAND2X1 U744 ( .A(\mem<11><0> ), .B(n1767), .Y(n2583) );
  OAI21X1 U745 ( .A(n1859), .B(n1765), .C(n2582), .Y(n2068) );
  NAND2X1 U746 ( .A(\mem<11><1> ), .B(n1767), .Y(n2582) );
  OAI21X1 U747 ( .A(n1856), .B(n1765), .C(n2581), .Y(n2067) );
  NAND2X1 U748 ( .A(\mem<11><2> ), .B(n1767), .Y(n2581) );
  OAI21X1 U749 ( .A(n1853), .B(n1765), .C(n2580), .Y(n2066) );
  NAND2X1 U750 ( .A(\mem<11><3> ), .B(n1767), .Y(n2580) );
  OAI21X1 U751 ( .A(n1850), .B(n1765), .C(n2579), .Y(n2065) );
  NAND2X1 U752 ( .A(\mem<11><4> ), .B(n1767), .Y(n2579) );
  OAI21X1 U753 ( .A(n1847), .B(n1765), .C(n2578), .Y(n2064) );
  NAND2X1 U754 ( .A(\mem<11><5> ), .B(n1767), .Y(n2578) );
  OAI21X1 U755 ( .A(n1844), .B(n1765), .C(n2577), .Y(n2063) );
  NAND2X1 U756 ( .A(\mem<11><6> ), .B(n1767), .Y(n2577) );
  OAI21X1 U757 ( .A(n1841), .B(n1765), .C(n2576), .Y(n2062) );
  NAND2X1 U758 ( .A(\mem<11><7> ), .B(n1767), .Y(n2576) );
  OAI21X1 U759 ( .A(n1839), .B(n1765), .C(n2575), .Y(n2061) );
  NAND2X1 U760 ( .A(\mem<11><8> ), .B(n1766), .Y(n2575) );
  OAI21X1 U761 ( .A(n1838), .B(n1765), .C(n2574), .Y(n2060) );
  NAND2X1 U762 ( .A(\mem<11><9> ), .B(n1766), .Y(n2574) );
  OAI21X1 U763 ( .A(n1837), .B(n1765), .C(n2573), .Y(n2059) );
  NAND2X1 U764 ( .A(\mem<11><10> ), .B(n1766), .Y(n2573) );
  OAI21X1 U765 ( .A(n1836), .B(n1765), .C(n2572), .Y(n2058) );
  NAND2X1 U766 ( .A(\mem<11><11> ), .B(n1766), .Y(n2572) );
  OAI21X1 U767 ( .A(n1835), .B(n1765), .C(n2571), .Y(n2057) );
  NAND2X1 U768 ( .A(\mem<11><12> ), .B(n1766), .Y(n2571) );
  OAI21X1 U769 ( .A(n1834), .B(n1765), .C(n2570), .Y(n2056) );
  NAND2X1 U770 ( .A(\mem<11><13> ), .B(n1766), .Y(n2570) );
  OAI21X1 U771 ( .A(n1833), .B(n1765), .C(n2569), .Y(n2055) );
  NAND2X1 U772 ( .A(\mem<11><14> ), .B(n1766), .Y(n2569) );
  OAI21X1 U773 ( .A(n1832), .B(n1765), .C(n2568), .Y(n2054) );
  NAND2X1 U774 ( .A(\mem<11><15> ), .B(n1766), .Y(n2568) );
  OAI21X1 U777 ( .A(n1862), .B(n1762), .C(n2567), .Y(n2053) );
  NAND2X1 U778 ( .A(\mem<10><0> ), .B(n1764), .Y(n2567) );
  OAI21X1 U779 ( .A(n1859), .B(n1762), .C(n2566), .Y(n2052) );
  NAND2X1 U780 ( .A(\mem<10><1> ), .B(n1764), .Y(n2566) );
  OAI21X1 U781 ( .A(n1856), .B(n1762), .C(n2565), .Y(n2051) );
  NAND2X1 U782 ( .A(\mem<10><2> ), .B(n1764), .Y(n2565) );
  OAI21X1 U783 ( .A(n1853), .B(n1762), .C(n2564), .Y(n2050) );
  NAND2X1 U784 ( .A(\mem<10><3> ), .B(n1764), .Y(n2564) );
  OAI21X1 U785 ( .A(n1850), .B(n1762), .C(n2563), .Y(n2049) );
  NAND2X1 U786 ( .A(\mem<10><4> ), .B(n1764), .Y(n2563) );
  OAI21X1 U787 ( .A(n1847), .B(n1762), .C(n2562), .Y(n2048) );
  NAND2X1 U788 ( .A(\mem<10><5> ), .B(n1764), .Y(n2562) );
  OAI21X1 U789 ( .A(n1844), .B(n1762), .C(n2561), .Y(n2047) );
  NAND2X1 U790 ( .A(\mem<10><6> ), .B(n1764), .Y(n2561) );
  OAI21X1 U791 ( .A(n1841), .B(n1762), .C(n2560), .Y(n2046) );
  NAND2X1 U792 ( .A(\mem<10><7> ), .B(n1764), .Y(n2560) );
  OAI21X1 U793 ( .A(n1839), .B(n1762), .C(n2559), .Y(n2045) );
  NAND2X1 U794 ( .A(\mem<10><8> ), .B(n1763), .Y(n2559) );
  OAI21X1 U795 ( .A(n1838), .B(n1762), .C(n2558), .Y(n2044) );
  NAND2X1 U796 ( .A(\mem<10><9> ), .B(n1763), .Y(n2558) );
  OAI21X1 U797 ( .A(n1837), .B(n1762), .C(n2557), .Y(n2043) );
  NAND2X1 U798 ( .A(\mem<10><10> ), .B(n1763), .Y(n2557) );
  OAI21X1 U799 ( .A(n1836), .B(n1762), .C(n2556), .Y(n2042) );
  NAND2X1 U800 ( .A(\mem<10><11> ), .B(n1763), .Y(n2556) );
  OAI21X1 U801 ( .A(n1835), .B(n1762), .C(n2555), .Y(n2041) );
  NAND2X1 U802 ( .A(\mem<10><12> ), .B(n1763), .Y(n2555) );
  OAI21X1 U803 ( .A(n1834), .B(n1762), .C(n2554), .Y(n2040) );
  NAND2X1 U804 ( .A(\mem<10><13> ), .B(n1763), .Y(n2554) );
  OAI21X1 U805 ( .A(n1833), .B(n1762), .C(n2553), .Y(n2039) );
  NAND2X1 U806 ( .A(\mem<10><14> ), .B(n1763), .Y(n2553) );
  OAI21X1 U807 ( .A(n1832), .B(n1762), .C(n2552), .Y(n2038) );
  NAND2X1 U808 ( .A(\mem<10><15> ), .B(n1763), .Y(n2552) );
  OAI21X1 U811 ( .A(n1862), .B(n1759), .C(n2551), .Y(n2037) );
  NAND2X1 U812 ( .A(\mem<9><0> ), .B(n1761), .Y(n2551) );
  OAI21X1 U813 ( .A(n1859), .B(n1759), .C(n2550), .Y(n2036) );
  NAND2X1 U814 ( .A(\mem<9><1> ), .B(n1761), .Y(n2550) );
  OAI21X1 U815 ( .A(n1856), .B(n1759), .C(n2549), .Y(n2035) );
  NAND2X1 U816 ( .A(\mem<9><2> ), .B(n1761), .Y(n2549) );
  OAI21X1 U817 ( .A(n1853), .B(n1759), .C(n2548), .Y(n2034) );
  NAND2X1 U818 ( .A(\mem<9><3> ), .B(n1761), .Y(n2548) );
  OAI21X1 U819 ( .A(n1850), .B(n1759), .C(n2547), .Y(n2033) );
  NAND2X1 U820 ( .A(\mem<9><4> ), .B(n1761), .Y(n2547) );
  OAI21X1 U821 ( .A(n1847), .B(n1759), .C(n2546), .Y(n2032) );
  NAND2X1 U822 ( .A(\mem<9><5> ), .B(n1761), .Y(n2546) );
  OAI21X1 U823 ( .A(n1844), .B(n1759), .C(n2545), .Y(n2031) );
  NAND2X1 U824 ( .A(\mem<9><6> ), .B(n1761), .Y(n2545) );
  OAI21X1 U825 ( .A(n1841), .B(n1759), .C(n2544), .Y(n2030) );
  NAND2X1 U826 ( .A(\mem<9><7> ), .B(n1761), .Y(n2544) );
  OAI21X1 U827 ( .A(n1839), .B(n1759), .C(n2543), .Y(n2029) );
  NAND2X1 U828 ( .A(\mem<9><8> ), .B(n1760), .Y(n2543) );
  OAI21X1 U829 ( .A(n1838), .B(n1759), .C(n2542), .Y(n2028) );
  NAND2X1 U830 ( .A(\mem<9><9> ), .B(n1760), .Y(n2542) );
  OAI21X1 U831 ( .A(n1837), .B(n1759), .C(n2541), .Y(n2027) );
  NAND2X1 U832 ( .A(\mem<9><10> ), .B(n1760), .Y(n2541) );
  OAI21X1 U833 ( .A(n1836), .B(n1759), .C(n2540), .Y(n2026) );
  NAND2X1 U834 ( .A(\mem<9><11> ), .B(n1760), .Y(n2540) );
  OAI21X1 U835 ( .A(n1835), .B(n1759), .C(n2539), .Y(n2025) );
  NAND2X1 U836 ( .A(\mem<9><12> ), .B(n1760), .Y(n2539) );
  OAI21X1 U837 ( .A(n1834), .B(n1759), .C(n2538), .Y(n2024) );
  NAND2X1 U838 ( .A(\mem<9><13> ), .B(n1760), .Y(n2538) );
  OAI21X1 U839 ( .A(n1833), .B(n1759), .C(n2537), .Y(n2023) );
  NAND2X1 U840 ( .A(\mem<9><14> ), .B(n1760), .Y(n2537) );
  OAI21X1 U841 ( .A(n1832), .B(n1759), .C(n2536), .Y(n2022) );
  NAND2X1 U842 ( .A(\mem<9><15> ), .B(n1760), .Y(n2536) );
  OAI21X1 U845 ( .A(n1862), .B(n1756), .C(n2535), .Y(n2021) );
  NAND2X1 U846 ( .A(\mem<8><0> ), .B(n1758), .Y(n2535) );
  OAI21X1 U847 ( .A(n1859), .B(n1756), .C(n2534), .Y(n2020) );
  NAND2X1 U848 ( .A(\mem<8><1> ), .B(n1758), .Y(n2534) );
  OAI21X1 U849 ( .A(n1856), .B(n1756), .C(n2533), .Y(n2019) );
  NAND2X1 U850 ( .A(\mem<8><2> ), .B(n1758), .Y(n2533) );
  OAI21X1 U851 ( .A(n1853), .B(n1756), .C(n2532), .Y(n2018) );
  NAND2X1 U852 ( .A(\mem<8><3> ), .B(n1758), .Y(n2532) );
  OAI21X1 U853 ( .A(n1850), .B(n1756), .C(n2531), .Y(n2017) );
  NAND2X1 U854 ( .A(\mem<8><4> ), .B(n1758), .Y(n2531) );
  OAI21X1 U855 ( .A(n1847), .B(n1756), .C(n2530), .Y(n2016) );
  NAND2X1 U856 ( .A(\mem<8><5> ), .B(n1758), .Y(n2530) );
  OAI21X1 U857 ( .A(n1844), .B(n1756), .C(n2529), .Y(n2015) );
  NAND2X1 U858 ( .A(\mem<8><6> ), .B(n1758), .Y(n2529) );
  OAI21X1 U859 ( .A(n1841), .B(n1756), .C(n2528), .Y(n2014) );
  NAND2X1 U860 ( .A(\mem<8><7> ), .B(n1758), .Y(n2528) );
  OAI21X1 U861 ( .A(n1839), .B(n1756), .C(n2527), .Y(n2013) );
  NAND2X1 U862 ( .A(\mem<8><8> ), .B(n1757), .Y(n2527) );
  OAI21X1 U863 ( .A(n1838), .B(n1756), .C(n2526), .Y(n2012) );
  NAND2X1 U864 ( .A(\mem<8><9> ), .B(n1757), .Y(n2526) );
  OAI21X1 U865 ( .A(n1837), .B(n1756), .C(n2525), .Y(n2011) );
  NAND2X1 U866 ( .A(\mem<8><10> ), .B(n1757), .Y(n2525) );
  OAI21X1 U867 ( .A(n1836), .B(n1756), .C(n2524), .Y(n2010) );
  NAND2X1 U868 ( .A(\mem<8><11> ), .B(n1757), .Y(n2524) );
  OAI21X1 U869 ( .A(n1835), .B(n1756), .C(n2523), .Y(n2009) );
  NAND2X1 U870 ( .A(\mem<8><12> ), .B(n1757), .Y(n2523) );
  OAI21X1 U871 ( .A(n1834), .B(n1756), .C(n2522), .Y(n2008) );
  NAND2X1 U872 ( .A(\mem<8><13> ), .B(n1757), .Y(n2522) );
  OAI21X1 U873 ( .A(n1833), .B(n1756), .C(n2521), .Y(n2007) );
  NAND2X1 U874 ( .A(\mem<8><14> ), .B(n1757), .Y(n2521) );
  OAI21X1 U875 ( .A(n1832), .B(n1756), .C(n2520), .Y(n2006) );
  NAND2X1 U876 ( .A(\mem<8><15> ), .B(n1757), .Y(n2520) );
  NAND3X1 U879 ( .A(n2777), .B(n1872), .C(n1870), .Y(n2519) );
  OAI21X1 U880 ( .A(n1862), .B(n1753), .C(n2518), .Y(n2005) );
  NAND2X1 U881 ( .A(\mem<7><0> ), .B(n1755), .Y(n2518) );
  OAI21X1 U882 ( .A(n1859), .B(n1753), .C(n2517), .Y(n2004) );
  NAND2X1 U883 ( .A(\mem<7><1> ), .B(n1755), .Y(n2517) );
  OAI21X1 U884 ( .A(n1856), .B(n1753), .C(n2516), .Y(n2003) );
  NAND2X1 U885 ( .A(\mem<7><2> ), .B(n1755), .Y(n2516) );
  OAI21X1 U886 ( .A(n1853), .B(n1753), .C(n2515), .Y(n2002) );
  NAND2X1 U887 ( .A(\mem<7><3> ), .B(n1755), .Y(n2515) );
  OAI21X1 U888 ( .A(n1850), .B(n1753), .C(n2514), .Y(n2001) );
  NAND2X1 U889 ( .A(\mem<7><4> ), .B(n1755), .Y(n2514) );
  OAI21X1 U890 ( .A(n1847), .B(n1753), .C(n2513), .Y(n2000) );
  NAND2X1 U891 ( .A(\mem<7><5> ), .B(n1755), .Y(n2513) );
  OAI21X1 U892 ( .A(n1844), .B(n1753), .C(n2512), .Y(n1999) );
  NAND2X1 U893 ( .A(\mem<7><6> ), .B(n1755), .Y(n2512) );
  OAI21X1 U894 ( .A(n1841), .B(n1753), .C(n2511), .Y(n1998) );
  NAND2X1 U895 ( .A(\mem<7><7> ), .B(n1755), .Y(n2511) );
  OAI21X1 U896 ( .A(n1839), .B(n1753), .C(n2510), .Y(n1997) );
  NAND2X1 U897 ( .A(\mem<7><8> ), .B(n1754), .Y(n2510) );
  OAI21X1 U898 ( .A(n1838), .B(n1753), .C(n2509), .Y(n1996) );
  NAND2X1 U899 ( .A(\mem<7><9> ), .B(n1754), .Y(n2509) );
  OAI21X1 U900 ( .A(n1837), .B(n1753), .C(n2508), .Y(n1995) );
  NAND2X1 U901 ( .A(\mem<7><10> ), .B(n1754), .Y(n2508) );
  OAI21X1 U902 ( .A(n1836), .B(n1753), .C(n2507), .Y(n1994) );
  NAND2X1 U903 ( .A(\mem<7><11> ), .B(n1754), .Y(n2507) );
  OAI21X1 U904 ( .A(n1835), .B(n1753), .C(n2506), .Y(n1993) );
  NAND2X1 U905 ( .A(\mem<7><12> ), .B(n1754), .Y(n2506) );
  OAI21X1 U906 ( .A(n1834), .B(n1753), .C(n2505), .Y(n1992) );
  NAND2X1 U907 ( .A(\mem<7><13> ), .B(n1754), .Y(n2505) );
  OAI21X1 U908 ( .A(n1833), .B(n1753), .C(n2504), .Y(n1991) );
  NAND2X1 U909 ( .A(\mem<7><14> ), .B(n1754), .Y(n2504) );
  OAI21X1 U910 ( .A(n1832), .B(n1753), .C(n2503), .Y(n1990) );
  NAND2X1 U911 ( .A(\mem<7><15> ), .B(n1754), .Y(n2503) );
  NOR3X1 U914 ( .A(n1867), .B(n1865), .C(n1869), .Y(n2898) );
  OAI21X1 U915 ( .A(n1862), .B(n1750), .C(n2502), .Y(n1989) );
  NAND2X1 U916 ( .A(\mem<6><0> ), .B(n1752), .Y(n2502) );
  OAI21X1 U917 ( .A(n1859), .B(n1750), .C(n2501), .Y(n1988) );
  NAND2X1 U918 ( .A(\mem<6><1> ), .B(n1752), .Y(n2501) );
  OAI21X1 U919 ( .A(n1856), .B(n1750), .C(n2500), .Y(n1987) );
  NAND2X1 U920 ( .A(\mem<6><2> ), .B(n1752), .Y(n2500) );
  OAI21X1 U921 ( .A(n1853), .B(n1750), .C(n2499), .Y(n1986) );
  NAND2X1 U922 ( .A(\mem<6><3> ), .B(n1752), .Y(n2499) );
  OAI21X1 U923 ( .A(n1850), .B(n1750), .C(n2498), .Y(n1985) );
  NAND2X1 U924 ( .A(\mem<6><4> ), .B(n1752), .Y(n2498) );
  OAI21X1 U925 ( .A(n1847), .B(n1750), .C(n2497), .Y(n1984) );
  NAND2X1 U926 ( .A(\mem<6><5> ), .B(n1752), .Y(n2497) );
  OAI21X1 U927 ( .A(n1844), .B(n1750), .C(n2496), .Y(n1983) );
  NAND2X1 U928 ( .A(\mem<6><6> ), .B(n1752), .Y(n2496) );
  OAI21X1 U929 ( .A(n1841), .B(n1750), .C(n2495), .Y(n1982) );
  NAND2X1 U930 ( .A(\mem<6><7> ), .B(n1752), .Y(n2495) );
  OAI21X1 U931 ( .A(n1839), .B(n1750), .C(n2494), .Y(n1981) );
  NAND2X1 U932 ( .A(\mem<6><8> ), .B(n1751), .Y(n2494) );
  OAI21X1 U933 ( .A(n1838), .B(n1750), .C(n2493), .Y(n1980) );
  NAND2X1 U934 ( .A(\mem<6><9> ), .B(n1751), .Y(n2493) );
  OAI21X1 U935 ( .A(n1837), .B(n1750), .C(n2492), .Y(n1979) );
  NAND2X1 U936 ( .A(\mem<6><10> ), .B(n1751), .Y(n2492) );
  OAI21X1 U937 ( .A(n1836), .B(n1750), .C(n2491), .Y(n1978) );
  NAND2X1 U938 ( .A(\mem<6><11> ), .B(n1751), .Y(n2491) );
  OAI21X1 U939 ( .A(n1835), .B(n1750), .C(n2490), .Y(n1977) );
  NAND2X1 U940 ( .A(\mem<6><12> ), .B(n1751), .Y(n2490) );
  OAI21X1 U941 ( .A(n1834), .B(n1750), .C(n2489), .Y(n1976) );
  NAND2X1 U942 ( .A(\mem<6><13> ), .B(n1751), .Y(n2489) );
  OAI21X1 U943 ( .A(n1833), .B(n1750), .C(n2488), .Y(n1975) );
  NAND2X1 U944 ( .A(\mem<6><14> ), .B(n1751), .Y(n2488) );
  OAI21X1 U945 ( .A(n1832), .B(n1750), .C(n2487), .Y(n1974) );
  NAND2X1 U946 ( .A(\mem<6><15> ), .B(n1751), .Y(n2487) );
  NOR3X1 U949 ( .A(n1867), .B(n1864), .C(n1869), .Y(n2881) );
  OAI21X1 U950 ( .A(n1863), .B(n1747), .C(n2486), .Y(n1973) );
  NAND2X1 U951 ( .A(\mem<5><0> ), .B(n1749), .Y(n2486) );
  OAI21X1 U952 ( .A(n1860), .B(n1747), .C(n2485), .Y(n1972) );
  NAND2X1 U953 ( .A(\mem<5><1> ), .B(n1749), .Y(n2485) );
  OAI21X1 U954 ( .A(n1857), .B(n1747), .C(n2484), .Y(n1971) );
  NAND2X1 U955 ( .A(\mem<5><2> ), .B(n1749), .Y(n2484) );
  OAI21X1 U956 ( .A(n1854), .B(n1747), .C(n2483), .Y(n1970) );
  NAND2X1 U957 ( .A(\mem<5><3> ), .B(n1749), .Y(n2483) );
  OAI21X1 U958 ( .A(n1851), .B(n1747), .C(n2482), .Y(n1969) );
  NAND2X1 U959 ( .A(\mem<5><4> ), .B(n1749), .Y(n2482) );
  OAI21X1 U960 ( .A(n1848), .B(n1747), .C(n2481), .Y(n1968) );
  NAND2X1 U961 ( .A(\mem<5><5> ), .B(n1749), .Y(n2481) );
  OAI21X1 U962 ( .A(n1845), .B(n1747), .C(n2480), .Y(n1967) );
  NAND2X1 U963 ( .A(\mem<5><6> ), .B(n1749), .Y(n2480) );
  OAI21X1 U964 ( .A(n1842), .B(n1747), .C(n2479), .Y(n1966) );
  NAND2X1 U965 ( .A(\mem<5><7> ), .B(n1749), .Y(n2479) );
  OAI21X1 U966 ( .A(n1839), .B(n1747), .C(n2478), .Y(n1965) );
  NAND2X1 U967 ( .A(\mem<5><8> ), .B(n1748), .Y(n2478) );
  OAI21X1 U968 ( .A(n1838), .B(n1747), .C(n2477), .Y(n1964) );
  NAND2X1 U969 ( .A(\mem<5><9> ), .B(n1748), .Y(n2477) );
  OAI21X1 U970 ( .A(n1837), .B(n1747), .C(n2476), .Y(n1963) );
  NAND2X1 U971 ( .A(\mem<5><10> ), .B(n1748), .Y(n2476) );
  OAI21X1 U972 ( .A(n1836), .B(n1747), .C(n2475), .Y(n1962) );
  NAND2X1 U973 ( .A(\mem<5><11> ), .B(n1748), .Y(n2475) );
  OAI21X1 U974 ( .A(n1835), .B(n1747), .C(n2474), .Y(n1961) );
  NAND2X1 U975 ( .A(\mem<5><12> ), .B(n1748), .Y(n2474) );
  OAI21X1 U976 ( .A(n1834), .B(n1747), .C(n2473), .Y(n1960) );
  NAND2X1 U977 ( .A(\mem<5><13> ), .B(n1748), .Y(n2473) );
  OAI21X1 U978 ( .A(n1833), .B(n1747), .C(n2472), .Y(n1959) );
  NAND2X1 U979 ( .A(\mem<5><14> ), .B(n1748), .Y(n2472) );
  OAI21X1 U980 ( .A(n1832), .B(n1747), .C(n2471), .Y(n1958) );
  NAND2X1 U981 ( .A(\mem<5><15> ), .B(n1748), .Y(n2471) );
  NOR3X1 U984 ( .A(n1865), .B(n1866), .C(n1869), .Y(n2864) );
  OAI21X1 U985 ( .A(n1863), .B(n1744), .C(n2470), .Y(n1957) );
  NAND2X1 U986 ( .A(\mem<4><0> ), .B(n1746), .Y(n2470) );
  OAI21X1 U987 ( .A(n1860), .B(n1744), .C(n2469), .Y(n1956) );
  NAND2X1 U988 ( .A(\mem<4><1> ), .B(n1746), .Y(n2469) );
  OAI21X1 U989 ( .A(n1857), .B(n1744), .C(n2468), .Y(n1955) );
  NAND2X1 U990 ( .A(\mem<4><2> ), .B(n1746), .Y(n2468) );
  OAI21X1 U991 ( .A(n1854), .B(n1744), .C(n2467), .Y(n1954) );
  NAND2X1 U992 ( .A(\mem<4><3> ), .B(n1746), .Y(n2467) );
  OAI21X1 U993 ( .A(n1851), .B(n1744), .C(n2466), .Y(n1953) );
  NAND2X1 U994 ( .A(\mem<4><4> ), .B(n1746), .Y(n2466) );
  OAI21X1 U995 ( .A(n1848), .B(n1744), .C(n2465), .Y(n1952) );
  NAND2X1 U996 ( .A(\mem<4><5> ), .B(n1746), .Y(n2465) );
  OAI21X1 U997 ( .A(n1845), .B(n1744), .C(n2464), .Y(n1951) );
  NAND2X1 U998 ( .A(\mem<4><6> ), .B(n1746), .Y(n2464) );
  OAI21X1 U999 ( .A(n1842), .B(n1744), .C(n2463), .Y(n1950) );
  NAND2X1 U1000 ( .A(\mem<4><7> ), .B(n1746), .Y(n2463) );
  OAI21X1 U1001 ( .A(n1839), .B(n1744), .C(n2462), .Y(n1949) );
  NAND2X1 U1002 ( .A(\mem<4><8> ), .B(n1745), .Y(n2462) );
  OAI21X1 U1003 ( .A(n1838), .B(n1744), .C(n2461), .Y(n1948) );
  NAND2X1 U1004 ( .A(\mem<4><9> ), .B(n1745), .Y(n2461) );
  OAI21X1 U1005 ( .A(n1837), .B(n1744), .C(n2460), .Y(n1947) );
  NAND2X1 U1006 ( .A(\mem<4><10> ), .B(n1745), .Y(n2460) );
  OAI21X1 U1007 ( .A(n1836), .B(n1744), .C(n2459), .Y(n1946) );
  NAND2X1 U1008 ( .A(\mem<4><11> ), .B(n1745), .Y(n2459) );
  OAI21X1 U1009 ( .A(n1835), .B(n1744), .C(n2458), .Y(n1945) );
  NAND2X1 U1010 ( .A(\mem<4><12> ), .B(n1745), .Y(n2458) );
  OAI21X1 U1011 ( .A(n1834), .B(n1744), .C(n2457), .Y(n1944) );
  NAND2X1 U1012 ( .A(\mem<4><13> ), .B(n1745), .Y(n2457) );
  OAI21X1 U1013 ( .A(n1833), .B(n1744), .C(n2456), .Y(n1943) );
  NAND2X1 U1014 ( .A(\mem<4><14> ), .B(n1745), .Y(n2456) );
  OAI21X1 U1015 ( .A(n1832), .B(n1744), .C(n2455), .Y(n1942) );
  NAND2X1 U1016 ( .A(\mem<4><15> ), .B(n1745), .Y(n2455) );
  NOR3X1 U1019 ( .A(n1864), .B(n1866), .C(n1869), .Y(n2847) );
  OAI21X1 U1020 ( .A(n1863), .B(n1741), .C(n2454), .Y(n1941) );
  NAND2X1 U1021 ( .A(\mem<3><0> ), .B(n1743), .Y(n2454) );
  OAI21X1 U1022 ( .A(n1860), .B(n1741), .C(n2453), .Y(n1940) );
  NAND2X1 U1023 ( .A(\mem<3><1> ), .B(n1743), .Y(n2453) );
  OAI21X1 U1024 ( .A(n1857), .B(n1741), .C(n2452), .Y(n1939) );
  NAND2X1 U1025 ( .A(\mem<3><2> ), .B(n1743), .Y(n2452) );
  OAI21X1 U1026 ( .A(n1854), .B(n1741), .C(n2451), .Y(n1938) );
  NAND2X1 U1027 ( .A(\mem<3><3> ), .B(n1743), .Y(n2451) );
  OAI21X1 U1028 ( .A(n1851), .B(n1741), .C(n2450), .Y(n1937) );
  NAND2X1 U1029 ( .A(\mem<3><4> ), .B(n1743), .Y(n2450) );
  OAI21X1 U1030 ( .A(n1848), .B(n1741), .C(n2449), .Y(n1936) );
  NAND2X1 U1031 ( .A(\mem<3><5> ), .B(n1743), .Y(n2449) );
  OAI21X1 U1032 ( .A(n1845), .B(n1741), .C(n2448), .Y(n1935) );
  NAND2X1 U1033 ( .A(\mem<3><6> ), .B(n1743), .Y(n2448) );
  OAI21X1 U1034 ( .A(n1842), .B(n1741), .C(n2447), .Y(n1934) );
  NAND2X1 U1035 ( .A(\mem<3><7> ), .B(n1743), .Y(n2447) );
  OAI21X1 U1036 ( .A(n1839), .B(n1741), .C(n2446), .Y(n1933) );
  NAND2X1 U1037 ( .A(\mem<3><8> ), .B(n1742), .Y(n2446) );
  OAI21X1 U1038 ( .A(n1838), .B(n1741), .C(n2445), .Y(n1932) );
  NAND2X1 U1039 ( .A(\mem<3><9> ), .B(n1742), .Y(n2445) );
  OAI21X1 U1040 ( .A(n1837), .B(n1741), .C(n2444), .Y(n1931) );
  NAND2X1 U1041 ( .A(\mem<3><10> ), .B(n1742), .Y(n2444) );
  OAI21X1 U1042 ( .A(n1836), .B(n1741), .C(n2443), .Y(n1930) );
  NAND2X1 U1043 ( .A(\mem<3><11> ), .B(n1742), .Y(n2443) );
  OAI21X1 U1044 ( .A(n1835), .B(n1741), .C(n2442), .Y(n1929) );
  NAND2X1 U1045 ( .A(\mem<3><12> ), .B(n1742), .Y(n2442) );
  OAI21X1 U1046 ( .A(n1834), .B(n1741), .C(n2441), .Y(n1928) );
  NAND2X1 U1047 ( .A(\mem<3><13> ), .B(n1742), .Y(n2441) );
  OAI21X1 U1048 ( .A(n1833), .B(n1741), .C(n2440), .Y(n1927) );
  NAND2X1 U1049 ( .A(\mem<3><14> ), .B(n1742), .Y(n2440) );
  OAI21X1 U1050 ( .A(n1832), .B(n1741), .C(n2439), .Y(n1926) );
  NAND2X1 U1051 ( .A(\mem<3><15> ), .B(n1742), .Y(n2439) );
  NOR3X1 U1054 ( .A(n1865), .B(n1868), .C(n1867), .Y(n2830) );
  OAI21X1 U1055 ( .A(n1863), .B(n1738), .C(n2438), .Y(n1925) );
  NAND2X1 U1056 ( .A(\mem<2><0> ), .B(n1740), .Y(n2438) );
  OAI21X1 U1057 ( .A(n1860), .B(n1738), .C(n2437), .Y(n1924) );
  NAND2X1 U1058 ( .A(\mem<2><1> ), .B(n1740), .Y(n2437) );
  OAI21X1 U1059 ( .A(n1857), .B(n1738), .C(n2436), .Y(n1923) );
  NAND2X1 U1060 ( .A(\mem<2><2> ), .B(n1740), .Y(n2436) );
  OAI21X1 U1061 ( .A(n1854), .B(n1738), .C(n2435), .Y(n1922) );
  NAND2X1 U1062 ( .A(\mem<2><3> ), .B(n1740), .Y(n2435) );
  OAI21X1 U1063 ( .A(n1851), .B(n1738), .C(n2434), .Y(n1921) );
  NAND2X1 U1064 ( .A(\mem<2><4> ), .B(n1740), .Y(n2434) );
  OAI21X1 U1065 ( .A(n1848), .B(n1738), .C(n2433), .Y(n1920) );
  NAND2X1 U1066 ( .A(\mem<2><5> ), .B(n1740), .Y(n2433) );
  OAI21X1 U1067 ( .A(n1845), .B(n1738), .C(n2432), .Y(n1919) );
  NAND2X1 U1068 ( .A(\mem<2><6> ), .B(n1740), .Y(n2432) );
  OAI21X1 U1069 ( .A(n1842), .B(n1738), .C(n2431), .Y(n1918) );
  NAND2X1 U1070 ( .A(\mem<2><7> ), .B(n1740), .Y(n2431) );
  OAI21X1 U1071 ( .A(n1839), .B(n1738), .C(n2430), .Y(n1917) );
  NAND2X1 U1072 ( .A(\mem<2><8> ), .B(n1739), .Y(n2430) );
  OAI21X1 U1073 ( .A(n1838), .B(n1738), .C(n2429), .Y(n1916) );
  NAND2X1 U1074 ( .A(\mem<2><9> ), .B(n1739), .Y(n2429) );
  OAI21X1 U1075 ( .A(n1837), .B(n1738), .C(n2428), .Y(n1915) );
  NAND2X1 U1076 ( .A(\mem<2><10> ), .B(n1739), .Y(n2428) );
  OAI21X1 U1077 ( .A(n1836), .B(n1738), .C(n2427), .Y(n1914) );
  NAND2X1 U1078 ( .A(\mem<2><11> ), .B(n1739), .Y(n2427) );
  OAI21X1 U1079 ( .A(n1835), .B(n1738), .C(n2426), .Y(n1913) );
  NAND2X1 U1080 ( .A(\mem<2><12> ), .B(n1739), .Y(n2426) );
  OAI21X1 U1081 ( .A(n1834), .B(n1738), .C(n2425), .Y(n1912) );
  NAND2X1 U1082 ( .A(\mem<2><13> ), .B(n1739), .Y(n2425) );
  OAI21X1 U1083 ( .A(n1833), .B(n1738), .C(n2424), .Y(n1911) );
  NAND2X1 U1084 ( .A(\mem<2><14> ), .B(n1739), .Y(n2424) );
  OAI21X1 U1085 ( .A(n1832), .B(n1738), .C(n2423), .Y(n1910) );
  NAND2X1 U1086 ( .A(\mem<2><15> ), .B(n1739), .Y(n2423) );
  NOR3X1 U1089 ( .A(n1864), .B(n1868), .C(n1867), .Y(n2813) );
  OAI21X1 U1090 ( .A(n1863), .B(n1735), .C(n2422), .Y(n1909) );
  NAND2X1 U1091 ( .A(\mem<1><0> ), .B(n1737), .Y(n2422) );
  OAI21X1 U1092 ( .A(n1860), .B(n1735), .C(n2421), .Y(n1908) );
  NAND2X1 U1093 ( .A(\mem<1><1> ), .B(n1737), .Y(n2421) );
  OAI21X1 U1094 ( .A(n1857), .B(n1735), .C(n2420), .Y(n1907) );
  NAND2X1 U1095 ( .A(\mem<1><2> ), .B(n1737), .Y(n2420) );
  OAI21X1 U1096 ( .A(n1854), .B(n1735), .C(n2419), .Y(n1906) );
  NAND2X1 U1097 ( .A(\mem<1><3> ), .B(n1737), .Y(n2419) );
  OAI21X1 U1098 ( .A(n1851), .B(n1735), .C(n2418), .Y(n1905) );
  NAND2X1 U1099 ( .A(\mem<1><4> ), .B(n1737), .Y(n2418) );
  OAI21X1 U1100 ( .A(n1848), .B(n1735), .C(n2417), .Y(n1904) );
  NAND2X1 U1101 ( .A(\mem<1><5> ), .B(n1737), .Y(n2417) );
  OAI21X1 U1102 ( .A(n1845), .B(n1735), .C(n2416), .Y(n1903) );
  NAND2X1 U1103 ( .A(\mem<1><6> ), .B(n1737), .Y(n2416) );
  OAI21X1 U1104 ( .A(n1842), .B(n1735), .C(n2415), .Y(n1902) );
  NAND2X1 U1105 ( .A(\mem<1><7> ), .B(n1737), .Y(n2415) );
  OAI21X1 U1106 ( .A(n1839), .B(n1735), .C(n2414), .Y(n1901) );
  NAND2X1 U1107 ( .A(\mem<1><8> ), .B(n1736), .Y(n2414) );
  OAI21X1 U1108 ( .A(n1838), .B(n1735), .C(n2413), .Y(n1900) );
  NAND2X1 U1109 ( .A(\mem<1><9> ), .B(n1736), .Y(n2413) );
  OAI21X1 U1110 ( .A(n1837), .B(n1735), .C(n2412), .Y(n1899) );
  NAND2X1 U1111 ( .A(\mem<1><10> ), .B(n1736), .Y(n2412) );
  OAI21X1 U1112 ( .A(n1836), .B(n1735), .C(n2411), .Y(n1898) );
  NAND2X1 U1113 ( .A(\mem<1><11> ), .B(n1736), .Y(n2411) );
  OAI21X1 U1114 ( .A(n1835), .B(n1735), .C(n2410), .Y(n1897) );
  NAND2X1 U1115 ( .A(\mem<1><12> ), .B(n1736), .Y(n2410) );
  OAI21X1 U1116 ( .A(n1834), .B(n1735), .C(n2409), .Y(n1896) );
  NAND2X1 U1117 ( .A(\mem<1><13> ), .B(n1736), .Y(n2409) );
  OAI21X1 U1118 ( .A(n1833), .B(n1735), .C(n2408), .Y(n1895) );
  NAND2X1 U1119 ( .A(\mem<1><14> ), .B(n1736), .Y(n2408) );
  OAI21X1 U1120 ( .A(n1832), .B(n1735), .C(n2407), .Y(n1894) );
  NAND2X1 U1121 ( .A(\mem<1><15> ), .B(n1736), .Y(n2407) );
  NOR3X1 U1124 ( .A(n1866), .B(n1868), .C(n1865), .Y(n2796) );
  OAI21X1 U1125 ( .A(n1863), .B(n1732), .C(n2406), .Y(n1893) );
  NAND2X1 U1126 ( .A(\mem<0><0> ), .B(n1734), .Y(n2406) );
  OAI21X1 U1128 ( .A(n1860), .B(n1732), .C(n2405), .Y(n1892) );
  NAND2X1 U1129 ( .A(\mem<0><1> ), .B(n1734), .Y(n2405) );
  OAI21X1 U1131 ( .A(n1857), .B(n1732), .C(n2404), .Y(n1891) );
  NAND2X1 U1132 ( .A(\mem<0><2> ), .B(n1734), .Y(n2404) );
  OAI21X1 U1134 ( .A(n1854), .B(n1732), .C(n2403), .Y(n1890) );
  NAND2X1 U1135 ( .A(\mem<0><3> ), .B(n1734), .Y(n2403) );
  OAI21X1 U1137 ( .A(n1851), .B(n1732), .C(n2402), .Y(n1889) );
  NAND2X1 U1138 ( .A(\mem<0><4> ), .B(n1734), .Y(n2402) );
  OAI21X1 U1140 ( .A(n1848), .B(n1732), .C(n2401), .Y(n1888) );
  NAND2X1 U1141 ( .A(\mem<0><5> ), .B(n1734), .Y(n2401) );
  OAI21X1 U1143 ( .A(n1845), .B(n1732), .C(n2400), .Y(n1887) );
  NAND2X1 U1144 ( .A(\mem<0><6> ), .B(n1734), .Y(n2400) );
  OAI21X1 U1146 ( .A(n1842), .B(n1732), .C(n2399), .Y(n1886) );
  NAND2X1 U1147 ( .A(\mem<0><7> ), .B(n1734), .Y(n2399) );
  OAI21X1 U1149 ( .A(n1839), .B(n1732), .C(n2398), .Y(n1885) );
  NAND2X1 U1150 ( .A(\mem<0><8> ), .B(n1733), .Y(n2398) );
  OAI21X1 U1152 ( .A(n1838), .B(n1732), .C(n2397), .Y(n1884) );
  NAND2X1 U1153 ( .A(\mem<0><9> ), .B(n1733), .Y(n2397) );
  OAI21X1 U1155 ( .A(n1837), .B(n1732), .C(n2396), .Y(n1883) );
  NAND2X1 U1156 ( .A(\mem<0><10> ), .B(n1733), .Y(n2396) );
  OAI21X1 U1158 ( .A(n1836), .B(n1732), .C(n2395), .Y(n1882) );
  NAND2X1 U1159 ( .A(\mem<0><11> ), .B(n1733), .Y(n2395) );
  OAI21X1 U1161 ( .A(n1835), .B(n1732), .C(n2394), .Y(n1881) );
  NAND2X1 U1162 ( .A(\mem<0><12> ), .B(n1733), .Y(n2394) );
  OAI21X1 U1164 ( .A(n1834), .B(n1732), .C(n2393), .Y(n1880) );
  NAND2X1 U1165 ( .A(\mem<0><13> ), .B(n1733), .Y(n2393) );
  OAI21X1 U1167 ( .A(n1833), .B(n1732), .C(n2392), .Y(n1879) );
  NAND2X1 U1168 ( .A(\mem<0><14> ), .B(n1733), .Y(n2392) );
  OAI21X1 U1170 ( .A(n1832), .B(n1732), .C(n2391), .Y(n1878) );
  NAND2X1 U1171 ( .A(\mem<0><15> ), .B(n1733), .Y(n2391) );
  NOR3X1 U1174 ( .A(n1866), .B(n1868), .C(n1864), .Y(n2779) );
  NAND3X1 U1175 ( .A(n1871), .B(n1872), .C(n2777), .Y(n2390) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2777) );
  INVX1 U3 ( .A(n8), .Y(n1) );
  INVX2 U4 ( .A(n1717), .Y(n1729) );
  INVX2 U5 ( .A(n1717), .Y(n1730) );
  INVX2 U6 ( .A(n1717), .Y(n1723) );
  INVX2 U7 ( .A(n1717), .Y(n1725) );
  INVX2 U8 ( .A(n1717), .Y(n1724) );
  AND2X2 U9 ( .A(\data_in<8> ), .B(n1830), .Y(n58) );
  AND2X2 U10 ( .A(\data_in<10> ), .B(n1830), .Y(n54) );
  AND2X2 U11 ( .A(\data_in<12> ), .B(n1830), .Y(n50) );
  AND2X2 U12 ( .A(\data_in<14> ), .B(n1830), .Y(n47) );
  AND2X2 U13 ( .A(\data_in<9> ), .B(n1829), .Y(n56) );
  AND2X2 U14 ( .A(\data_in<11> ), .B(n1829), .Y(n52) );
  AND2X2 U15 ( .A(\data_in<13> ), .B(n1829), .Y(n48) );
  AND2X2 U16 ( .A(\data_in<15> ), .B(n1829), .Y(n45) );
  INVX1 U17 ( .A(n10), .Y(n2) );
  INVX1 U18 ( .A(n1865), .Y(n1731) );
  INVX1 U19 ( .A(n1706), .Y(n1707) );
  INVX1 U20 ( .A(n1706), .Y(n1708) );
  INVX1 U21 ( .A(n1718), .Y(n1722) );
  INVX1 U22 ( .A(n1706), .Y(n1709) );
  INVX1 U23 ( .A(n1718), .Y(n1726) );
  INVX1 U24 ( .A(n1718), .Y(n1727) );
  INVX1 U25 ( .A(n1704), .Y(n1712) );
  INVX1 U26 ( .A(n1704), .Y(n1713) );
  INVX1 U27 ( .A(n1704), .Y(n1714) );
  INVX2 U28 ( .A(n1706), .Y(n1715) );
  INVX1 U29 ( .A(n1718), .Y(n1728) );
  INVX2 U30 ( .A(n1704), .Y(n1716) );
  INVX1 U31 ( .A(rst), .Y(n1873) );
  INVX1 U32 ( .A(n1699), .Y(n1701) );
  INVX1 U33 ( .A(n1866), .Y(n1705) );
  INVX2 U34 ( .A(n1705), .Y(n1710) );
  INVX1 U35 ( .A(n1705), .Y(n1711) );
  INVX1 U36 ( .A(n1731), .Y(n1718) );
  INVX2 U37 ( .A(n1717), .Y(n1720) );
  INVX2 U38 ( .A(n1717), .Y(n1719) );
  INVX2 U39 ( .A(n1718), .Y(n1721) );
  INVX1 U40 ( .A(n1865), .Y(n1864) );
  INVX2 U41 ( .A(n1864), .Y(n1717) );
  INVX1 U42 ( .A(N13), .Y(n1871) );
  INVX1 U43 ( .A(n1871), .Y(n1697) );
  INVX1 U44 ( .A(n1871), .Y(n1696) );
  INVX1 U45 ( .A(n1868), .Y(n1698) );
  INVX1 U46 ( .A(n1698), .Y(n1703) );
  INVX1 U47 ( .A(n1698), .Y(n1702) );
  INVX1 U48 ( .A(n1867), .Y(n1866) );
  INVX1 U49 ( .A(N14), .Y(n1872) );
  INVX1 U50 ( .A(n101), .Y(n1732) );
  INVX1 U51 ( .A(n118), .Y(n1735) );
  INVX1 U52 ( .A(n177), .Y(n1756) );
  INVX1 U53 ( .A(n194), .Y(n1759) );
  INVX1 U54 ( .A(n253), .Y(n1780) );
  INVX1 U55 ( .A(n269), .Y(n1783) );
  INVX1 U56 ( .A(n1872), .Y(n1695) );
  INVX1 U57 ( .A(n287), .Y(n1789) );
  INVX1 U58 ( .A(n289), .Y(n1792) );
  INVX1 U59 ( .A(n305), .Y(n1795) );
  INVX1 U60 ( .A(n307), .Y(n1798) );
  INVX1 U93 ( .A(n323), .Y(n1801) );
  INVX1 U94 ( .A(n325), .Y(n1804) );
  INVX1 U127 ( .A(n341), .Y(n1807) );
  INVX1 U128 ( .A(n343), .Y(n1810) );
  INVX1 U161 ( .A(n360), .Y(n1813) );
  INVX1 U162 ( .A(n362), .Y(n1816) );
  INVX1 U195 ( .A(n378), .Y(n1819) );
  INVX1 U196 ( .A(n380), .Y(n1822) );
  INVX1 U229 ( .A(n396), .Y(n1825) );
  INVX4 U230 ( .A(n2899), .Y(n1831) );
  INVX1 U263 ( .A(n120), .Y(n1738) );
  INVX1 U264 ( .A(n137), .Y(n1741) );
  INVX1 U297 ( .A(n139), .Y(n1744) );
  INVX1 U298 ( .A(n156), .Y(n1747) );
  INVX1 U331 ( .A(n158), .Y(n1750) );
  INVX1 U332 ( .A(n175), .Y(n1753) );
  INVX1 U366 ( .A(n196), .Y(n1762) );
  INVX1 U367 ( .A(n215), .Y(n1765) );
  INVX1 U400 ( .A(n217), .Y(n1768) );
  INVX1 U401 ( .A(n233), .Y(n1771) );
  INVX1 U434 ( .A(n235), .Y(n1774) );
  INVX1 U435 ( .A(n251), .Y(n1777) );
  INVX1 U468 ( .A(n271), .Y(n1786) );
  INVX1 U469 ( .A(n1868), .Y(n1699) );
  INVX1 U502 ( .A(n1699), .Y(n1700) );
  INVX1 U503 ( .A(n1866), .Y(n1704) );
  INVX1 U536 ( .A(n1866), .Y(n1706) );
  INVX1 U537 ( .A(n8), .Y(n3) );
  INVX1 U570 ( .A(write), .Y(n4) );
  INVX1 U571 ( .A(n10), .Y(n5) );
  INVX1 U604 ( .A(n8), .Y(n6) );
  INVX1 U605 ( .A(n8), .Y(n7) );
  AND2X2 U639 ( .A(n9), .B(n1873), .Y(n8) );
  INVX1 U640 ( .A(write), .Y(n9) );
  AND2X2 U673 ( .A(n4), .B(n1873), .Y(n10) );
  INVX1 U674 ( .A(n10), .Y(n11) );
  INVX1 U707 ( .A(n10), .Y(n12) );
  OR2X2 U708 ( .A(n3), .B(n1694), .Y(n43) );
  OR2X2 U741 ( .A(n7), .B(n1693), .Y(n41) );
  OR2X2 U742 ( .A(n6), .B(n1679), .Y(n13) );
  INVX1 U775 ( .A(n13), .Y(\data_out<0> ) );
  OR2X2 U776 ( .A(n11), .B(n1680), .Y(n15) );
  INVX1 U809 ( .A(n15), .Y(\data_out<1> ) );
  OR2X2 U810 ( .A(n1), .B(n1681), .Y(n17) );
  INVX1 U843 ( .A(n17), .Y(\data_out<2> ) );
  OR2X2 U844 ( .A(n6), .B(n1682), .Y(n19) );
  INVX1 U877 ( .A(n19), .Y(\data_out<3> ) );
  OR2X2 U878 ( .A(n2), .B(n1683), .Y(n21) );
  INVX1 U912 ( .A(n21), .Y(\data_out<4> ) );
  OR2X2 U913 ( .A(n7), .B(n1684), .Y(n23) );
  INVX1 U947 ( .A(n23), .Y(\data_out<5> ) );
  OR2X2 U948 ( .A(n12), .B(n1685), .Y(n25) );
  INVX1 U982 ( .A(n25), .Y(\data_out<6> ) );
  OR2X2 U983 ( .A(n2), .B(n1686), .Y(n27) );
  INVX1 U1017 ( .A(n27), .Y(\data_out<7> ) );
  OR2X2 U1018 ( .A(n12), .B(n1687), .Y(n29) );
  INVX1 U1052 ( .A(n29), .Y(\data_out<8> ) );
  OR2X2 U1053 ( .A(n5), .B(n1688), .Y(n31) );
  INVX1 U1087 ( .A(n31), .Y(\data_out<9> ) );
  OR2X2 U1088 ( .A(n3), .B(n1689), .Y(n33) );
  INVX1 U1122 ( .A(n33), .Y(\data_out<10> ) );
  OR2X2 U1123 ( .A(n11), .B(n1690), .Y(n35) );
  INVX1 U1127 ( .A(n35), .Y(\data_out<11> ) );
  OR2X2 U1130 ( .A(n1), .B(n1691), .Y(n37) );
  INVX1 U1133 ( .A(n37), .Y(\data_out<12> ) );
  OR2X2 U1136 ( .A(n5), .B(n1692), .Y(n39) );
  INVX1 U1139 ( .A(n39), .Y(\data_out<13> ) );
  INVX1 U1142 ( .A(n41), .Y(\data_out<14> ) );
  INVX1 U1145 ( .A(n43), .Y(\data_out<15> ) );
  BUFX2 U1148 ( .A(n414), .Y(n1733) );
  BUFX2 U1151 ( .A(n414), .Y(n1734) );
  BUFX2 U1154 ( .A(n432), .Y(n1736) );
  BUFX2 U1157 ( .A(n432), .Y(n1737) );
  BUFX2 U1160 ( .A(n450), .Y(n1739) );
  BUFX2 U1163 ( .A(n450), .Y(n1740) );
  BUFX2 U1166 ( .A(n468), .Y(n1742) );
  BUFX2 U1169 ( .A(n468), .Y(n1743) );
  BUFX2 U1172 ( .A(n486), .Y(n1745) );
  BUFX2 U1173 ( .A(n486), .Y(n1746) );
  BUFX2 U1177 ( .A(n505), .Y(n1748) );
  BUFX2 U1178 ( .A(n505), .Y(n1749) );
  BUFX2 U1179 ( .A(n523), .Y(n1751) );
  BUFX2 U1180 ( .A(n523), .Y(n1752) );
  BUFX2 U1181 ( .A(n541), .Y(n1754) );
  BUFX2 U1182 ( .A(n541), .Y(n1755) );
  BUFX2 U1183 ( .A(n559), .Y(n1757) );
  BUFX2 U1184 ( .A(n559), .Y(n1758) );
  BUFX2 U1185 ( .A(n577), .Y(n1760) );
  BUFX2 U1186 ( .A(n577), .Y(n1761) );
  BUFX2 U1187 ( .A(n595), .Y(n1763) );
  BUFX2 U1188 ( .A(n595), .Y(n1764) );
  BUFX2 U1189 ( .A(n613), .Y(n1766) );
  BUFX2 U1190 ( .A(n613), .Y(n1767) );
  BUFX2 U1191 ( .A(n631), .Y(n1769) );
  BUFX2 U1192 ( .A(n631), .Y(n1770) );
  BUFX2 U1193 ( .A(n650), .Y(n1772) );
  BUFX2 U1194 ( .A(n650), .Y(n1773) );
  BUFX2 U1195 ( .A(n1164), .Y(n1775) );
  BUFX2 U1196 ( .A(n1164), .Y(n1776) );
  BUFX2 U1197 ( .A(n1166), .Y(n1778) );
  BUFX2 U1198 ( .A(n1166), .Y(n1779) );
  BUFX2 U1199 ( .A(n1168), .Y(n1781) );
  BUFX2 U1200 ( .A(n1168), .Y(n1782) );
  BUFX2 U1201 ( .A(n1170), .Y(n1784) );
  BUFX2 U1202 ( .A(n1170), .Y(n1785) );
  BUFX2 U1203 ( .A(n1172), .Y(n1787) );
  BUFX2 U1204 ( .A(n1172), .Y(n1788) );
  BUFX2 U1205 ( .A(n1174), .Y(n1790) );
  BUFX2 U1206 ( .A(n1174), .Y(n1791) );
  BUFX2 U1207 ( .A(n1176), .Y(n1793) );
  BUFX2 U1208 ( .A(n1176), .Y(n1794) );
  BUFX2 U1209 ( .A(n1178), .Y(n1796) );
  BUFX2 U1210 ( .A(n1178), .Y(n1797) );
  BUFX2 U1211 ( .A(n1180), .Y(n1799) );
  BUFX2 U1212 ( .A(n1180), .Y(n1800) );
  BUFX2 U1213 ( .A(n1182), .Y(n1802) );
  BUFX2 U1214 ( .A(n1182), .Y(n1803) );
  BUFX2 U1215 ( .A(n1184), .Y(n1805) );
  BUFX2 U1216 ( .A(n1184), .Y(n1806) );
  BUFX2 U1217 ( .A(n1186), .Y(n1808) );
  BUFX2 U1218 ( .A(n1186), .Y(n1809) );
  BUFX2 U1219 ( .A(n1188), .Y(n1811) );
  BUFX2 U1220 ( .A(n1188), .Y(n1812) );
  BUFX2 U1221 ( .A(n1190), .Y(n1814) );
  BUFX2 U1222 ( .A(n1190), .Y(n1815) );
  BUFX2 U1223 ( .A(n1192), .Y(n1817) );
  BUFX2 U1224 ( .A(n1192), .Y(n1818) );
  BUFX2 U1225 ( .A(n1194), .Y(n1820) );
  BUFX2 U1226 ( .A(n1194), .Y(n1821) );
  BUFX2 U1227 ( .A(n1196), .Y(n1823) );
  BUFX2 U1228 ( .A(n1196), .Y(n1824) );
  BUFX2 U1229 ( .A(n1198), .Y(n1826) );
  BUFX2 U1230 ( .A(n1198), .Y(n1827) );
  INVX1 U1231 ( .A(n1871), .Y(n1870) );
  AND2X1 U1232 ( .A(\data_in<7> ), .B(n1830), .Y(n60) );
  AND2X1 U1233 ( .A(\data_in<6> ), .B(n1830), .Y(n62) );
  AND2X1 U1234 ( .A(\data_in<5> ), .B(n1830), .Y(n64) );
  AND2X1 U1235 ( .A(\data_in<4> ), .B(n1830), .Y(n66) );
  AND2X1 U1236 ( .A(\data_in<3> ), .B(n1830), .Y(n68) );
  AND2X1 U1237 ( .A(\data_in<2> ), .B(n1830), .Y(n70) );
  AND2X1 U1238 ( .A(\data_in<1> ), .B(n1830), .Y(n72) );
  AND2X1 U1239 ( .A(\data_in<0> ), .B(n1830), .Y(n74) );
  BUFX2 U1240 ( .A(n2390), .Y(n76) );
  INVX1 U1241 ( .A(n76), .Y(n1874) );
  BUFX2 U1242 ( .A(n2519), .Y(n80) );
  INVX1 U1243 ( .A(n80), .Y(n1877) );
  BUFX2 U1244 ( .A(n2648), .Y(n82) );
  INVX1 U1245 ( .A(n82), .Y(n1875) );
  BUFX2 U1246 ( .A(n2778), .Y(n99) );
  INVX1 U1247 ( .A(n99), .Y(n1876) );
  AND2X1 U1248 ( .A(n1874), .B(n2779), .Y(n101) );
  INVX1 U1249 ( .A(n60), .Y(n1842) );
  INVX2 U1250 ( .A(n60), .Y(n1841) );
  INVX2 U1251 ( .A(n60), .Y(n1840) );
  INVX1 U1252 ( .A(n62), .Y(n1845) );
  INVX2 U1253 ( .A(n62), .Y(n1844) );
  INVX2 U1254 ( .A(n62), .Y(n1843) );
  INVX1 U1255 ( .A(n64), .Y(n1848) );
  INVX2 U1256 ( .A(n64), .Y(n1847) );
  INVX2 U1257 ( .A(n64), .Y(n1846) );
  INVX1 U1258 ( .A(n66), .Y(n1851) );
  INVX2 U1259 ( .A(n66), .Y(n1850) );
  INVX2 U1260 ( .A(n66), .Y(n1849) );
  INVX1 U1261 ( .A(n68), .Y(n1854) );
  INVX2 U1262 ( .A(n68), .Y(n1853) );
  INVX2 U1263 ( .A(n68), .Y(n1852) );
  INVX1 U1264 ( .A(n70), .Y(n1857) );
  INVX2 U1265 ( .A(n70), .Y(n1856) );
  INVX2 U1266 ( .A(n70), .Y(n1855) );
  INVX1 U1267 ( .A(n72), .Y(n1860) );
  INVX2 U1268 ( .A(n72), .Y(n1859) );
  INVX2 U1269 ( .A(n72), .Y(n1858) );
  INVX1 U1270 ( .A(n74), .Y(n1863) );
  INVX2 U1271 ( .A(n74), .Y(n1862) );
  INVX2 U1272 ( .A(n74), .Y(n1861) );
  AND2X1 U1273 ( .A(n1874), .B(n2796), .Y(n118) );
  AND2X1 U1274 ( .A(n1874), .B(n2813), .Y(n120) );
  AND2X1 U1275 ( .A(n1874), .B(n2830), .Y(n137) );
  AND2X1 U1276 ( .A(n1874), .B(n2847), .Y(n139) );
  AND2X1 U1277 ( .A(n1874), .B(n2864), .Y(n156) );
  AND2X1 U1278 ( .A(n1874), .B(n2881), .Y(n158) );
  AND2X1 U1279 ( .A(n1874), .B(n2898), .Y(n175) );
  AND2X1 U1280 ( .A(n1877), .B(n2779), .Y(n177) );
  AND2X1 U1281 ( .A(n1877), .B(n2796), .Y(n194) );
  AND2X1 U1282 ( .A(n1877), .B(n2813), .Y(n196) );
  AND2X1 U1283 ( .A(n1877), .B(n2830), .Y(n215) );
  AND2X1 U1284 ( .A(n1877), .B(n2847), .Y(n217) );
  AND2X1 U1285 ( .A(n1877), .B(n2864), .Y(n233) );
  AND2X1 U1286 ( .A(n1877), .B(n2881), .Y(n235) );
  AND2X1 U1287 ( .A(n1877), .B(n2898), .Y(n251) );
  AND2X1 U1288 ( .A(n1875), .B(n2779), .Y(n253) );
  AND2X1 U1289 ( .A(n1875), .B(n2796), .Y(n269) );
  AND2X1 U1290 ( .A(n1875), .B(n2813), .Y(n271) );
  AND2X1 U1291 ( .A(n1875), .B(n2830), .Y(n287) );
  AND2X1 U1292 ( .A(n1875), .B(n2847), .Y(n289) );
  AND2X1 U1293 ( .A(n1875), .B(n2864), .Y(n305) );
  AND2X1 U1294 ( .A(n1875), .B(n2881), .Y(n307) );
  AND2X1 U1295 ( .A(n1875), .B(n2898), .Y(n323) );
  AND2X1 U1296 ( .A(n2779), .B(n1876), .Y(n325) );
  AND2X1 U1297 ( .A(n2796), .B(n1876), .Y(n341) );
  AND2X1 U1298 ( .A(n2813), .B(n1876), .Y(n343) );
  AND2X1 U1299 ( .A(n2830), .B(n1876), .Y(n360) );
  AND2X1 U1300 ( .A(n2847), .B(n1876), .Y(n362) );
  AND2X1 U1301 ( .A(n2864), .B(n1876), .Y(n378) );
  AND2X1 U1302 ( .A(n2881), .B(n1876), .Y(n380) );
  AND2X1 U1303 ( .A(n2898), .B(n1876), .Y(n396) );
  AND2X2 U1304 ( .A(n101), .B(n1829), .Y(n398) );
  INVX1 U1305 ( .A(n398), .Y(n414) );
  AND2X2 U1306 ( .A(n118), .B(n1830), .Y(n416) );
  INVX1 U1307 ( .A(n416), .Y(n432) );
  AND2X2 U1308 ( .A(n120), .B(n1830), .Y(n434) );
  INVX1 U1309 ( .A(n434), .Y(n450) );
  AND2X2 U1310 ( .A(n137), .B(n1830), .Y(n452) );
  INVX1 U1311 ( .A(n452), .Y(n468) );
  AND2X2 U1312 ( .A(n139), .B(n1830), .Y(n470) );
  INVX1 U1313 ( .A(n470), .Y(n486) );
  AND2X2 U1314 ( .A(n156), .B(n1830), .Y(n488) );
  INVX1 U1315 ( .A(n488), .Y(n505) );
  AND2X2 U1316 ( .A(n158), .B(n1829), .Y(n507) );
  INVX1 U1317 ( .A(n507), .Y(n523) );
  AND2X2 U1318 ( .A(n175), .B(n1829), .Y(n525) );
  INVX1 U1319 ( .A(n525), .Y(n541) );
  AND2X2 U1320 ( .A(n177), .B(n1829), .Y(n543) );
  INVX1 U1321 ( .A(n543), .Y(n559) );
  AND2X2 U1322 ( .A(n194), .B(n1829), .Y(n561) );
  INVX1 U1323 ( .A(n561), .Y(n577) );
  AND2X2 U1324 ( .A(n196), .B(n1829), .Y(n579) );
  INVX1 U1325 ( .A(n579), .Y(n595) );
  AND2X2 U1326 ( .A(n215), .B(n1829), .Y(n597) );
  INVX1 U1327 ( .A(n597), .Y(n613) );
  AND2X2 U1328 ( .A(n217), .B(n1829), .Y(n615) );
  INVX1 U1329 ( .A(n615), .Y(n631) );
  AND2X2 U1330 ( .A(n233), .B(n1829), .Y(n633) );
  INVX1 U1331 ( .A(n633), .Y(n650) );
  AND2X2 U1332 ( .A(n235), .B(n1829), .Y(n1163) );
  INVX1 U1333 ( .A(n1163), .Y(n1164) );
  AND2X2 U1334 ( .A(n251), .B(n1829), .Y(n1165) );
  INVX1 U1335 ( .A(n1165), .Y(n1166) );
  AND2X2 U1336 ( .A(n253), .B(n1829), .Y(n1167) );
  INVX1 U1337 ( .A(n1167), .Y(n1168) );
  AND2X2 U1338 ( .A(n269), .B(n1829), .Y(n1169) );
  INVX1 U1339 ( .A(n1169), .Y(n1170) );
  AND2X2 U1340 ( .A(n271), .B(n1829), .Y(n1171) );
  INVX1 U1341 ( .A(n1171), .Y(n1172) );
  AND2X1 U1342 ( .A(n287), .B(n1828), .Y(n1173) );
  INVX1 U1343 ( .A(n1173), .Y(n1174) );
  AND2X1 U1344 ( .A(n289), .B(n1828), .Y(n1175) );
  INVX1 U1345 ( .A(n1175), .Y(n1176) );
  AND2X1 U1346 ( .A(n305), .B(n1828), .Y(n1177) );
  INVX1 U1347 ( .A(n1177), .Y(n1178) );
  AND2X1 U1348 ( .A(n307), .B(n1828), .Y(n1179) );
  INVX1 U1349 ( .A(n1179), .Y(n1180) );
  AND2X1 U1350 ( .A(n323), .B(n1828), .Y(n1181) );
  INVX1 U1351 ( .A(n1181), .Y(n1182) );
  AND2X1 U1352 ( .A(n325), .B(n1828), .Y(n1183) );
  INVX1 U1353 ( .A(n1183), .Y(n1184) );
  AND2X1 U1354 ( .A(n341), .B(n1828), .Y(n1185) );
  INVX1 U1355 ( .A(n1185), .Y(n1186) );
  AND2X1 U1356 ( .A(n343), .B(n1828), .Y(n1187) );
  INVX1 U1357 ( .A(n1187), .Y(n1188) );
  AND2X1 U1358 ( .A(n360), .B(n1828), .Y(n1189) );
  INVX1 U1359 ( .A(n1189), .Y(n1190) );
  AND2X1 U1360 ( .A(n362), .B(n1828), .Y(n1191) );
  INVX1 U1361 ( .A(n1191), .Y(n1192) );
  AND2X1 U1362 ( .A(n378), .B(n1828), .Y(n1193) );
  INVX1 U1363 ( .A(n1193), .Y(n1194) );
  AND2X1 U1364 ( .A(n380), .B(n1828), .Y(n1195) );
  INVX1 U1365 ( .A(n1195), .Y(n1196) );
  AND2X1 U1366 ( .A(n396), .B(n1828), .Y(n1197) );
  INVX1 U1367 ( .A(n1197), .Y(n1198) );
  MUX2X1 U1368 ( .B(n1200), .A(n1201), .S(n1707), .Y(n1199) );
  MUX2X1 U1369 ( .B(n1203), .A(n1204), .S(n1707), .Y(n1202) );
  MUX2X1 U1370 ( .B(n1206), .A(n1207), .S(n1707), .Y(n1205) );
  MUX2X1 U1371 ( .B(n1209), .A(n1210), .S(n1707), .Y(n1208) );
  MUX2X1 U1372 ( .B(n1212), .A(n1213), .S(n1697), .Y(n1211) );
  MUX2X1 U1373 ( .B(n1215), .A(n1216), .S(n1707), .Y(n1214) );
  MUX2X1 U1374 ( .B(n1218), .A(n1219), .S(n1707), .Y(n1217) );
  MUX2X1 U1375 ( .B(n1221), .A(n1222), .S(n1707), .Y(n1220) );
  MUX2X1 U1376 ( .B(n1224), .A(n1225), .S(n1707), .Y(n1223) );
  MUX2X1 U1377 ( .B(n1227), .A(n1228), .S(n1697), .Y(n1226) );
  MUX2X1 U1378 ( .B(n1230), .A(n1231), .S(n1708), .Y(n1229) );
  MUX2X1 U1379 ( .B(n1233), .A(n1234), .S(n1708), .Y(n1232) );
  MUX2X1 U1380 ( .B(n1236), .A(n1237), .S(n1708), .Y(n1235) );
  MUX2X1 U1381 ( .B(n1239), .A(n1240), .S(n1708), .Y(n1238) );
  MUX2X1 U1382 ( .B(n1242), .A(n1243), .S(n1697), .Y(n1241) );
  MUX2X1 U1383 ( .B(n1245), .A(n1246), .S(n1708), .Y(n1244) );
  MUX2X1 U1384 ( .B(n1248), .A(n1249), .S(n1708), .Y(n1247) );
  MUX2X1 U1385 ( .B(n1251), .A(n1252), .S(n1708), .Y(n1250) );
  MUX2X1 U1386 ( .B(n1254), .A(n1255), .S(n1708), .Y(n1253) );
  MUX2X1 U1387 ( .B(n1257), .A(n1258), .S(n1697), .Y(n1256) );
  MUX2X1 U1388 ( .B(n1260), .A(n1261), .S(n1708), .Y(n1259) );
  MUX2X1 U1389 ( .B(n1263), .A(n1264), .S(n1708), .Y(n1262) );
  MUX2X1 U1390 ( .B(n1266), .A(n1267), .S(n1708), .Y(n1265) );
  MUX2X1 U1391 ( .B(n1269), .A(n1270), .S(n1708), .Y(n1268) );
  MUX2X1 U1392 ( .B(n1272), .A(n1273), .S(n1697), .Y(n1271) );
  MUX2X1 U1393 ( .B(n1275), .A(n1276), .S(n1709), .Y(n1274) );
  MUX2X1 U1394 ( .B(n1278), .A(n1279), .S(n1709), .Y(n1277) );
  MUX2X1 U1395 ( .B(n1281), .A(n1282), .S(n1709), .Y(n1280) );
  MUX2X1 U1396 ( .B(n1284), .A(n1285), .S(n1709), .Y(n1283) );
  MUX2X1 U1397 ( .B(n1287), .A(n1288), .S(n1697), .Y(n1286) );
  MUX2X1 U1398 ( .B(n1290), .A(n1291), .S(n1709), .Y(n1289) );
  MUX2X1 U1399 ( .B(n1293), .A(n1294), .S(n1709), .Y(n1292) );
  MUX2X1 U1400 ( .B(n1296), .A(n1297), .S(n1709), .Y(n1295) );
  MUX2X1 U1401 ( .B(n1299), .A(n1300), .S(n1709), .Y(n1298) );
  MUX2X1 U1402 ( .B(n1302), .A(n1303), .S(n1697), .Y(n1301) );
  MUX2X1 U1403 ( .B(n1305), .A(n1306), .S(n1709), .Y(n1304) );
  MUX2X1 U1404 ( .B(n1308), .A(n1309), .S(n1709), .Y(n1307) );
  MUX2X1 U1405 ( .B(n1311), .A(n1312), .S(n1709), .Y(n1310) );
  MUX2X1 U1406 ( .B(n1314), .A(n1315), .S(n1709), .Y(n1313) );
  MUX2X1 U1407 ( .B(n1317), .A(n1318), .S(n1697), .Y(n1316) );
  MUX2X1 U1408 ( .B(n1320), .A(n1321), .S(n1710), .Y(n1319) );
  MUX2X1 U1409 ( .B(n1323), .A(n1324), .S(n1710), .Y(n1322) );
  MUX2X1 U1410 ( .B(n1326), .A(n1327), .S(n1710), .Y(n1325) );
  MUX2X1 U1411 ( .B(n1329), .A(n1330), .S(n1710), .Y(n1328) );
  MUX2X1 U1412 ( .B(n1332), .A(n1333), .S(n1697), .Y(n1331) );
  MUX2X1 U1413 ( .B(n1335), .A(n1336), .S(n1710), .Y(n1334) );
  MUX2X1 U1414 ( .B(n1338), .A(n1339), .S(n1710), .Y(n1337) );
  MUX2X1 U1415 ( .B(n1341), .A(n1342), .S(n1710), .Y(n1340) );
  MUX2X1 U1416 ( .B(n1344), .A(n1345), .S(n1710), .Y(n1343) );
  MUX2X1 U1417 ( .B(n1347), .A(n1348), .S(n1697), .Y(n1346) );
  MUX2X1 U1418 ( .B(n1350), .A(n1351), .S(n1710), .Y(n1349) );
  MUX2X1 U1419 ( .B(n1353), .A(n1354), .S(n1710), .Y(n1352) );
  MUX2X1 U1420 ( .B(n1356), .A(n1357), .S(n1710), .Y(n1355) );
  MUX2X1 U1421 ( .B(n1359), .A(n1360), .S(n1710), .Y(n1358) );
  MUX2X1 U1422 ( .B(n1362), .A(n1363), .S(n1697), .Y(n1361) );
  MUX2X1 U1423 ( .B(n1365), .A(n1366), .S(n1711), .Y(n1364) );
  MUX2X1 U1424 ( .B(n1368), .A(n1369), .S(n1711), .Y(n1367) );
  MUX2X1 U1425 ( .B(n1371), .A(n1372), .S(n1711), .Y(n1370) );
  MUX2X1 U1426 ( .B(n1374), .A(n1375), .S(n1711), .Y(n1373) );
  MUX2X1 U1427 ( .B(n1377), .A(n1378), .S(n1697), .Y(n1376) );
  MUX2X1 U1428 ( .B(n1380), .A(n1381), .S(n1711), .Y(n1379) );
  MUX2X1 U1429 ( .B(n1383), .A(n1384), .S(n1711), .Y(n1382) );
  MUX2X1 U1430 ( .B(n1386), .A(n1387), .S(n1711), .Y(n1385) );
  MUX2X1 U1431 ( .B(n1389), .A(n1390), .S(n1711), .Y(n1388) );
  MUX2X1 U1432 ( .B(n1392), .A(n1393), .S(n1696), .Y(n1391) );
  MUX2X1 U1433 ( .B(n1395), .A(n1396), .S(n1711), .Y(n1394) );
  MUX2X1 U1434 ( .B(n1398), .A(n1399), .S(n1711), .Y(n1397) );
  MUX2X1 U1435 ( .B(n1401), .A(n1402), .S(n1711), .Y(n1400) );
  MUX2X1 U1436 ( .B(n1404), .A(n1405), .S(n1711), .Y(n1403) );
  MUX2X1 U1437 ( .B(n1407), .A(n1408), .S(n1696), .Y(n1406) );
  MUX2X1 U1438 ( .B(n1410), .A(n1411), .S(n1710), .Y(n1409) );
  MUX2X1 U1439 ( .B(n1413), .A(n1414), .S(n1711), .Y(n1412) );
  MUX2X1 U1440 ( .B(n1416), .A(n1417), .S(n1711), .Y(n1415) );
  MUX2X1 U1441 ( .B(n1419), .A(n1420), .S(n1710), .Y(n1418) );
  MUX2X1 U1442 ( .B(n1422), .A(n1423), .S(n1696), .Y(n1421) );
  MUX2X1 U1443 ( .B(n1425), .A(n1426), .S(n1710), .Y(n1424) );
  MUX2X1 U1444 ( .B(n1428), .A(n1429), .S(n1710), .Y(n1427) );
  MUX2X1 U1445 ( .B(n1431), .A(n1432), .S(n1711), .Y(n1430) );
  MUX2X1 U1446 ( .B(n1434), .A(n1435), .S(n1710), .Y(n1433) );
  MUX2X1 U1447 ( .B(n1437), .A(n1438), .S(n1696), .Y(n1436) );
  MUX2X1 U1448 ( .B(n1440), .A(n1441), .S(n1711), .Y(n1439) );
  MUX2X1 U1449 ( .B(n1443), .A(n1444), .S(n1710), .Y(n1442) );
  MUX2X1 U1450 ( .B(n1446), .A(n1447), .S(n1710), .Y(n1445) );
  MUX2X1 U1451 ( .B(n1449), .A(n1450), .S(n1710), .Y(n1448) );
  MUX2X1 U1452 ( .B(n1452), .A(n1453), .S(n1696), .Y(n1451) );
  MUX2X1 U1453 ( .B(n1455), .A(n1456), .S(n1712), .Y(n1454) );
  MUX2X1 U1454 ( .B(n1458), .A(n1459), .S(n1712), .Y(n1457) );
  MUX2X1 U1455 ( .B(n1461), .A(n1462), .S(n1712), .Y(n1460) );
  MUX2X1 U1456 ( .B(n1464), .A(n1465), .S(n1712), .Y(n1463) );
  MUX2X1 U1457 ( .B(n1467), .A(n1468), .S(n1696), .Y(n1466) );
  MUX2X1 U1458 ( .B(n1470), .A(n1471), .S(n1712), .Y(n1469) );
  MUX2X1 U1459 ( .B(n1473), .A(n1474), .S(n1712), .Y(n1472) );
  MUX2X1 U1460 ( .B(n1476), .A(n1477), .S(n1712), .Y(n1475) );
  MUX2X1 U1461 ( .B(n1479), .A(n1480), .S(n1712), .Y(n1478) );
  MUX2X1 U1462 ( .B(n1482), .A(n1483), .S(n1696), .Y(n1481) );
  MUX2X1 U1463 ( .B(n1485), .A(n1486), .S(n1712), .Y(n1484) );
  MUX2X1 U1464 ( .B(n1488), .A(n1489), .S(n1712), .Y(n1487) );
  MUX2X1 U1465 ( .B(n1491), .A(n1492), .S(n1712), .Y(n1490) );
  MUX2X1 U1466 ( .B(n1494), .A(n1495), .S(n1712), .Y(n1493) );
  MUX2X1 U1467 ( .B(n1497), .A(n1498), .S(n1696), .Y(n1496) );
  MUX2X1 U1468 ( .B(n1500), .A(n1501), .S(n1713), .Y(n1499) );
  MUX2X1 U1469 ( .B(n1503), .A(n1504), .S(n1713), .Y(n1502) );
  MUX2X1 U1470 ( .B(n1506), .A(n1507), .S(n1713), .Y(n1505) );
  MUX2X1 U1471 ( .B(n1509), .A(n1510), .S(n1713), .Y(n1508) );
  MUX2X1 U1472 ( .B(n1512), .A(n1513), .S(n1696), .Y(n1511) );
  MUX2X1 U1473 ( .B(n1515), .A(n1516), .S(n1713), .Y(n1514) );
  MUX2X1 U1474 ( .B(n1518), .A(n1519), .S(n1713), .Y(n1517) );
  MUX2X1 U1475 ( .B(n1521), .A(n1522), .S(n1713), .Y(n1520) );
  MUX2X1 U1476 ( .B(n1524), .A(n1525), .S(n1713), .Y(n1523) );
  MUX2X1 U1477 ( .B(n1527), .A(n1528), .S(n1696), .Y(n1526) );
  MUX2X1 U1478 ( .B(n1530), .A(n1531), .S(n1713), .Y(n1529) );
  MUX2X1 U1479 ( .B(n1533), .A(n1534), .S(n1713), .Y(n1532) );
  MUX2X1 U1480 ( .B(n1536), .A(n1537), .S(n1713), .Y(n1535) );
  MUX2X1 U1481 ( .B(n1539), .A(n1540), .S(n1713), .Y(n1538) );
  MUX2X1 U1482 ( .B(n1542), .A(n1543), .S(n1696), .Y(n1541) );
  MUX2X1 U1483 ( .B(n1545), .A(n1546), .S(n1714), .Y(n1544) );
  MUX2X1 U1484 ( .B(n1548), .A(n1549), .S(n1714), .Y(n1547) );
  MUX2X1 U1485 ( .B(n1551), .A(n1552), .S(n1714), .Y(n1550) );
  MUX2X1 U1486 ( .B(n1554), .A(n1555), .S(n1714), .Y(n1553) );
  MUX2X1 U1487 ( .B(n1557), .A(n1558), .S(n1696), .Y(n1556) );
  MUX2X1 U1488 ( .B(n1560), .A(n1561), .S(n1714), .Y(n1559) );
  MUX2X1 U1489 ( .B(n1563), .A(n1564), .S(n1714), .Y(n1562) );
  MUX2X1 U1490 ( .B(n1566), .A(n1567), .S(n1714), .Y(n1565) );
  MUX2X1 U1491 ( .B(n1569), .A(n1570), .S(n1714), .Y(n1568) );
  MUX2X1 U1492 ( .B(n1572), .A(n1573), .S(n1697), .Y(n1571) );
  MUX2X1 U1493 ( .B(n1575), .A(n1576), .S(n1714), .Y(n1574) );
  MUX2X1 U1494 ( .B(n1578), .A(n1579), .S(n1714), .Y(n1577) );
  MUX2X1 U1495 ( .B(n1581), .A(n1582), .S(n1714), .Y(n1580) );
  MUX2X1 U1496 ( .B(n1584), .A(n1585), .S(n1714), .Y(n1583) );
  MUX2X1 U1497 ( .B(n1587), .A(n1588), .S(n1697), .Y(n1586) );
  MUX2X1 U1498 ( .B(n1590), .A(n1591), .S(n1715), .Y(n1589) );
  MUX2X1 U1499 ( .B(n1593), .A(n1594), .S(n1715), .Y(n1592) );
  MUX2X1 U1500 ( .B(n1596), .A(n1597), .S(n1715), .Y(n1595) );
  MUX2X1 U1501 ( .B(n1599), .A(n1600), .S(n1715), .Y(n1598) );
  MUX2X1 U1502 ( .B(n1602), .A(n1603), .S(n1697), .Y(n1601) );
  MUX2X1 U1503 ( .B(n1605), .A(n1606), .S(n1715), .Y(n1604) );
  MUX2X1 U1504 ( .B(n1608), .A(n1609), .S(n1715), .Y(n1607) );
  MUX2X1 U1505 ( .B(n1611), .A(n1612), .S(n1715), .Y(n1610) );
  MUX2X1 U1506 ( .B(n1614), .A(n1615), .S(n1715), .Y(n1613) );
  MUX2X1 U1507 ( .B(n1617), .A(n1618), .S(n1697), .Y(n1616) );
  MUX2X1 U1508 ( .B(n1620), .A(n1621), .S(n1715), .Y(n1619) );
  MUX2X1 U1509 ( .B(n1623), .A(n1624), .S(n1715), .Y(n1622) );
  MUX2X1 U1510 ( .B(n1626), .A(n1627), .S(n1715), .Y(n1625) );
  MUX2X1 U1511 ( .B(n1629), .A(n1630), .S(n1715), .Y(n1628) );
  MUX2X1 U1512 ( .B(n1632), .A(n1633), .S(n1696), .Y(n1631) );
  MUX2X1 U1513 ( .B(n1635), .A(n1636), .S(n1716), .Y(n1634) );
  MUX2X1 U1514 ( .B(n1638), .A(n1639), .S(n1716), .Y(n1637) );
  MUX2X1 U1515 ( .B(n1641), .A(n1642), .S(n1716), .Y(n1640) );
  MUX2X1 U1516 ( .B(n1644), .A(n1645), .S(n1716), .Y(n1643) );
  MUX2X1 U1517 ( .B(n1647), .A(n1648), .S(n1696), .Y(n1646) );
  MUX2X1 U1518 ( .B(n1650), .A(n1651), .S(n1716), .Y(n1649) );
  MUX2X1 U1519 ( .B(n1653), .A(n1654), .S(n1716), .Y(n1652) );
  MUX2X1 U1520 ( .B(n1656), .A(n1657), .S(n1716), .Y(n1655) );
  MUX2X1 U1521 ( .B(n1659), .A(n1660), .S(n1716), .Y(n1658) );
  MUX2X1 U1522 ( .B(n1662), .A(n1663), .S(n1696), .Y(n1661) );
  MUX2X1 U1523 ( .B(n1665), .A(n1666), .S(n1716), .Y(n1664) );
  MUX2X1 U1524 ( .B(n1668), .A(n1669), .S(n1716), .Y(n1667) );
  MUX2X1 U1525 ( .B(n1671), .A(n1672), .S(n1716), .Y(n1670) );
  MUX2X1 U1526 ( .B(n1674), .A(n1675), .S(n1716), .Y(n1673) );
  MUX2X1 U1527 ( .B(n1677), .A(n1678), .S(n1696), .Y(n1676) );
  MUX2X1 U1528 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1729), .Y(n1201) );
  MUX2X1 U1529 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1727), .Y(n1200) );
  MUX2X1 U1530 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1721), .Y(n1204) );
  MUX2X1 U1531 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1719), .Y(n1203) );
  MUX2X1 U1532 ( .B(n1202), .A(n1199), .S(n1703), .Y(n1213) );
  MUX2X1 U1533 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1719), .Y(n1207) );
  MUX2X1 U1534 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1719), .Y(n1206) );
  MUX2X1 U1535 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1719), .Y(n1210) );
  MUX2X1 U1536 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1719), .Y(n1209) );
  MUX2X1 U1537 ( .B(n1208), .A(n1205), .S(n1703), .Y(n1212) );
  MUX2X1 U1538 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1719), .Y(n1216) );
  MUX2X1 U1539 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1719), .Y(n1215) );
  MUX2X1 U1540 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1719), .Y(n1219) );
  MUX2X1 U1541 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1719), .Y(n1218) );
  MUX2X1 U1542 ( .B(n1217), .A(n1214), .S(n1703), .Y(n1228) );
  MUX2X1 U1543 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1719), .Y(n1222) );
  MUX2X1 U1544 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1719), .Y(n1221) );
  MUX2X1 U1545 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1719), .Y(n1225) );
  MUX2X1 U1546 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1719), .Y(n1224) );
  MUX2X1 U1547 ( .B(n1223), .A(n1220), .S(n1703), .Y(n1227) );
  MUX2X1 U1548 ( .B(n1226), .A(n1211), .S(n1695), .Y(n1679) );
  MUX2X1 U1549 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1720), .Y(n1231) );
  MUX2X1 U1550 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1720), .Y(n1230) );
  MUX2X1 U1551 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1720), .Y(n1234) );
  MUX2X1 U1552 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1720), .Y(n1233) );
  MUX2X1 U1553 ( .B(n1232), .A(n1229), .S(n1703), .Y(n1243) );
  MUX2X1 U1554 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1720), .Y(n1237) );
  MUX2X1 U1555 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1720), .Y(n1236) );
  MUX2X1 U1556 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1720), .Y(n1240) );
  MUX2X1 U1557 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1720), .Y(n1239) );
  MUX2X1 U1558 ( .B(n1238), .A(n1235), .S(n1703), .Y(n1242) );
  MUX2X1 U1559 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1720), .Y(n1246) );
  MUX2X1 U1560 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1720), .Y(n1245) );
  MUX2X1 U1561 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1720), .Y(n1249) );
  MUX2X1 U1562 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1720), .Y(n1248) );
  MUX2X1 U1563 ( .B(n1247), .A(n1244), .S(n1703), .Y(n1258) );
  MUX2X1 U1564 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1721), .Y(n1252) );
  MUX2X1 U1565 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1721), .Y(n1251) );
  MUX2X1 U1566 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1721), .Y(n1255) );
  MUX2X1 U1567 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1721), .Y(n1254) );
  MUX2X1 U1568 ( .B(n1253), .A(n1250), .S(n1703), .Y(n1257) );
  MUX2X1 U1569 ( .B(n1256), .A(n1241), .S(n1695), .Y(n1680) );
  MUX2X1 U1570 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1721), .Y(n1261) );
  MUX2X1 U1571 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1721), .Y(n1260) );
  MUX2X1 U1572 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1721), .Y(n1264) );
  MUX2X1 U1573 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1721), .Y(n1263) );
  MUX2X1 U1574 ( .B(n1262), .A(n1259), .S(n1703), .Y(n1273) );
  MUX2X1 U1575 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1721), .Y(n1267) );
  MUX2X1 U1576 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1721), .Y(n1266) );
  MUX2X1 U1577 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1721), .Y(n1270) );
  MUX2X1 U1578 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1721), .Y(n1269) );
  MUX2X1 U1579 ( .B(n1268), .A(n1265), .S(n1703), .Y(n1272) );
  MUX2X1 U1580 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1722), .Y(n1276) );
  MUX2X1 U1581 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1722), .Y(n1275) );
  MUX2X1 U1582 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1722), .Y(n1279) );
  MUX2X1 U1583 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1722), .Y(n1278) );
  MUX2X1 U1584 ( .B(n1277), .A(n1274), .S(n1703), .Y(n1288) );
  MUX2X1 U1585 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1722), .Y(n1282) );
  MUX2X1 U1586 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1722), .Y(n1281) );
  MUX2X1 U1587 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1722), .Y(n1285) );
  MUX2X1 U1588 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1722), .Y(n1284) );
  MUX2X1 U1589 ( .B(n1283), .A(n1280), .S(n1703), .Y(n1287) );
  MUX2X1 U1590 ( .B(n1286), .A(n1271), .S(n1695), .Y(n1681) );
  MUX2X1 U1591 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1722), .Y(n1291) );
  MUX2X1 U1592 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1722), .Y(n1290) );
  MUX2X1 U1593 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1722), .Y(n1294) );
  MUX2X1 U1594 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1722), .Y(n1293) );
  MUX2X1 U1595 ( .B(n1292), .A(n1289), .S(n1702), .Y(n1303) );
  MUX2X1 U1596 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1720), .Y(n1297) );
  MUX2X1 U1597 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1719), .Y(n1296) );
  MUX2X1 U1598 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1720), .Y(n1300) );
  MUX2X1 U1599 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1719), .Y(n1299) );
  MUX2X1 U1600 ( .B(n1298), .A(n1295), .S(n1702), .Y(n1302) );
  MUX2X1 U1601 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1720), .Y(n1306) );
  MUX2X1 U1602 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1720), .Y(n1305) );
  MUX2X1 U1603 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1720), .Y(n1309) );
  MUX2X1 U1604 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1720), .Y(n1308) );
  MUX2X1 U1605 ( .B(n1307), .A(n1304), .S(n1702), .Y(n1318) );
  MUX2X1 U1606 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1719), .Y(n1312) );
  MUX2X1 U1607 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1721), .Y(n1311) );
  MUX2X1 U1608 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1720), .Y(n1315) );
  MUX2X1 U1609 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1720), .Y(n1314) );
  MUX2X1 U1610 ( .B(n1313), .A(n1310), .S(n1702), .Y(n1317) );
  MUX2X1 U1611 ( .B(n1316), .A(n1301), .S(n1695), .Y(n1682) );
  MUX2X1 U1612 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1723), .Y(n1321) );
  MUX2X1 U1613 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1723), .Y(n1320) );
  MUX2X1 U1614 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1723), .Y(n1324) );
  MUX2X1 U1615 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1723), .Y(n1323) );
  MUX2X1 U1616 ( .B(n1322), .A(n1319), .S(n1702), .Y(n1333) );
  MUX2X1 U1617 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1723), .Y(n1327) );
  MUX2X1 U1618 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1723), .Y(n1326) );
  MUX2X1 U1619 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1723), .Y(n1330) );
  MUX2X1 U1620 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1723), .Y(n1329) );
  MUX2X1 U1621 ( .B(n1328), .A(n1325), .S(n1702), .Y(n1332) );
  MUX2X1 U1622 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1723), .Y(n1336) );
  MUX2X1 U1623 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1723), .Y(n1335) );
  MUX2X1 U1624 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1723), .Y(n1339) );
  MUX2X1 U1625 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1723), .Y(n1338) );
  MUX2X1 U1626 ( .B(n1337), .A(n1334), .S(n1702), .Y(n1348) );
  MUX2X1 U1627 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1724), .Y(n1342) );
  MUX2X1 U1628 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1724), .Y(n1341) );
  MUX2X1 U1629 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1724), .Y(n1345) );
  MUX2X1 U1630 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1724), .Y(n1344) );
  MUX2X1 U1631 ( .B(n1343), .A(n1340), .S(n1702), .Y(n1347) );
  MUX2X1 U1632 ( .B(n1346), .A(n1331), .S(n1695), .Y(n1683) );
  MUX2X1 U1633 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1724), .Y(n1351) );
  MUX2X1 U1634 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1724), .Y(n1350) );
  MUX2X1 U1635 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1724), .Y(n1354) );
  MUX2X1 U1636 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1724), .Y(n1353) );
  MUX2X1 U1637 ( .B(n1352), .A(n1349), .S(n1702), .Y(n1363) );
  MUX2X1 U1638 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1724), .Y(n1357) );
  MUX2X1 U1639 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1724), .Y(n1356) );
  MUX2X1 U1640 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1724), .Y(n1360) );
  MUX2X1 U1641 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1724), .Y(n1359) );
  MUX2X1 U1642 ( .B(n1358), .A(n1355), .S(n1702), .Y(n1362) );
  MUX2X1 U1643 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1725), .Y(n1366) );
  MUX2X1 U1644 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1725), .Y(n1365) );
  MUX2X1 U1645 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1725), .Y(n1369) );
  MUX2X1 U1646 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1725), .Y(n1368) );
  MUX2X1 U1647 ( .B(n1367), .A(n1364), .S(n1702), .Y(n1378) );
  MUX2X1 U1648 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1725), .Y(n1372) );
  MUX2X1 U1649 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1725), .Y(n1371) );
  MUX2X1 U1650 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1725), .Y(n1375) );
  MUX2X1 U1651 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1725), .Y(n1374) );
  MUX2X1 U1652 ( .B(n1373), .A(n1370), .S(n1702), .Y(n1377) );
  MUX2X1 U1653 ( .B(n1376), .A(n1361), .S(n1695), .Y(n1684) );
  MUX2X1 U1654 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1725), .Y(n1381) );
  MUX2X1 U1655 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1725), .Y(n1380) );
  MUX2X1 U1656 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1725), .Y(n1384) );
  MUX2X1 U1657 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1725), .Y(n1383) );
  MUX2X1 U1658 ( .B(n1382), .A(n1379), .S(n1702), .Y(n1393) );
  MUX2X1 U1659 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1726), .Y(n1387) );
  MUX2X1 U1660 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1726), .Y(n1386) );
  MUX2X1 U1661 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1726), .Y(n1390) );
  MUX2X1 U1662 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1726), .Y(n1389) );
  MUX2X1 U1663 ( .B(n1388), .A(n1385), .S(n1702), .Y(n1392) );
  MUX2X1 U1664 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1726), .Y(n1396) );
  MUX2X1 U1665 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1726), .Y(n1395) );
  MUX2X1 U1666 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1726), .Y(n1399) );
  MUX2X1 U1667 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1726), .Y(n1398) );
  MUX2X1 U1668 ( .B(n1397), .A(n1394), .S(n1703), .Y(n1408) );
  MUX2X1 U1669 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1726), .Y(n1402) );
  MUX2X1 U1670 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1726), .Y(n1401) );
  MUX2X1 U1671 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1726), .Y(n1405) );
  MUX2X1 U1672 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1726), .Y(n1404) );
  MUX2X1 U1673 ( .B(n1403), .A(n1400), .S(n1702), .Y(n1407) );
  MUX2X1 U1674 ( .B(n1406), .A(n1391), .S(n1695), .Y(n1685) );
  MUX2X1 U1675 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1724), .Y(n1411) );
  MUX2X1 U1676 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1721), .Y(n1410) );
  MUX2X1 U1677 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1725), .Y(n1414) );
  MUX2X1 U1678 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1721), .Y(n1413) );
  MUX2X1 U1679 ( .B(n1412), .A(n1409), .S(n1702), .Y(n1423) );
  MUX2X1 U1680 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1721), .Y(n1417) );
  MUX2X1 U1681 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1721), .Y(n1416) );
  MUX2X1 U1682 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1730), .Y(n1420) );
  MUX2X1 U1683 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1721), .Y(n1419) );
  MUX2X1 U1684 ( .B(n1418), .A(n1415), .S(n1703), .Y(n1422) );
  MUX2X1 U1685 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1723), .Y(n1426) );
  MUX2X1 U1686 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1729), .Y(n1425) );
  MUX2X1 U1687 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1721), .Y(n1429) );
  MUX2X1 U1688 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1719), .Y(n1428) );
  MUX2X1 U1689 ( .B(n1427), .A(n1424), .S(n1703), .Y(n1438) );
  MUX2X1 U1690 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1730), .Y(n1432) );
  MUX2X1 U1691 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1729), .Y(n1431) );
  MUX2X1 U1692 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1723), .Y(n1435) );
  MUX2X1 U1693 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1730), .Y(n1434) );
  MUX2X1 U1694 ( .B(n1433), .A(n1430), .S(n1703), .Y(n1437) );
  MUX2X1 U1695 ( .B(n1436), .A(n1421), .S(n1695), .Y(n1686) );
  MUX2X1 U1696 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1730), .Y(n1441) );
  MUX2X1 U1697 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1730), .Y(n1440) );
  MUX2X1 U1698 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1723), .Y(n1444) );
  MUX2X1 U1699 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1723), .Y(n1443) );
  MUX2X1 U1700 ( .B(n1442), .A(n1439), .S(n1702), .Y(n1453) );
  MUX2X1 U1701 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1729), .Y(n1447) );
  MUX2X1 U1702 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1723), .Y(n1446) );
  MUX2X1 U1703 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1730), .Y(n1450) );
  MUX2X1 U1704 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1729), .Y(n1449) );
  MUX2X1 U1705 ( .B(n1448), .A(n1445), .S(n1702), .Y(n1452) );
  MUX2X1 U1706 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1727), .Y(n1456) );
  MUX2X1 U1707 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1727), .Y(n1455) );
  MUX2X1 U1708 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1727), .Y(n1459) );
  MUX2X1 U1709 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1727), .Y(n1458) );
  MUX2X1 U1710 ( .B(n1457), .A(n1454), .S(n1702), .Y(n1468) );
  MUX2X1 U1711 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1727), .Y(n1462) );
  MUX2X1 U1712 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1727), .Y(n1461) );
  MUX2X1 U1713 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1727), .Y(n1465) );
  MUX2X1 U1714 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1727), .Y(n1464) );
  MUX2X1 U1715 ( .B(n1463), .A(n1460), .S(n1702), .Y(n1467) );
  MUX2X1 U1716 ( .B(n1466), .A(n1451), .S(n1695), .Y(n1687) );
  MUX2X1 U1717 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1727), .Y(n1471) );
  MUX2X1 U1718 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1727), .Y(n1470) );
  MUX2X1 U1719 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1727), .Y(n1474) );
  MUX2X1 U1720 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1727), .Y(n1473) );
  MUX2X1 U1721 ( .B(n1472), .A(n1469), .S(n1701), .Y(n1483) );
  MUX2X1 U1722 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1728), .Y(n1477) );
  MUX2X1 U1723 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1728), .Y(n1476) );
  MUX2X1 U1724 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1728), .Y(n1480) );
  MUX2X1 U1725 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1728), .Y(n1479) );
  MUX2X1 U1726 ( .B(n1478), .A(n1475), .S(n1701), .Y(n1482) );
  MUX2X1 U1727 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1728), .Y(n1486) );
  MUX2X1 U1728 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1728), .Y(n1485) );
  MUX2X1 U1729 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1728), .Y(n1489) );
  MUX2X1 U1730 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1728), .Y(n1488) );
  MUX2X1 U1731 ( .B(n1487), .A(n1484), .S(n1701), .Y(n1498) );
  MUX2X1 U1732 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1728), .Y(n1492) );
  MUX2X1 U1733 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1728), .Y(n1491) );
  MUX2X1 U1734 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1728), .Y(n1495) );
  MUX2X1 U1735 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1728), .Y(n1494) );
  MUX2X1 U1736 ( .B(n1493), .A(n1490), .S(n1701), .Y(n1497) );
  MUX2X1 U1737 ( .B(n1496), .A(n1481), .S(n1695), .Y(n1688) );
  MUX2X1 U1738 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1721), .Y(n1501) );
  MUX2X1 U1739 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1725), .Y(n1500) );
  MUX2X1 U1740 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1720), .Y(n1504) );
  MUX2X1 U1741 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1723), .Y(n1503) );
  MUX2X1 U1742 ( .B(n1502), .A(n1499), .S(n1701), .Y(n1513) );
  MUX2X1 U1743 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1720), .Y(n1507) );
  MUX2X1 U1744 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1725), .Y(n1506) );
  MUX2X1 U1745 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1719), .Y(n1510) );
  MUX2X1 U1746 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1724), .Y(n1509) );
  MUX2X1 U1747 ( .B(n1508), .A(n1505), .S(n1701), .Y(n1512) );
  MUX2X1 U1748 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1730), .Y(n1516) );
  MUX2X1 U1749 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1726), .Y(n1515) );
  MUX2X1 U1750 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1723), .Y(n1519) );
  MUX2X1 U1751 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1729), .Y(n1518) );
  MUX2X1 U1752 ( .B(n1517), .A(n1514), .S(n1701), .Y(n1528) );
  MUX2X1 U1753 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1723), .Y(n1522) );
  MUX2X1 U1754 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1726), .Y(n1521) );
  MUX2X1 U1755 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1730), .Y(n1525) );
  MUX2X1 U1756 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1724), .Y(n1524) );
  MUX2X1 U1757 ( .B(n1523), .A(n1520), .S(n1701), .Y(n1527) );
  MUX2X1 U1758 ( .B(n1526), .A(n1511), .S(n1695), .Y(n1689) );
  MUX2X1 U1759 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1721), .Y(n1531) );
  MUX2X1 U1760 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1724), .Y(n1530) );
  MUX2X1 U1761 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1723), .Y(n1534) );
  MUX2X1 U1762 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1722), .Y(n1533) );
  MUX2X1 U1763 ( .B(n1532), .A(n1529), .S(n1701), .Y(n1543) );
  MUX2X1 U1764 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1721), .Y(n1537) );
  MUX2X1 U1765 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1726), .Y(n1536) );
  MUX2X1 U1766 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1725), .Y(n1540) );
  MUX2X1 U1767 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1719), .Y(n1539) );
  MUX2X1 U1768 ( .B(n1538), .A(n1535), .S(n1701), .Y(n1542) );
  MUX2X1 U1769 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1730), .Y(n1546) );
  MUX2X1 U1770 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1722), .Y(n1545) );
  MUX2X1 U1771 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1721), .Y(n1549) );
  MUX2X1 U1772 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1729), .Y(n1548) );
  MUX2X1 U1773 ( .B(n1547), .A(n1544), .S(n1701), .Y(n1558) );
  MUX2X1 U1774 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1720), .Y(n1552) );
  MUX2X1 U1775 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1719), .Y(n1551) );
  MUX2X1 U1776 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1725), .Y(n1555) );
  MUX2X1 U1777 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1724), .Y(n1554) );
  MUX2X1 U1778 ( .B(n1553), .A(n1550), .S(n1701), .Y(n1557) );
  MUX2X1 U1779 ( .B(n1556), .A(n1541), .S(n1695), .Y(n1690) );
  MUX2X1 U1780 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1719), .Y(n1561) );
  MUX2X1 U1781 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1725), .Y(n1560) );
  MUX2X1 U1782 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1721), .Y(n1564) );
  MUX2X1 U1783 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1729), .Y(n1563) );
  MUX2X1 U1784 ( .B(n1562), .A(n1559), .S(n1700), .Y(n1573) );
  MUX2X1 U1785 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1729), .Y(n1567) );
  MUX2X1 U1786 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1724), .Y(n1566) );
  MUX2X1 U1787 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1725), .Y(n1570) );
  MUX2X1 U1788 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1723), .Y(n1569) );
  MUX2X1 U1789 ( .B(n1568), .A(n1565), .S(n1700), .Y(n1572) );
  MUX2X1 U1790 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1729), .Y(n1576) );
  MUX2X1 U1791 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1730), .Y(n1575) );
  MUX2X1 U1792 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1730), .Y(n1579) );
  MUX2X1 U1793 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1725), .Y(n1578) );
  MUX2X1 U1794 ( .B(n1577), .A(n1574), .S(n1700), .Y(n1588) );
  MUX2X1 U1795 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1721), .Y(n1582) );
  MUX2X1 U1796 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1727), .Y(n1581) );
  MUX2X1 U1797 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1729), .Y(n1585) );
  MUX2X1 U1798 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1730), .Y(n1584) );
  MUX2X1 U1799 ( .B(n1583), .A(n1580), .S(n1700), .Y(n1587) );
  MUX2X1 U1800 ( .B(n1586), .A(n1571), .S(n1695), .Y(n1691) );
  MUX2X1 U1801 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1729), .Y(n1591) );
  MUX2X1 U1802 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1729), .Y(n1590) );
  MUX2X1 U1803 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1729), .Y(n1594) );
  MUX2X1 U1804 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1729), .Y(n1593) );
  MUX2X1 U1805 ( .B(n1592), .A(n1589), .S(n1700), .Y(n1603) );
  MUX2X1 U1806 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1729), .Y(n1597) );
  MUX2X1 U1807 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1729), .Y(n1596) );
  MUX2X1 U1808 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1729), .Y(n1600) );
  MUX2X1 U1809 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1729), .Y(n1599) );
  MUX2X1 U1810 ( .B(n1598), .A(n1595), .S(n1700), .Y(n1602) );
  MUX2X1 U1811 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1729), .Y(n1606) );
  MUX2X1 U1812 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1729), .Y(n1605) );
  MUX2X1 U1813 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1729), .Y(n1609) );
  MUX2X1 U1814 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1729), .Y(n1608) );
  MUX2X1 U1815 ( .B(n1607), .A(n1604), .S(n1700), .Y(n1618) );
  MUX2X1 U1816 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1721), .Y(n1612) );
  MUX2X1 U1817 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1725), .Y(n1611) );
  MUX2X1 U1818 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1725), .Y(n1615) );
  MUX2X1 U1819 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1724), .Y(n1614) );
  MUX2X1 U1820 ( .B(n1613), .A(n1610), .S(n1700), .Y(n1617) );
  MUX2X1 U1821 ( .B(n1616), .A(n1601), .S(n1695), .Y(n1692) );
  MUX2X1 U1822 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1725), .Y(n1621) );
  MUX2X1 U1823 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1719), .Y(n1620) );
  MUX2X1 U1824 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1724), .Y(n1624) );
  MUX2X1 U1825 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1729), .Y(n1623) );
  MUX2X1 U1826 ( .B(n1622), .A(n1619), .S(n1700), .Y(n1633) );
  MUX2X1 U1827 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1721), .Y(n1627) );
  MUX2X1 U1828 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1721), .Y(n1626) );
  MUX2X1 U1829 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1725), .Y(n1630) );
  MUX2X1 U1830 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1724), .Y(n1629) );
  MUX2X1 U1831 ( .B(n1628), .A(n1625), .S(n1700), .Y(n1632) );
  MUX2X1 U1832 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1730), .Y(n1636) );
  MUX2X1 U1833 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1730), .Y(n1635) );
  MUX2X1 U1834 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1730), .Y(n1639) );
  MUX2X1 U1835 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1730), .Y(n1638) );
  MUX2X1 U1836 ( .B(n1637), .A(n1634), .S(n1700), .Y(n1648) );
  MUX2X1 U1837 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1730), .Y(n1642) );
  MUX2X1 U1838 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1730), .Y(n1641) );
  MUX2X1 U1839 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1730), .Y(n1645) );
  MUX2X1 U1840 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1730), .Y(n1644) );
  MUX2X1 U1841 ( .B(n1643), .A(n1640), .S(n1700), .Y(n1647) );
  MUX2X1 U1842 ( .B(n1646), .A(n1631), .S(n1695), .Y(n1693) );
  MUX2X1 U1843 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1730), .Y(n1651) );
  MUX2X1 U1844 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1730), .Y(n1650) );
  MUX2X1 U1845 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1730), .Y(n1654) );
  MUX2X1 U1846 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1730), .Y(n1653) );
  MUX2X1 U1847 ( .B(n1652), .A(n1649), .S(n1700), .Y(n1663) );
  MUX2X1 U1848 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1724), .Y(n1657) );
  MUX2X1 U1849 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1728), .Y(n1656) );
  MUX2X1 U1850 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1728), .Y(n1660) );
  MUX2X1 U1851 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1719), .Y(n1659) );
  MUX2X1 U1852 ( .B(n1658), .A(n1655), .S(n1700), .Y(n1662) );
  MUX2X1 U1853 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1721), .Y(n1666) );
  MUX2X1 U1854 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1728), .Y(n1665) );
  MUX2X1 U1855 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1722), .Y(n1669) );
  MUX2X1 U1856 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1724), .Y(n1668) );
  MUX2X1 U1857 ( .B(n1667), .A(n1664), .S(n1700), .Y(n1678) );
  MUX2X1 U1858 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1723), .Y(n1672) );
  MUX2X1 U1859 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1727), .Y(n1671) );
  MUX2X1 U1860 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1723), .Y(n1675) );
  MUX2X1 U1861 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1720), .Y(n1674) );
  MUX2X1 U1862 ( .B(n1673), .A(n1670), .S(n1700), .Y(n1677) );
  MUX2X1 U1863 ( .B(n1676), .A(n1661), .S(n1695), .Y(n1694) );
  INVX1 U1864 ( .A(N11), .Y(n1867) );
  INVX1 U1865 ( .A(N10), .Y(n1865) );
  INVX8 U1866 ( .A(n1831), .Y(n1828) );
  INVX8 U1867 ( .A(n1831), .Y(n1829) );
  INVX8 U1868 ( .A(n1831), .Y(n1830) );
  INVX8 U1869 ( .A(n45), .Y(n1832) );
  INVX8 U1870 ( .A(n47), .Y(n1833) );
  INVX8 U1871 ( .A(n48), .Y(n1834) );
  INVX8 U1872 ( .A(n50), .Y(n1835) );
  INVX8 U1873 ( .A(n52), .Y(n1836) );
  INVX8 U1874 ( .A(n54), .Y(n1837) );
  INVX8 U1875 ( .A(n56), .Y(n1838) );
  INVX8 U1876 ( .A(n58), .Y(n1839) );
  INVX8 U1877 ( .A(n1869), .Y(n1868) );
  INVX8 U1878 ( .A(N12), .Y(n1869) );
endmodule


module memc_Size16_4 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1800), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1801), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1802), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1803), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1804), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1805), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1806), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1807), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1808), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1809), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1810), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1811), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1812), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1813), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1814), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1815), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1816), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1817), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1818), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1819), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1820), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1821), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1822), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1823), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1824), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1825), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1826), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1827), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1828), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1829), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1830), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1831), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1832), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1833), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1834), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1835), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1836), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1837), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1838), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1839), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1840), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1841), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1842), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1843), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1844), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1845), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1846), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1847), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1848), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1849), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1850), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1851), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1852), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1853), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1854), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1855), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1856), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1857), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1858), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1859), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1860), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1861), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1862), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1863), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1864), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1865), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1866), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1867), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1868), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1869), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1870), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1871), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1872), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1873), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1874), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1875), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1876), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1877), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1878), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1879), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1880), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1881), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1882), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1883), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1884), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1885), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1886), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1887), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1888), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1889), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1890), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1891), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1892), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1893), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1894), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1895), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1896), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1897), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1898), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1899), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1900), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1901), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1902), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1903), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1904), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1905), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1906), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1907), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1908), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1909), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1910), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1911), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1912), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1913), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1914), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1915), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1916), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1917), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1918), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1919), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1920), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1921), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1922), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1923), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1924), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1925), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1926), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1927), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1928), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1929), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1930), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1931), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1932), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1933), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1934), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1935), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1936), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1937), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1938), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1939), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1940), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1941), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1942), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1943), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1944), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1945), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1946), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1947), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1948), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1949), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1950), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1951), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1952), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1953), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1954), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1955), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1956), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1957), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1958), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1959), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1960), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1961), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1962), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n1963), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n1964), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n1965), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n1966), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n1967), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1968), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1969), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1970), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1971), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1972), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1973), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1974), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1975), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n1976), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n1977), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n1978), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n1979), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n1980), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n1981), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n1982), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n1983), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1984), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1985), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1986), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1987), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1988), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1989), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1990), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1991), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n1992), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n1993), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n1994), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n1995), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n1996), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n1997), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n1998), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n1999), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2000), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2001), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2002), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2003), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2004), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2005), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2006), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2007), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2008), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2009), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2010), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2011), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2012), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2013), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2014), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2015), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2016), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2017), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2018), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2019), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2020), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2021), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2022), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2023), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2024), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2025), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2026), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2027), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2028), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2029), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2030), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2031), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2032), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2033), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2034), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2035), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2036), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2037), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2038), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2039), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2040), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2041), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2042), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2043), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2044), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2045), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2046), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2047), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2048), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2049), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2050), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2051), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2052), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2053), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2054), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2055), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2056), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2057), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2058), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2059), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2060), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2061), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2062), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2063), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2064), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2065), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2066), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2067), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2068), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2069), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2070), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2071), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2072), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2073), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2074), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2075), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2076), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2077), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2078), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2079), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2080), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2081), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2082), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2083), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2084), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2085), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2086), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2087), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2088), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2089), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2090), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2091), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2092), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2093), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2094), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2095), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2096), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2097), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2098), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2099), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2100), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2101), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2102), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2103), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2104), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2105), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2106), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2107), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2108), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2109), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2110), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2111), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2112), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2113), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2114), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2115), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2116), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2117), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2118), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2119), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2120), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2121), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2122), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2123), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2124), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2125), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2126), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2127), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2128), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2129), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2130), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2131), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2132), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2133), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2134), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2135), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2136), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2137), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2138), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2139), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2140), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2141), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2142), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2143), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2144), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2145), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2146), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2147), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2148), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2149), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2150), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2151), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2152), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2153), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2154), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2155), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2156), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2157), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2158), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2159), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2160), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2161), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2162), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2163), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2164), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2165), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2166), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2167), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2168), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2169), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2170), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2171), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2172), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2173), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2174), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2175), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2176), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2177), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2178), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2179), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2180), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2181), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2182), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2183), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2184), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2185), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2186), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2187), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2188), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2189), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2190), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2191), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2192), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2193), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2194), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2195), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2196), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2197), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2198), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2199), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2200), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2201), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2202), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2203), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2204), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2205), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2206), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2207), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2208), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2209), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2210), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2211), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2212), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2213), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2214), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2215), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2216), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2217), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2218), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2219), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2220), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2221), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2222), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2223), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2224), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2225), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2226), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2227), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2228), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2229), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2230), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2231), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2232), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2233), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2234), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2235), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2236), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2237), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2238), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2239), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2240), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2241), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2242), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2243), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2244), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2245), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2246), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2247), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2248), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2249), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2250), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2251), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2252), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2253), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2254), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2255), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2256), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2257), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2258), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2259), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2260), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2261), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2262), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2263), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2264), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2265), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2266), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2267), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2268), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2269), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2270), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2271), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2272), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2273), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2274), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2275), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2276), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2277), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2278), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2279), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2280), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2281), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2282), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2283), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2284), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2285), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2286), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2287), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2288), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2289), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2290), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2291), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2292), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2293), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2295), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2296), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2297), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2298), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2299), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2300), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2301), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2302), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2303), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2304), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2305), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2306), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2307), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2308), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2309), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2310), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2311), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2312) );
  INVX1 U2 ( .A(n1200), .Y(n1209) );
  INVX1 U3 ( .A(n1199), .Y(n1211) );
  INVX1 U4 ( .A(n1199), .Y(n1212) );
  INVX2 U5 ( .A(N10), .Y(n1264) );
  INVX1 U6 ( .A(n8), .Y(n5) );
  INVX1 U7 ( .A(n1272), .Y(n1271) );
  INVX1 U8 ( .A(n1215), .Y(n1200) );
  INVX1 U9 ( .A(n1265), .Y(n1187) );
  INVX1 U10 ( .A(n1199), .Y(n1214) );
  INVX2 U11 ( .A(n1201), .Y(n1202) );
  INVX1 U12 ( .A(n1187), .Y(n1188) );
  INVX2 U13 ( .A(n1201), .Y(n1203) );
  INVX1 U14 ( .A(n1187), .Y(n1189) );
  INVX1 U15 ( .A(n1264), .Y(n1205) );
  INVX1 U16 ( .A(n1264), .Y(n1206) );
  INVX1 U17 ( .A(n1187), .Y(n1190) );
  INVX2 U18 ( .A(n1201), .Y(n1207) );
  INVX1 U19 ( .A(n1187), .Y(n1191) );
  INVX1 U20 ( .A(n1187), .Y(n1192) );
  INVX1 U21 ( .A(n1200), .Y(n1208) );
  INVX1 U22 ( .A(n1187), .Y(n1193) );
  INVX1 U23 ( .A(n1264), .Y(n1210) );
  INVX1 U24 ( .A(n1186), .Y(n1194) );
  INVX1 U25 ( .A(n1186), .Y(n1195) );
  INVX1 U26 ( .A(n1186), .Y(n1196) );
  INVX2 U27 ( .A(n1199), .Y(n1213) );
  INVX2 U28 ( .A(n1264), .Y(n1204) );
  INVX2 U29 ( .A(n1187), .Y(n1198) );
  INVX1 U30 ( .A(n1186), .Y(n1197) );
  INVX1 U31 ( .A(n1163), .Y(N32) );
  INVX1 U32 ( .A(n1164), .Y(N31) );
  INVX1 U33 ( .A(n1165), .Y(N30) );
  INVX1 U34 ( .A(n1167), .Y(N28) );
  INVX1 U35 ( .A(n1168), .Y(N27) );
  INVX1 U36 ( .A(n1169), .Y(N26) );
  INVX1 U37 ( .A(n1170), .Y(N25) );
  INVX1 U38 ( .A(n1173), .Y(N22) );
  INVX1 U39 ( .A(n1174), .Y(N21) );
  INVX1 U40 ( .A(n1175), .Y(N20) );
  INVX1 U41 ( .A(n1176), .Y(N19) );
  INVX1 U42 ( .A(n1177), .Y(N18) );
  INVX1 U43 ( .A(n1178), .Y(N17) );
  INVX1 U44 ( .A(n1166), .Y(N29) );
  INVX1 U45 ( .A(n1171), .Y(N24) );
  INVX1 U46 ( .A(n1172), .Y(N23) );
  INVX2 U47 ( .A(n1267), .Y(n1182) );
  INVX1 U48 ( .A(n1215), .Y(n1199) );
  INVX1 U49 ( .A(n1267), .Y(n1184) );
  INVX1 U50 ( .A(N12), .Y(n1267) );
  INVX1 U51 ( .A(n1267), .Y(n1183) );
  INVX1 U52 ( .A(n1267), .Y(n1185) );
  INVX1 U53 ( .A(N14), .Y(n1270) );
  INVX1 U54 ( .A(n1270), .Y(n1179) );
  INVX1 U55 ( .A(N13), .Y(n1268) );
  INVX1 U56 ( .A(n1268), .Y(n1181) );
  INVX1 U57 ( .A(n1268), .Y(n1180) );
  INVX1 U58 ( .A(n1265), .Y(n1186) );
  INVX1 U59 ( .A(n1264), .Y(n1215) );
  INVX1 U60 ( .A(n78), .Y(n1216) );
  INVX1 U61 ( .A(n79), .Y(n1219) );
  INVX1 U62 ( .A(n80), .Y(n1222) );
  INVX1 U63 ( .A(n81), .Y(n1225) );
  INVX1 U64 ( .A(n1263), .Y(n1201) );
  INVX4 U65 ( .A(n60), .Y(n165) );
  INVX4 U66 ( .A(n57), .Y(n156) );
  INVX4 U67 ( .A(n54), .Y(n147) );
  INVX4 U68 ( .A(n12), .Y(n84) );
  INVX4 U69 ( .A(n28), .Y(n87) );
  INVX4 U70 ( .A(n59), .Y(n162) );
  INVX4 U71 ( .A(n58), .Y(n159) );
  INVX4 U72 ( .A(n56), .Y(n153) );
  INVX4 U73 ( .A(n55), .Y(n150) );
  INVX4 U74 ( .A(n42), .Y(n123) );
  INVX4 U75 ( .A(n41), .Y(n120) );
  INVX4 U76 ( .A(n43), .Y(n124) );
  INVX4 U77 ( .A(n34), .Y(n103) );
  INVX4 U78 ( .A(n29), .Y(n90) );
  INVX4 U79 ( .A(n51), .Y(n144) );
  INVX4 U80 ( .A(n50), .Y(n141) );
  INVX4 U81 ( .A(n49), .Y(n138) );
  INVX4 U82 ( .A(n48), .Y(n135) );
  INVX4 U83 ( .A(n47), .Y(n132) );
  INVX4 U84 ( .A(n46), .Y(n129) );
  INVX4 U85 ( .A(n38), .Y(n115) );
  INVX4 U86 ( .A(n37), .Y(n112) );
  INVX4 U87 ( .A(n36), .Y(n109) );
  INVX4 U88 ( .A(n35), .Y(n106) );
  INVX4 U89 ( .A(n33), .Y(n102) );
  INVX4 U90 ( .A(n32), .Y(n99) );
  INVX4 U91 ( .A(n31), .Y(n96) );
  INVX4 U92 ( .A(n30), .Y(n93) );
  INVX1 U93 ( .A(n1231), .Y(n1230) );
  INVX4 U94 ( .A(n10), .Y(n1231) );
  BUFX2 U95 ( .A(n45), .Y(n1) );
  BUFX2 U96 ( .A(n40), .Y(n2) );
  BUFX2 U97 ( .A(n62), .Y(n3) );
  BUFX2 U98 ( .A(n53), .Y(n4) );
  OR2X2 U99 ( .A(n166), .B(n66), .Y(n6) );
  INVX1 U100 ( .A(n6), .Y(\data_out<15> ) );
  OR2X2 U101 ( .A(write), .B(n1271), .Y(n8) );
  INVX1 U102 ( .A(n8), .Y(n9) );
  AND2X2 U103 ( .A(n166), .B(n1272), .Y(n10) );
  AND2X2 U104 ( .A(\data_in<0> ), .B(n1229), .Y(n11) );
  AND2X2 U105 ( .A(n1229), .B(n82), .Y(n12) );
  AND2X2 U106 ( .A(\data_in<1> ), .B(n1228), .Y(n13) );
  AND2X2 U107 ( .A(\data_in<2> ), .B(n1228), .Y(n14) );
  AND2X2 U108 ( .A(\data_in<3> ), .B(n1229), .Y(n15) );
  AND2X2 U109 ( .A(\data_in<4> ), .B(n1228), .Y(n16) );
  AND2X2 U110 ( .A(\data_in<5> ), .B(n1229), .Y(n17) );
  AND2X2 U111 ( .A(\data_in<6> ), .B(n1228), .Y(n18) );
  AND2X2 U112 ( .A(\data_in<7> ), .B(n1228), .Y(n19) );
  AND2X2 U113 ( .A(\data_in<8> ), .B(n1228), .Y(n20) );
  AND2X2 U114 ( .A(\data_in<9> ), .B(n1228), .Y(n21) );
  AND2X2 U115 ( .A(\data_in<10> ), .B(n1229), .Y(n22) );
  AND2X2 U116 ( .A(\data_in<11> ), .B(n1229), .Y(n23) );
  AND2X2 U117 ( .A(\data_in<12> ), .B(n1228), .Y(n24) );
  AND2X2 U118 ( .A(\data_in<13> ), .B(n1228), .Y(n25) );
  AND2X2 U119 ( .A(\data_in<14> ), .B(n1228), .Y(n26) );
  AND2X2 U120 ( .A(\data_in<15> ), .B(n1228), .Y(n27) );
  AND2X2 U121 ( .A(n1228), .B(n85), .Y(n28) );
  AND2X2 U122 ( .A(n1228), .B(n88), .Y(n29) );
  AND2X2 U123 ( .A(n1228), .B(n91), .Y(n30) );
  AND2X2 U124 ( .A(n1229), .B(n94), .Y(n31) );
  AND2X2 U125 ( .A(n1228), .B(n97), .Y(n32) );
  AND2X2 U126 ( .A(n1229), .B(n100), .Y(n33) );
  AND2X2 U127 ( .A(n1229), .B(n78), .Y(n34) );
  AND2X2 U128 ( .A(n1229), .B(n104), .Y(n35) );
  AND2X2 U129 ( .A(n1228), .B(n107), .Y(n36) );
  AND2X2 U130 ( .A(n1228), .B(n110), .Y(n37) );
  AND2X2 U131 ( .A(n1228), .B(n113), .Y(n38) );
  AND2X2 U132 ( .A(n1230), .B(n116), .Y(n39) );
  INVX1 U133 ( .A(n39), .Y(n40) );
  AND2X2 U134 ( .A(n1228), .B(n118), .Y(n41) );
  AND2X2 U135 ( .A(n1229), .B(n121), .Y(n42) );
  AND2X2 U136 ( .A(n1228), .B(n79), .Y(n43) );
  AND2X2 U137 ( .A(n1230), .B(n125), .Y(n44) );
  INVX1 U138 ( .A(n44), .Y(n45) );
  AND2X2 U139 ( .A(n1228), .B(n127), .Y(n46) );
  AND2X2 U140 ( .A(n1229), .B(n130), .Y(n47) );
  AND2X2 U141 ( .A(n1228), .B(n133), .Y(n48) );
  AND2X2 U142 ( .A(n1228), .B(n136), .Y(n49) );
  AND2X2 U143 ( .A(n1229), .B(n139), .Y(n50) );
  AND2X2 U144 ( .A(n1228), .B(n142), .Y(n51) );
  AND2X2 U145 ( .A(n1230), .B(n80), .Y(n52) );
  INVX1 U146 ( .A(n52), .Y(n53) );
  AND2X2 U147 ( .A(n1228), .B(n145), .Y(n54) );
  AND2X2 U148 ( .A(n1229), .B(n148), .Y(n55) );
  AND2X2 U149 ( .A(n1228), .B(n151), .Y(n56) );
  AND2X2 U150 ( .A(n1228), .B(n154), .Y(n57) );
  AND2X2 U151 ( .A(n1229), .B(n157), .Y(n58) );
  AND2X2 U152 ( .A(n1228), .B(n160), .Y(n59) );
  AND2X2 U153 ( .A(n1228), .B(n163), .Y(n60) );
  AND2X2 U154 ( .A(n1230), .B(n81), .Y(n61) );
  INVX1 U155 ( .A(n61), .Y(n62) );
  BUFX2 U156 ( .A(n40), .Y(n1217) );
  BUFX2 U157 ( .A(n40), .Y(n1218) );
  BUFX2 U158 ( .A(n45), .Y(n1220) );
  BUFX2 U159 ( .A(n45), .Y(n1221) );
  BUFX2 U160 ( .A(n53), .Y(n1223) );
  BUFX2 U161 ( .A(n53), .Y(n1224) );
  BUFX2 U162 ( .A(n62), .Y(n1226) );
  BUFX2 U163 ( .A(n62), .Y(n1227) );
  INVX1 U164 ( .A(n1264), .Y(n1263) );
  AND2X1 U165 ( .A(n1184), .B(n1265), .Y(n63) );
  INVX1 U166 ( .A(n1266), .Y(n1265) );
  AND2X1 U167 ( .A(n2312), .B(n1269), .Y(n64) );
  INVX1 U168 ( .A(n1270), .Y(n1269) );
  AND2X1 U169 ( .A(N17), .B(n1272), .Y(n65) );
  INVX1 U170 ( .A(n65), .Y(n66) );
  BUFX2 U171 ( .A(n1305), .Y(n67) );
  INVX1 U172 ( .A(n67), .Y(n1697) );
  BUFX2 U173 ( .A(n1322), .Y(n68) );
  INVX1 U174 ( .A(n68), .Y(n1714) );
  BUFX2 U175 ( .A(n1339), .Y(n69) );
  INVX1 U176 ( .A(n69), .Y(n1731) );
  BUFX2 U177 ( .A(n1356), .Y(n70) );
  INVX1 U178 ( .A(n70), .Y(n1748) );
  BUFX2 U179 ( .A(n1373), .Y(n71) );
  INVX1 U180 ( .A(n71), .Y(n1765) );
  BUFX2 U181 ( .A(n1534), .Y(n72) );
  INVX1 U182 ( .A(n72), .Y(n1647) );
  BUFX2 U183 ( .A(n1664), .Y(n73) );
  INVX1 U184 ( .A(n73), .Y(n1782) );
  AND2X1 U185 ( .A(n1263), .B(n63), .Y(n74) );
  AND2X1 U186 ( .A(n1180), .B(n64), .Y(n75) );
  AND2X1 U187 ( .A(n1264), .B(n63), .Y(n76) );
  AND2X1 U188 ( .A(n1268), .B(n64), .Y(n77) );
  AND2X1 U189 ( .A(n75), .B(n1783), .Y(n78) );
  AND2X1 U190 ( .A(n1783), .B(n77), .Y(n79) );
  AND2X1 U191 ( .A(n1783), .B(n1647), .Y(n80) );
  AND2X1 U192 ( .A(n1783), .B(n1782), .Y(n81) );
  AND2X1 U193 ( .A(n74), .B(n75), .Y(n82) );
  INVX1 U194 ( .A(n82), .Y(n83) );
  AND2X1 U195 ( .A(n75), .B(n76), .Y(n85) );
  INVX1 U196 ( .A(n85), .Y(n86) );
  AND2X1 U197 ( .A(n75), .B(n1697), .Y(n88) );
  INVX1 U198 ( .A(n88), .Y(n89) );
  AND2X1 U199 ( .A(n75), .B(n1714), .Y(n91) );
  INVX1 U200 ( .A(n91), .Y(n92) );
  AND2X1 U201 ( .A(n75), .B(n1731), .Y(n94) );
  INVX1 U202 ( .A(n94), .Y(n95) );
  AND2X1 U203 ( .A(n75), .B(n1748), .Y(n97) );
  INVX1 U204 ( .A(n97), .Y(n98) );
  AND2X1 U205 ( .A(n75), .B(n1765), .Y(n100) );
  INVX1 U206 ( .A(n100), .Y(n101) );
  AND2X1 U207 ( .A(n74), .B(n77), .Y(n104) );
  INVX1 U208 ( .A(n104), .Y(n105) );
  AND2X1 U209 ( .A(n76), .B(n77), .Y(n107) );
  INVX1 U210 ( .A(n107), .Y(n108) );
  AND2X1 U211 ( .A(n1697), .B(n77), .Y(n110) );
  INVX1 U212 ( .A(n110), .Y(n111) );
  AND2X1 U213 ( .A(n1714), .B(n77), .Y(n113) );
  INVX1 U214 ( .A(n113), .Y(n114) );
  AND2X1 U215 ( .A(n1731), .B(n77), .Y(n116) );
  INVX1 U216 ( .A(n116), .Y(n117) );
  AND2X1 U217 ( .A(n1748), .B(n77), .Y(n118) );
  INVX1 U218 ( .A(n118), .Y(n119) );
  AND2X1 U219 ( .A(n1765), .B(n77), .Y(n121) );
  INVX1 U220 ( .A(n121), .Y(n122) );
  AND2X1 U221 ( .A(n74), .B(n1647), .Y(n125) );
  INVX1 U222 ( .A(n125), .Y(n126) );
  AND2X1 U223 ( .A(n76), .B(n1647), .Y(n127) );
  INVX1 U224 ( .A(n127), .Y(n128) );
  AND2X1 U225 ( .A(n1697), .B(n1647), .Y(n130) );
  INVX1 U226 ( .A(n130), .Y(n131) );
  AND2X1 U227 ( .A(n1714), .B(n1647), .Y(n133) );
  INVX1 U228 ( .A(n133), .Y(n134) );
  AND2X1 U229 ( .A(n1731), .B(n1647), .Y(n136) );
  INVX1 U230 ( .A(n136), .Y(n137) );
  AND2X1 U231 ( .A(n1748), .B(n1647), .Y(n139) );
  INVX1 U232 ( .A(n139), .Y(n140) );
  AND2X1 U233 ( .A(n1765), .B(n1647), .Y(n142) );
  INVX1 U234 ( .A(n142), .Y(n143) );
  AND2X1 U235 ( .A(n74), .B(n1782), .Y(n145) );
  INVX1 U236 ( .A(n145), .Y(n146) );
  AND2X1 U237 ( .A(n76), .B(n1782), .Y(n148) );
  INVX1 U238 ( .A(n148), .Y(n149) );
  AND2X1 U239 ( .A(n1697), .B(n1782), .Y(n151) );
  INVX1 U240 ( .A(n151), .Y(n152) );
  AND2X1 U241 ( .A(n1714), .B(n1782), .Y(n154) );
  INVX1 U242 ( .A(n154), .Y(n155) );
  AND2X1 U243 ( .A(n1731), .B(n1782), .Y(n157) );
  INVX1 U244 ( .A(n157), .Y(n158) );
  AND2X1 U245 ( .A(n1748), .B(n1782), .Y(n160) );
  INVX1 U246 ( .A(n160), .Y(n161) );
  AND2X1 U247 ( .A(n1765), .B(n1782), .Y(n163) );
  INVX1 U248 ( .A(n163), .Y(n164) );
  INVX1 U249 ( .A(rst), .Y(n1272) );
  BUFX2 U250 ( .A(write), .Y(n166) );
  INVX1 U251 ( .A(n8), .Y(n167) );
  INVX1 U252 ( .A(n8), .Y(n168) );
  INVX1 U253 ( .A(n8), .Y(n169) );
  MUX2X1 U254 ( .B(n171), .A(n172), .S(n1188), .Y(n170) );
  MUX2X1 U255 ( .B(n174), .A(n175), .S(n1188), .Y(n173) );
  MUX2X1 U256 ( .B(n177), .A(n178), .S(n1188), .Y(n176) );
  MUX2X1 U257 ( .B(n180), .A(n181), .S(n1188), .Y(n179) );
  MUX2X1 U258 ( .B(n183), .A(n184), .S(n1181), .Y(n182) );
  MUX2X1 U259 ( .B(n186), .A(n187), .S(n1188), .Y(n185) );
  MUX2X1 U260 ( .B(n189), .A(n190), .S(n1188), .Y(n188) );
  MUX2X1 U261 ( .B(n192), .A(n193), .S(n1188), .Y(n191) );
  MUX2X1 U262 ( .B(n195), .A(n196), .S(n1188), .Y(n194) );
  MUX2X1 U263 ( .B(n198), .A(n199), .S(n1181), .Y(n197) );
  MUX2X1 U264 ( .B(n201), .A(n202), .S(n1189), .Y(n200) );
  MUX2X1 U265 ( .B(n204), .A(n205), .S(n1189), .Y(n203) );
  MUX2X1 U266 ( .B(n207), .A(n208), .S(n1189), .Y(n206) );
  MUX2X1 U267 ( .B(n210), .A(n211), .S(n1189), .Y(n209) );
  MUX2X1 U268 ( .B(n213), .A(n215), .S(n1181), .Y(n212) );
  MUX2X1 U269 ( .B(n217), .A(n218), .S(n1189), .Y(n216) );
  MUX2X1 U270 ( .B(n220), .A(n221), .S(n1189), .Y(n219) );
  MUX2X1 U271 ( .B(n223), .A(n224), .S(n1189), .Y(n222) );
  MUX2X1 U272 ( .B(n226), .A(n227), .S(n1189), .Y(n225) );
  MUX2X1 U273 ( .B(n229), .A(n230), .S(n1181), .Y(n228) );
  MUX2X1 U274 ( .B(n232), .A(n233), .S(n1189), .Y(n231) );
  MUX2X1 U275 ( .B(n235), .A(n236), .S(n1189), .Y(n234) );
  MUX2X1 U276 ( .B(n238), .A(n239), .S(n1189), .Y(n237) );
  MUX2X1 U277 ( .B(n241), .A(n242), .S(n1189), .Y(n240) );
  MUX2X1 U278 ( .B(n244), .A(n245), .S(n1181), .Y(n243) );
  MUX2X1 U279 ( .B(n247), .A(n248), .S(n1190), .Y(n246) );
  MUX2X1 U280 ( .B(n250), .A(n251), .S(n1190), .Y(n249) );
  MUX2X1 U281 ( .B(n253), .A(n254), .S(n1190), .Y(n252) );
  MUX2X1 U282 ( .B(n256), .A(n257), .S(n1190), .Y(n255) );
  MUX2X1 U283 ( .B(n259), .A(n260), .S(n1181), .Y(n258) );
  MUX2X1 U284 ( .B(n262), .A(n263), .S(n1190), .Y(n261) );
  MUX2X1 U285 ( .B(n265), .A(n266), .S(n1190), .Y(n264) );
  MUX2X1 U286 ( .B(n268), .A(n269), .S(n1190), .Y(n267) );
  MUX2X1 U287 ( .B(n271), .A(n272), .S(n1190), .Y(n270) );
  MUX2X1 U288 ( .B(n274), .A(n275), .S(n1181), .Y(n273) );
  MUX2X1 U289 ( .B(n277), .A(n278), .S(n1190), .Y(n276) );
  MUX2X1 U290 ( .B(n280), .A(n281), .S(n1190), .Y(n279) );
  MUX2X1 U291 ( .B(n283), .A(n284), .S(n1190), .Y(n282) );
  MUX2X1 U292 ( .B(n286), .A(n287), .S(n1190), .Y(n285) );
  MUX2X1 U293 ( .B(n289), .A(n290), .S(n1181), .Y(n288) );
  MUX2X1 U294 ( .B(n292), .A(n293), .S(n1191), .Y(n291) );
  MUX2X1 U295 ( .B(n295), .A(n296), .S(n1191), .Y(n294) );
  MUX2X1 U296 ( .B(n298), .A(n299), .S(n1191), .Y(n297) );
  MUX2X1 U297 ( .B(n301), .A(n302), .S(n1191), .Y(n300) );
  MUX2X1 U298 ( .B(n304), .A(n305), .S(n1181), .Y(n303) );
  MUX2X1 U299 ( .B(n307), .A(n308), .S(n1191), .Y(n306) );
  MUX2X1 U300 ( .B(n310), .A(n311), .S(n1191), .Y(n309) );
  MUX2X1 U301 ( .B(n313), .A(n314), .S(n1191), .Y(n312) );
  MUX2X1 U302 ( .B(n316), .A(n317), .S(n1191), .Y(n315) );
  MUX2X1 U303 ( .B(n319), .A(n320), .S(n1181), .Y(n318) );
  MUX2X1 U304 ( .B(n322), .A(n323), .S(n1191), .Y(n321) );
  MUX2X1 U305 ( .B(n325), .A(n326), .S(n1191), .Y(n324) );
  MUX2X1 U306 ( .B(n328), .A(n329), .S(n1191), .Y(n327) );
  MUX2X1 U307 ( .B(n331), .A(n332), .S(n1191), .Y(n330) );
  MUX2X1 U308 ( .B(n334), .A(n335), .S(n1181), .Y(n333) );
  MUX2X1 U309 ( .B(n337), .A(n338), .S(n1192), .Y(n336) );
  MUX2X1 U310 ( .B(n340), .A(n341), .S(n1192), .Y(n339) );
  MUX2X1 U311 ( .B(n343), .A(n344), .S(n1192), .Y(n342) );
  MUX2X1 U312 ( .B(n346), .A(n347), .S(n1192), .Y(n345) );
  MUX2X1 U313 ( .B(n349), .A(n350), .S(n1181), .Y(n348) );
  MUX2X1 U314 ( .B(n352), .A(n353), .S(n1192), .Y(n351) );
  MUX2X1 U315 ( .B(n355), .A(n356), .S(n1192), .Y(n354) );
  MUX2X1 U316 ( .B(n358), .A(n359), .S(n1192), .Y(n357) );
  MUX2X1 U317 ( .B(n361), .A(n362), .S(n1192), .Y(n360) );
  MUX2X1 U318 ( .B(n364), .A(n365), .S(n1180), .Y(n363) );
  MUX2X1 U319 ( .B(n367), .A(n368), .S(n1192), .Y(n366) );
  MUX2X1 U320 ( .B(n370), .A(n371), .S(n1192), .Y(n369) );
  MUX2X1 U321 ( .B(n373), .A(n374), .S(n1192), .Y(n372) );
  MUX2X1 U322 ( .B(n376), .A(n377), .S(n1192), .Y(n375) );
  MUX2X1 U323 ( .B(n379), .A(n380), .S(n1180), .Y(n378) );
  MUX2X1 U324 ( .B(n382), .A(n383), .S(n1193), .Y(n381) );
  MUX2X1 U325 ( .B(n385), .A(n386), .S(n1193), .Y(n384) );
  MUX2X1 U326 ( .B(n388), .A(n389), .S(n1193), .Y(n387) );
  MUX2X1 U327 ( .B(n391), .A(n392), .S(n1193), .Y(n390) );
  MUX2X1 U328 ( .B(n394), .A(n395), .S(n1180), .Y(n393) );
  MUX2X1 U329 ( .B(n397), .A(n398), .S(n1193), .Y(n396) );
  MUX2X1 U330 ( .B(n400), .A(n401), .S(n1193), .Y(n399) );
  MUX2X1 U331 ( .B(n403), .A(n404), .S(n1193), .Y(n402) );
  MUX2X1 U332 ( .B(n406), .A(n407), .S(n1193), .Y(n405) );
  MUX2X1 U333 ( .B(n409), .A(n410), .S(n1180), .Y(n408) );
  MUX2X1 U334 ( .B(n412), .A(n413), .S(n1193), .Y(n411) );
  MUX2X1 U335 ( .B(n415), .A(n416), .S(n1193), .Y(n414) );
  MUX2X1 U336 ( .B(n418), .A(n419), .S(n1193), .Y(n417) );
  MUX2X1 U337 ( .B(n421), .A(n422), .S(n1193), .Y(n420) );
  MUX2X1 U338 ( .B(n424), .A(n425), .S(n1180), .Y(n423) );
  MUX2X1 U339 ( .B(n427), .A(n428), .S(n1194), .Y(n426) );
  MUX2X1 U340 ( .B(n430), .A(n431), .S(n1194), .Y(n429) );
  MUX2X1 U341 ( .B(n433), .A(n434), .S(n1194), .Y(n432) );
  MUX2X1 U342 ( .B(n436), .A(n437), .S(n1194), .Y(n435) );
  MUX2X1 U343 ( .B(n439), .A(n440), .S(n1180), .Y(n438) );
  MUX2X1 U344 ( .B(n442), .A(n443), .S(n1194), .Y(n441) );
  MUX2X1 U345 ( .B(n445), .A(n446), .S(n1194), .Y(n444) );
  MUX2X1 U346 ( .B(n448), .A(n449), .S(n1194), .Y(n447) );
  MUX2X1 U347 ( .B(n451), .A(n452), .S(n1194), .Y(n450) );
  MUX2X1 U348 ( .B(n454), .A(n455), .S(n1180), .Y(n453) );
  MUX2X1 U349 ( .B(n457), .A(n458), .S(n1194), .Y(n456) );
  MUX2X1 U350 ( .B(n460), .A(n461), .S(n1194), .Y(n459) );
  MUX2X1 U351 ( .B(n463), .A(n464), .S(n1194), .Y(n462) );
  MUX2X1 U352 ( .B(n466), .A(n467), .S(n1194), .Y(n465) );
  MUX2X1 U353 ( .B(n469), .A(n470), .S(n1180), .Y(n468) );
  MUX2X1 U354 ( .B(n472), .A(n473), .S(n1195), .Y(n471) );
  MUX2X1 U355 ( .B(n475), .A(n476), .S(n1195), .Y(n474) );
  MUX2X1 U356 ( .B(n478), .A(n479), .S(n1195), .Y(n477) );
  MUX2X1 U357 ( .B(n481), .A(n482), .S(n1195), .Y(n480) );
  MUX2X1 U358 ( .B(n484), .A(n485), .S(n1180), .Y(n483) );
  MUX2X1 U359 ( .B(n487), .A(n488), .S(n1195), .Y(n486) );
  MUX2X1 U360 ( .B(n490), .A(n491), .S(n1195), .Y(n489) );
  MUX2X1 U361 ( .B(n493), .A(n494), .S(n1195), .Y(n492) );
  MUX2X1 U362 ( .B(n496), .A(n497), .S(n1195), .Y(n495) );
  MUX2X1 U363 ( .B(n499), .A(n500), .S(n1180), .Y(n498) );
  MUX2X1 U364 ( .B(n502), .A(n503), .S(n1195), .Y(n501) );
  MUX2X1 U365 ( .B(n505), .A(n506), .S(n1195), .Y(n504) );
  MUX2X1 U366 ( .B(n508), .A(n509), .S(n1195), .Y(n507) );
  MUX2X1 U367 ( .B(n511), .A(n512), .S(n1195), .Y(n510) );
  MUX2X1 U368 ( .B(n514), .A(n515), .S(n1180), .Y(n513) );
  MUX2X1 U369 ( .B(n517), .A(n518), .S(n1196), .Y(n516) );
  MUX2X1 U370 ( .B(n520), .A(n521), .S(n1196), .Y(n519) );
  MUX2X1 U371 ( .B(n523), .A(n524), .S(n1196), .Y(n522) );
  MUX2X1 U372 ( .B(n526), .A(n527), .S(n1196), .Y(n525) );
  MUX2X1 U373 ( .B(n529), .A(n530), .S(n1180), .Y(n528) );
  MUX2X1 U374 ( .B(n532), .A(n533), .S(n1196), .Y(n531) );
  MUX2X1 U375 ( .B(n535), .A(n536), .S(n1196), .Y(n534) );
  MUX2X1 U376 ( .B(n538), .A(n539), .S(n1196), .Y(n537) );
  MUX2X1 U377 ( .B(n541), .A(n542), .S(n1196), .Y(n540) );
  MUX2X1 U378 ( .B(n544), .A(n545), .S(n1181), .Y(n543) );
  MUX2X1 U379 ( .B(n547), .A(n548), .S(n1196), .Y(n546) );
  MUX2X1 U380 ( .B(n550), .A(n551), .S(n1196), .Y(n549) );
  MUX2X1 U381 ( .B(n553), .A(n554), .S(n1196), .Y(n552) );
  MUX2X1 U382 ( .B(n556), .A(n557), .S(n1196), .Y(n555) );
  MUX2X1 U383 ( .B(n559), .A(n560), .S(n1181), .Y(n558) );
  MUX2X1 U384 ( .B(n562), .A(n563), .S(n1197), .Y(n561) );
  MUX2X1 U385 ( .B(n565), .A(n566), .S(n1197), .Y(n564) );
  MUX2X1 U386 ( .B(n568), .A(n569), .S(n1197), .Y(n567) );
  MUX2X1 U387 ( .B(n571), .A(n572), .S(n1197), .Y(n570) );
  MUX2X1 U388 ( .B(n574), .A(n575), .S(n1180), .Y(n573) );
  MUX2X1 U389 ( .B(n577), .A(n578), .S(n1197), .Y(n576) );
  MUX2X1 U390 ( .B(n580), .A(n581), .S(n1197), .Y(n579) );
  MUX2X1 U391 ( .B(n583), .A(n584), .S(n1197), .Y(n582) );
  MUX2X1 U392 ( .B(n586), .A(n587), .S(n1197), .Y(n585) );
  MUX2X1 U393 ( .B(n589), .A(n590), .S(n1181), .Y(n588) );
  MUX2X1 U394 ( .B(n592), .A(n593), .S(n1197), .Y(n591) );
  MUX2X1 U395 ( .B(n595), .A(n596), .S(n1197), .Y(n594) );
  MUX2X1 U396 ( .B(n598), .A(n599), .S(n1197), .Y(n597) );
  MUX2X1 U397 ( .B(n601), .A(n602), .S(n1197), .Y(n600) );
  MUX2X1 U398 ( .B(n604), .A(n605), .S(n1181), .Y(n603) );
  MUX2X1 U399 ( .B(n607), .A(n608), .S(n1198), .Y(n606) );
  MUX2X1 U400 ( .B(n610), .A(n611), .S(n1198), .Y(n609) );
  MUX2X1 U401 ( .B(n613), .A(n614), .S(n1198), .Y(n612) );
  MUX2X1 U402 ( .B(n616), .A(n617), .S(n1198), .Y(n615) );
  MUX2X1 U403 ( .B(n619), .A(n620), .S(n1181), .Y(n618) );
  MUX2X1 U404 ( .B(n622), .A(n623), .S(n1198), .Y(n621) );
  MUX2X1 U405 ( .B(n625), .A(n626), .S(n1198), .Y(n624) );
  MUX2X1 U406 ( .B(n628), .A(n629), .S(n1198), .Y(n627) );
  MUX2X1 U407 ( .B(n631), .A(n632), .S(n1198), .Y(n630) );
  MUX2X1 U408 ( .B(n634), .A(n635), .S(n1180), .Y(n633) );
  MUX2X1 U409 ( .B(n637), .A(n638), .S(n1198), .Y(n636) );
  MUX2X1 U410 ( .B(n640), .A(n641), .S(n1198), .Y(n639) );
  MUX2X1 U411 ( .B(n643), .A(n644), .S(n1198), .Y(n642) );
  MUX2X1 U412 ( .B(n646), .A(n647), .S(n1198), .Y(n645) );
  MUX2X1 U413 ( .B(n649), .A(n650), .S(n1180), .Y(n648) );
  MUX2X1 U414 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1208), .Y(n172) );
  MUX2X1 U415 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1204), .Y(n171) );
  MUX2X1 U416 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1211), .Y(n175) );
  MUX2X1 U417 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1206), .Y(n174) );
  MUX2X1 U418 ( .B(n173), .A(n170), .S(n1185), .Y(n184) );
  MUX2X1 U419 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1202), .Y(n178) );
  MUX2X1 U420 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1202), .Y(n177) );
  MUX2X1 U421 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1202), .Y(n181) );
  MUX2X1 U422 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1202), .Y(n180) );
  MUX2X1 U423 ( .B(n179), .A(n176), .S(n1185), .Y(n183) );
  MUX2X1 U424 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1202), .Y(n187) );
  MUX2X1 U425 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1202), .Y(n186) );
  MUX2X1 U426 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1202), .Y(n190) );
  MUX2X1 U427 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1202), .Y(n189) );
  MUX2X1 U428 ( .B(n188), .A(n185), .S(n1185), .Y(n199) );
  MUX2X1 U429 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1202), .Y(n193) );
  MUX2X1 U430 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1202), .Y(n192) );
  MUX2X1 U431 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1202), .Y(n196) );
  MUX2X1 U432 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1202), .Y(n195) );
  MUX2X1 U433 ( .B(n194), .A(n191), .S(n1185), .Y(n198) );
  MUX2X1 U434 ( .B(n197), .A(n182), .S(n1179), .Y(n1163) );
  MUX2X1 U435 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1203), .Y(n202) );
  MUX2X1 U436 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1203), .Y(n201) );
  MUX2X1 U437 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1203), .Y(n205) );
  MUX2X1 U438 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1203), .Y(n204) );
  MUX2X1 U439 ( .B(n203), .A(n200), .S(n1185), .Y(n215) );
  MUX2X1 U440 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1203), .Y(n208) );
  MUX2X1 U441 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1203), .Y(n207) );
  MUX2X1 U442 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1203), .Y(n211) );
  MUX2X1 U443 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1203), .Y(n210) );
  MUX2X1 U444 ( .B(n209), .A(n206), .S(n1185), .Y(n213) );
  MUX2X1 U445 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1203), .Y(n218) );
  MUX2X1 U446 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1203), .Y(n217) );
  MUX2X1 U447 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1203), .Y(n221) );
  MUX2X1 U448 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1203), .Y(n220) );
  MUX2X1 U449 ( .B(n219), .A(n216), .S(n1185), .Y(n230) );
  MUX2X1 U450 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1204), .Y(n224) );
  MUX2X1 U451 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1204), .Y(n223) );
  MUX2X1 U452 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1204), .Y(n227) );
  MUX2X1 U453 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1204), .Y(n226) );
  MUX2X1 U454 ( .B(n225), .A(n222), .S(n1185), .Y(n229) );
  MUX2X1 U455 ( .B(n228), .A(n212), .S(n1179), .Y(n1164) );
  MUX2X1 U456 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1204), .Y(n233) );
  MUX2X1 U457 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1204), .Y(n232) );
  MUX2X1 U458 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1204), .Y(n236) );
  MUX2X1 U459 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1204), .Y(n235) );
  MUX2X1 U460 ( .B(n234), .A(n231), .S(n1185), .Y(n245) );
  MUX2X1 U461 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1204), .Y(n239) );
  MUX2X1 U462 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1204), .Y(n238) );
  MUX2X1 U463 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1204), .Y(n242) );
  MUX2X1 U464 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1204), .Y(n241) );
  MUX2X1 U465 ( .B(n240), .A(n237), .S(n1185), .Y(n244) );
  MUX2X1 U466 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1205), .Y(n248) );
  MUX2X1 U467 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1205), .Y(n247) );
  MUX2X1 U468 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1205), .Y(n251) );
  MUX2X1 U469 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1205), .Y(n250) );
  MUX2X1 U470 ( .B(n249), .A(n246), .S(n1185), .Y(n260) );
  MUX2X1 U471 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1205), .Y(n254) );
  MUX2X1 U472 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1205), .Y(n253) );
  MUX2X1 U473 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1205), .Y(n257) );
  MUX2X1 U474 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1205), .Y(n256) );
  MUX2X1 U475 ( .B(n255), .A(n252), .S(n1185), .Y(n259) );
  MUX2X1 U476 ( .B(n258), .A(n243), .S(n1179), .Y(n1165) );
  MUX2X1 U477 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1205), .Y(n263) );
  MUX2X1 U478 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1205), .Y(n262) );
  MUX2X1 U479 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1205), .Y(n266) );
  MUX2X1 U480 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1205), .Y(n265) );
  MUX2X1 U481 ( .B(n264), .A(n261), .S(n1184), .Y(n275) );
  MUX2X1 U482 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1206), .Y(n269) );
  MUX2X1 U483 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1206), .Y(n268) );
  MUX2X1 U484 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1206), .Y(n272) );
  MUX2X1 U485 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1206), .Y(n271) );
  MUX2X1 U486 ( .B(n270), .A(n267), .S(n1184), .Y(n274) );
  MUX2X1 U487 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1206), .Y(n278) );
  MUX2X1 U488 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1206), .Y(n277) );
  MUX2X1 U489 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1206), .Y(n281) );
  MUX2X1 U490 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1206), .Y(n280) );
  MUX2X1 U491 ( .B(n279), .A(n276), .S(n1184), .Y(n290) );
  MUX2X1 U492 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1206), .Y(n284) );
  MUX2X1 U493 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1206), .Y(n283) );
  MUX2X1 U494 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1206), .Y(n287) );
  MUX2X1 U495 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1206), .Y(n286) );
  MUX2X1 U496 ( .B(n285), .A(n282), .S(n1184), .Y(n289) );
  MUX2X1 U497 ( .B(n288), .A(n273), .S(n1179), .Y(n1166) );
  MUX2X1 U498 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1207), .Y(n293) );
  MUX2X1 U499 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1207), .Y(n292) );
  MUX2X1 U500 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1207), .Y(n296) );
  MUX2X1 U501 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1207), .Y(n295) );
  MUX2X1 U502 ( .B(n294), .A(n291), .S(n1184), .Y(n305) );
  MUX2X1 U503 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1207), .Y(n299) );
  MUX2X1 U504 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1207), .Y(n298) );
  MUX2X1 U505 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1207), .Y(n302) );
  MUX2X1 U506 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1207), .Y(n301) );
  MUX2X1 U507 ( .B(n300), .A(n297), .S(n1184), .Y(n304) );
  MUX2X1 U508 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1207), .Y(n308) );
  MUX2X1 U509 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1207), .Y(n307) );
  MUX2X1 U510 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1207), .Y(n311) );
  MUX2X1 U511 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1207), .Y(n310) );
  MUX2X1 U512 ( .B(n309), .A(n306), .S(n1184), .Y(n320) );
  MUX2X1 U513 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1213), .Y(n314) );
  MUX2X1 U514 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1213), .Y(n313) );
  MUX2X1 U515 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1213), .Y(n317) );
  MUX2X1 U516 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1213), .Y(n316) );
  MUX2X1 U517 ( .B(n315), .A(n312), .S(n1184), .Y(n319) );
  MUX2X1 U518 ( .B(n318), .A(n303), .S(n1179), .Y(n1167) );
  MUX2X1 U519 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1213), .Y(n323) );
  MUX2X1 U520 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1213), .Y(n322) );
  MUX2X1 U521 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1213), .Y(n326) );
  MUX2X1 U522 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1213), .Y(n325) );
  MUX2X1 U523 ( .B(n324), .A(n321), .S(n1184), .Y(n335) );
  MUX2X1 U524 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1213), .Y(n329) );
  MUX2X1 U525 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1213), .Y(n328) );
  MUX2X1 U526 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1213), .Y(n332) );
  MUX2X1 U527 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1213), .Y(n331) );
  MUX2X1 U528 ( .B(n330), .A(n327), .S(n1184), .Y(n334) );
  MUX2X1 U529 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1207), .Y(n338) );
  MUX2X1 U530 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1213), .Y(n337) );
  MUX2X1 U531 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1213), .Y(n341) );
  MUX2X1 U532 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1213), .Y(n340) );
  MUX2X1 U533 ( .B(n339), .A(n336), .S(n1184), .Y(n350) );
  MUX2X1 U534 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1207), .Y(n344) );
  MUX2X1 U535 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1213), .Y(n343) );
  MUX2X1 U536 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1213), .Y(n347) );
  MUX2X1 U537 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1213), .Y(n346) );
  MUX2X1 U538 ( .B(n345), .A(n342), .S(n1184), .Y(n349) );
  MUX2X1 U539 ( .B(n348), .A(n333), .S(n1179), .Y(n1168) );
  MUX2X1 U540 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1213), .Y(n353) );
  MUX2X1 U541 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1213), .Y(n352) );
  MUX2X1 U542 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1202), .Y(n356) );
  MUX2X1 U543 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1207), .Y(n355) );
  MUX2X1 U544 ( .B(n354), .A(n351), .S(n1183), .Y(n365) );
  MUX2X1 U545 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1209), .Y(n359) );
  MUX2X1 U546 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1204), .Y(n358) );
  MUX2X1 U547 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1204), .Y(n362) );
  MUX2X1 U548 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1212), .Y(n361) );
  MUX2X1 U549 ( .B(n360), .A(n357), .S(n1183), .Y(n364) );
  MUX2X1 U550 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1212), .Y(n368) );
  MUX2X1 U551 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1211), .Y(n367) );
  MUX2X1 U552 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1204), .Y(n371) );
  MUX2X1 U553 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1204), .Y(n370) );
  MUX2X1 U554 ( .B(n369), .A(n366), .S(n1183), .Y(n380) );
  MUX2X1 U555 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1209), .Y(n374) );
  MUX2X1 U556 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1204), .Y(n373) );
  MUX2X1 U557 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1212), .Y(n377) );
  MUX2X1 U558 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1211), .Y(n376) );
  MUX2X1 U559 ( .B(n375), .A(n372), .S(n1183), .Y(n379) );
  MUX2X1 U560 ( .B(n378), .A(n363), .S(n1179), .Y(n1169) );
  MUX2X1 U561 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1208), .Y(n383) );
  MUX2X1 U562 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1208), .Y(n382) );
  MUX2X1 U563 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1208), .Y(n386) );
  MUX2X1 U564 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1208), .Y(n385) );
  MUX2X1 U565 ( .B(n384), .A(n381), .S(n1183), .Y(n395) );
  MUX2X1 U566 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1208), .Y(n389) );
  MUX2X1 U567 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1208), .Y(n388) );
  MUX2X1 U568 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1208), .Y(n392) );
  MUX2X1 U569 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1208), .Y(n391) );
  MUX2X1 U570 ( .B(n390), .A(n387), .S(n1183), .Y(n394) );
  MUX2X1 U571 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1208), .Y(n398) );
  MUX2X1 U572 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1208), .Y(n397) );
  MUX2X1 U573 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1208), .Y(n401) );
  MUX2X1 U574 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1208), .Y(n400) );
  MUX2X1 U575 ( .B(n399), .A(n396), .S(n1183), .Y(n410) );
  MUX2X1 U576 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1209), .Y(n404) );
  MUX2X1 U577 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1209), .Y(n403) );
  MUX2X1 U578 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1209), .Y(n407) );
  MUX2X1 U579 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1209), .Y(n406) );
  MUX2X1 U580 ( .B(n405), .A(n402), .S(n1183), .Y(n409) );
  MUX2X1 U581 ( .B(n408), .A(n393), .S(n1179), .Y(n1170) );
  MUX2X1 U582 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1209), .Y(n413) );
  MUX2X1 U583 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1209), .Y(n412) );
  MUX2X1 U584 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1209), .Y(n416) );
  MUX2X1 U585 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1209), .Y(n415) );
  MUX2X1 U586 ( .B(n414), .A(n411), .S(n1183), .Y(n425) );
  MUX2X1 U587 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1209), .Y(n419) );
  MUX2X1 U588 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1209), .Y(n418) );
  MUX2X1 U589 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1209), .Y(n422) );
  MUX2X1 U590 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1209), .Y(n421) );
  MUX2X1 U591 ( .B(n420), .A(n417), .S(n1183), .Y(n424) );
  MUX2X1 U592 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1210), .Y(n428) );
  MUX2X1 U593 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1210), .Y(n427) );
  MUX2X1 U594 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1210), .Y(n431) );
  MUX2X1 U595 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1210), .Y(n430) );
  MUX2X1 U596 ( .B(n429), .A(n426), .S(n1183), .Y(n440) );
  MUX2X1 U597 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1210), .Y(n434) );
  MUX2X1 U598 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1210), .Y(n433) );
  MUX2X1 U599 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1210), .Y(n437) );
  MUX2X1 U600 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1210), .Y(n436) );
  MUX2X1 U601 ( .B(n435), .A(n432), .S(n1183), .Y(n439) );
  MUX2X1 U602 ( .B(n438), .A(n423), .S(n1179), .Y(n1171) );
  MUX2X1 U603 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1210), .Y(n443) );
  MUX2X1 U604 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1210), .Y(n442) );
  MUX2X1 U605 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1210), .Y(n446) );
  MUX2X1 U606 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1210), .Y(n445) );
  MUX2X1 U607 ( .B(n444), .A(n441), .S(n1182), .Y(n455) );
  MUX2X1 U608 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1210), .Y(n449) );
  MUX2X1 U609 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1204), .Y(n448) );
  MUX2X1 U610 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1210), .Y(n452) );
  MUX2X1 U611 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1204), .Y(n451) );
  MUX2X1 U612 ( .B(n450), .A(n447), .S(n1182), .Y(n454) );
  MUX2X1 U613 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1204), .Y(n458) );
  MUX2X1 U614 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1208), .Y(n457) );
  MUX2X1 U615 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1204), .Y(n461) );
  MUX2X1 U616 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1204), .Y(n460) );
  MUX2X1 U617 ( .B(n459), .A(n456), .S(n1182), .Y(n470) );
  MUX2X1 U618 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1204), .Y(n464) );
  MUX2X1 U619 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1208), .Y(n463) );
  MUX2X1 U620 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1204), .Y(n467) );
  MUX2X1 U621 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1204), .Y(n466) );
  MUX2X1 U622 ( .B(n465), .A(n462), .S(n1182), .Y(n469) );
  MUX2X1 U623 ( .B(n468), .A(n453), .S(n1179), .Y(n1172) );
  MUX2X1 U624 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1203), .Y(n473) );
  MUX2X1 U625 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1202), .Y(n472) );
  MUX2X1 U626 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1206), .Y(n476) );
  MUX2X1 U627 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1210), .Y(n475) );
  MUX2X1 U628 ( .B(n474), .A(n471), .S(n1182), .Y(n485) );
  MUX2X1 U629 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1205), .Y(n479) );
  MUX2X1 U630 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1202), .Y(n478) );
  MUX2X1 U631 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1204), .Y(n482) );
  MUX2X1 U632 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1205), .Y(n481) );
  MUX2X1 U633 ( .B(n480), .A(n477), .S(n1182), .Y(n484) );
  MUX2X1 U634 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1205), .Y(n488) );
  MUX2X1 U635 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1206), .Y(n487) );
  MUX2X1 U636 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1204), .Y(n491) );
  MUX2X1 U637 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1208), .Y(n490) );
  MUX2X1 U638 ( .B(n489), .A(n486), .S(n1182), .Y(n500) );
  MUX2X1 U639 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1204), .Y(n494) );
  MUX2X1 U640 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1204), .Y(n493) );
  MUX2X1 U641 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1206), .Y(n497) );
  MUX2X1 U642 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1214), .Y(n496) );
  MUX2X1 U643 ( .B(n495), .A(n492), .S(n1182), .Y(n499) );
  MUX2X1 U644 ( .B(n498), .A(n483), .S(n1179), .Y(n1173) );
  MUX2X1 U645 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1210), .Y(n503) );
  MUX2X1 U646 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1212), .Y(n502) );
  MUX2X1 U647 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1263), .Y(n506) );
  MUX2X1 U648 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1208), .Y(n505) );
  MUX2X1 U649 ( .B(n504), .A(n501), .S(n1182), .Y(n515) );
  MUX2X1 U650 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1211), .Y(n509) );
  MUX2X1 U651 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1204), .Y(n508) );
  MUX2X1 U652 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1203), .Y(n512) );
  MUX2X1 U653 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1205), .Y(n511) );
  MUX2X1 U654 ( .B(n510), .A(n507), .S(n1182), .Y(n514) );
  MUX2X1 U655 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1211), .Y(n518) );
  MUX2X1 U656 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1211), .Y(n517) );
  MUX2X1 U657 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1211), .Y(n521) );
  MUX2X1 U658 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1211), .Y(n520) );
  MUX2X1 U659 ( .B(n519), .A(n516), .S(n1182), .Y(n530) );
  MUX2X1 U660 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1211), .Y(n524) );
  MUX2X1 U661 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1211), .Y(n523) );
  MUX2X1 U662 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1211), .Y(n527) );
  MUX2X1 U663 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1211), .Y(n526) );
  MUX2X1 U664 ( .B(n525), .A(n522), .S(n1182), .Y(n529) );
  MUX2X1 U665 ( .B(n528), .A(n513), .S(n1179), .Y(n1174) );
  MUX2X1 U666 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1211), .Y(n533) );
  MUX2X1 U667 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1211), .Y(n532) );
  MUX2X1 U668 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1211), .Y(n536) );
  MUX2X1 U669 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1211), .Y(n535) );
  MUX2X1 U670 ( .B(n534), .A(n531), .S(n1185), .Y(n545) );
  MUX2X1 U671 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1212), .Y(n539) );
  MUX2X1 U672 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1212), .Y(n538) );
  MUX2X1 U673 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1212), .Y(n542) );
  MUX2X1 U674 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1212), .Y(n541) );
  MUX2X1 U675 ( .B(n540), .A(n537), .S(n1183), .Y(n544) );
  MUX2X1 U676 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1212), .Y(n548) );
  MUX2X1 U677 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1212), .Y(n547) );
  MUX2X1 U678 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1212), .Y(n551) );
  MUX2X1 U679 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1212), .Y(n550) );
  MUX2X1 U680 ( .B(n549), .A(n546), .S(n1182), .Y(n560) );
  MUX2X1 U681 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1212), .Y(n554) );
  MUX2X1 U682 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1212), .Y(n553) );
  MUX2X1 U683 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1212), .Y(n557) );
  MUX2X1 U684 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1212), .Y(n556) );
  MUX2X1 U685 ( .B(n555), .A(n552), .S(n1182), .Y(n559) );
  MUX2X1 U686 ( .B(n558), .A(n543), .S(n1179), .Y(n1175) );
  MUX2X1 U687 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1213), .Y(n563) );
  MUX2X1 U688 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1213), .Y(n562) );
  MUX2X1 U689 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1213), .Y(n566) );
  MUX2X1 U690 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1213), .Y(n565) );
  MUX2X1 U691 ( .B(n564), .A(n561), .S(n1185), .Y(n575) );
  MUX2X1 U692 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1213), .Y(n569) );
  MUX2X1 U693 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1213), .Y(n568) );
  MUX2X1 U694 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1213), .Y(n572) );
  MUX2X1 U695 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1213), .Y(n571) );
  MUX2X1 U696 ( .B(n570), .A(n567), .S(n1183), .Y(n574) );
  MUX2X1 U697 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1213), .Y(n578) );
  MUX2X1 U698 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1213), .Y(n577) );
  MUX2X1 U699 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1213), .Y(n581) );
  MUX2X1 U700 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1213), .Y(n580) );
  MUX2X1 U701 ( .B(n579), .A(n576), .S(n1182), .Y(n590) );
  MUX2X1 U702 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1204), .Y(n584) );
  MUX2X1 U703 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1206), .Y(n583) );
  MUX2X1 U704 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1204), .Y(n587) );
  MUX2X1 U705 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1210), .Y(n586) );
  MUX2X1 U706 ( .B(n585), .A(n582), .S(n1184), .Y(n589) );
  MUX2X1 U707 ( .B(n588), .A(n573), .S(n1179), .Y(n1176) );
  MUX2X1 U708 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1206), .Y(n593) );
  MUX2X1 U709 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1206), .Y(n592) );
  MUX2X1 U710 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1204), .Y(n596) );
  MUX2X1 U711 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1210), .Y(n595) );
  MUX2X1 U712 ( .B(n594), .A(n591), .S(n1184), .Y(n605) );
  MUX2X1 U713 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1204), .Y(n599) );
  MUX2X1 U714 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1204), .Y(n598) );
  MUX2X1 U715 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1205), .Y(n602) );
  MUX2X1 U716 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1205), .Y(n601) );
  MUX2X1 U717 ( .B(n600), .A(n597), .S(n1182), .Y(n604) );
  MUX2X1 U718 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1209), .Y(n608) );
  MUX2X1 U719 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1211), .Y(n607) );
  MUX2X1 U720 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1205), .Y(n611) );
  MUX2X1 U721 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1210), .Y(n610) );
  MUX2X1 U722 ( .B(n609), .A(n606), .S(n1183), .Y(n620) );
  MUX2X1 U723 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1204), .Y(n614) );
  MUX2X1 U724 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1209), .Y(n613) );
  MUX2X1 U725 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1204), .Y(n617) );
  MUX2X1 U726 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1209), .Y(n616) );
  MUX2X1 U727 ( .B(n615), .A(n612), .S(n1182), .Y(n619) );
  MUX2X1 U728 ( .B(n618), .A(n603), .S(n1179), .Y(n1177) );
  MUX2X1 U729 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1263), .Y(n623) );
  MUX2X1 U730 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1263), .Y(n622) );
  MUX2X1 U731 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1263), .Y(n626) );
  MUX2X1 U732 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1263), .Y(n625) );
  MUX2X1 U733 ( .B(n624), .A(n621), .S(n1182), .Y(n635) );
  MUX2X1 U734 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1214), .Y(n629) );
  MUX2X1 U735 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1214), .Y(n628) );
  MUX2X1 U736 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1214), .Y(n632) );
  MUX2X1 U737 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1214), .Y(n631) );
  MUX2X1 U738 ( .B(n630), .A(n627), .S(n1182), .Y(n634) );
  MUX2X1 U739 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1214), .Y(n638) );
  MUX2X1 U740 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1214), .Y(n637) );
  MUX2X1 U741 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1214), .Y(n641) );
  MUX2X1 U742 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1214), .Y(n640) );
  MUX2X1 U743 ( .B(n639), .A(n636), .S(n1182), .Y(n650) );
  MUX2X1 U744 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1214), .Y(n644) );
  MUX2X1 U745 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1214), .Y(n643) );
  MUX2X1 U746 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1214), .Y(n647) );
  MUX2X1 U747 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1214), .Y(n646) );
  MUX2X1 U748 ( .B(n645), .A(n642), .S(n1182), .Y(n649) );
  MUX2X1 U749 ( .B(n648), .A(n633), .S(n1269), .Y(n1178) );
  INVX1 U750 ( .A(N11), .Y(n1266) );
  INVX8 U751 ( .A(n1231), .Y(n1228) );
  INVX8 U752 ( .A(n1231), .Y(n1229) );
  INVX8 U753 ( .A(n11), .Y(n1232) );
  INVX8 U754 ( .A(n11), .Y(n1233) );
  INVX8 U755 ( .A(n13), .Y(n1234) );
  INVX8 U756 ( .A(n13), .Y(n1235) );
  INVX8 U757 ( .A(n14), .Y(n1236) );
  INVX8 U758 ( .A(n14), .Y(n1237) );
  INVX8 U759 ( .A(n15), .Y(n1238) );
  INVX8 U760 ( .A(n15), .Y(n1239) );
  INVX8 U761 ( .A(n16), .Y(n1240) );
  INVX8 U762 ( .A(n16), .Y(n1241) );
  INVX8 U763 ( .A(n17), .Y(n1242) );
  INVX8 U764 ( .A(n17), .Y(n1243) );
  INVX8 U765 ( .A(n18), .Y(n1244) );
  INVX8 U766 ( .A(n18), .Y(n1245) );
  INVX8 U767 ( .A(n19), .Y(n1246) );
  INVX8 U768 ( .A(n19), .Y(n1247) );
  INVX8 U769 ( .A(n20), .Y(n1248) );
  INVX8 U770 ( .A(n20), .Y(n1249) );
  INVX8 U771 ( .A(n21), .Y(n1250) );
  INVX8 U772 ( .A(n21), .Y(n1251) );
  INVX8 U773 ( .A(n22), .Y(n1252) );
  INVX8 U774 ( .A(n22), .Y(n1253) );
  INVX8 U775 ( .A(n23), .Y(n1254) );
  INVX8 U776 ( .A(n24), .Y(n1255) );
  INVX8 U777 ( .A(n24), .Y(n1256) );
  INVX8 U778 ( .A(n25), .Y(n1257) );
  INVX8 U779 ( .A(n25), .Y(n1258) );
  INVX8 U780 ( .A(n26), .Y(n1259) );
  INVX8 U781 ( .A(n26), .Y(n1260) );
  INVX8 U782 ( .A(n27), .Y(n1261) );
  INVX8 U783 ( .A(n27), .Y(n1262) );
  AND2X2 U784 ( .A(n5), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U785 ( .A(n9), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U786 ( .A(n9), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U787 ( .A(N29), .B(n169), .Y(\data_out<3> ) );
  AND2X2 U788 ( .A(n168), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U789 ( .A(n167), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U790 ( .A(n5), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U791 ( .A(N25), .B(n167), .Y(\data_out<7> ) );
  AND2X2 U792 ( .A(n169), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U793 ( .A(n168), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U794 ( .A(n168), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U795 ( .A(n5), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U796 ( .A(n5), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U797 ( .A(N19), .B(n9), .Y(\data_out<13> ) );
  AND2X2 U798 ( .A(n169), .B(N18), .Y(\data_out<14> ) );
  NAND2X1 U799 ( .A(\mem<31><0> ), .B(n84), .Y(n1273) );
  OAI21X1 U800 ( .A(n83), .B(n1232), .C(n1273), .Y(n2311) );
  NAND2X1 U801 ( .A(\mem<31><1> ), .B(n84), .Y(n1274) );
  OAI21X1 U802 ( .A(n1235), .B(n83), .C(n1274), .Y(n2310) );
  NAND2X1 U803 ( .A(\mem<31><2> ), .B(n84), .Y(n1275) );
  OAI21X1 U804 ( .A(n1237), .B(n83), .C(n1275), .Y(n2309) );
  NAND2X1 U805 ( .A(\mem<31><3> ), .B(n84), .Y(n1276) );
  OAI21X1 U806 ( .A(n1239), .B(n83), .C(n1276), .Y(n2308) );
  NAND2X1 U807 ( .A(\mem<31><4> ), .B(n84), .Y(n1277) );
  OAI21X1 U808 ( .A(n1241), .B(n83), .C(n1277), .Y(n2307) );
  NAND2X1 U809 ( .A(\mem<31><5> ), .B(n84), .Y(n1278) );
  OAI21X1 U810 ( .A(n1243), .B(n83), .C(n1278), .Y(n2306) );
  NAND2X1 U811 ( .A(\mem<31><6> ), .B(n84), .Y(n1279) );
  OAI21X1 U812 ( .A(n1245), .B(n83), .C(n1279), .Y(n2305) );
  NAND2X1 U813 ( .A(\mem<31><7> ), .B(n84), .Y(n1280) );
  OAI21X1 U814 ( .A(n1247), .B(n83), .C(n1280), .Y(n2304) );
  NAND2X1 U815 ( .A(\mem<31><8> ), .B(n84), .Y(n1281) );
  OAI21X1 U816 ( .A(n1249), .B(n83), .C(n1281), .Y(n2303) );
  NAND2X1 U817 ( .A(\mem<31><9> ), .B(n84), .Y(n1282) );
  OAI21X1 U818 ( .A(n1251), .B(n83), .C(n1282), .Y(n2302) );
  NAND2X1 U819 ( .A(\mem<31><10> ), .B(n84), .Y(n1283) );
  OAI21X1 U820 ( .A(n1253), .B(n83), .C(n1283), .Y(n2301) );
  NAND2X1 U821 ( .A(\mem<31><11> ), .B(n84), .Y(n1284) );
  OAI21X1 U822 ( .A(n1254), .B(n83), .C(n1284), .Y(n2300) );
  NAND2X1 U823 ( .A(\mem<31><12> ), .B(n84), .Y(n1285) );
  OAI21X1 U824 ( .A(n1255), .B(n83), .C(n1285), .Y(n2299) );
  NAND2X1 U825 ( .A(\mem<31><13> ), .B(n84), .Y(n1286) );
  OAI21X1 U826 ( .A(n1257), .B(n83), .C(n1286), .Y(n2298) );
  NAND2X1 U827 ( .A(\mem<31><14> ), .B(n84), .Y(n1287) );
  OAI21X1 U828 ( .A(n1259), .B(n83), .C(n1287), .Y(n2297) );
  NAND2X1 U829 ( .A(\mem<31><15> ), .B(n84), .Y(n1288) );
  OAI21X1 U830 ( .A(n1261), .B(n83), .C(n1288), .Y(n2296) );
  NAND2X1 U831 ( .A(\mem<30><0> ), .B(n87), .Y(n1289) );
  OAI21X1 U832 ( .A(n86), .B(n1232), .C(n1289), .Y(n2295) );
  NAND2X1 U833 ( .A(\mem<30><1> ), .B(n87), .Y(n1290) );
  OAI21X1 U834 ( .A(n86), .B(n1235), .C(n1290), .Y(n2294) );
  NAND2X1 U835 ( .A(\mem<30><2> ), .B(n87), .Y(n1291) );
  OAI21X1 U836 ( .A(n86), .B(n1237), .C(n1291), .Y(n2293) );
  NAND2X1 U837 ( .A(\mem<30><3> ), .B(n87), .Y(n1292) );
  OAI21X1 U838 ( .A(n86), .B(n1239), .C(n1292), .Y(n2292) );
  NAND2X1 U839 ( .A(\mem<30><4> ), .B(n87), .Y(n1293) );
  OAI21X1 U840 ( .A(n86), .B(n1241), .C(n1293), .Y(n2291) );
  NAND2X1 U841 ( .A(\mem<30><5> ), .B(n87), .Y(n1294) );
  OAI21X1 U842 ( .A(n86), .B(n1243), .C(n1294), .Y(n2290) );
  NAND2X1 U843 ( .A(\mem<30><6> ), .B(n87), .Y(n1295) );
  OAI21X1 U844 ( .A(n86), .B(n1245), .C(n1295), .Y(n2289) );
  NAND2X1 U845 ( .A(\mem<30><7> ), .B(n87), .Y(n1296) );
  OAI21X1 U846 ( .A(n86), .B(n1247), .C(n1296), .Y(n2288) );
  NAND2X1 U847 ( .A(\mem<30><8> ), .B(n87), .Y(n1297) );
  OAI21X1 U848 ( .A(n86), .B(n1248), .C(n1297), .Y(n2287) );
  NAND2X1 U849 ( .A(\mem<30><9> ), .B(n87), .Y(n1298) );
  OAI21X1 U850 ( .A(n86), .B(n1250), .C(n1298), .Y(n2286) );
  NAND2X1 U851 ( .A(\mem<30><10> ), .B(n87), .Y(n1299) );
  OAI21X1 U852 ( .A(n86), .B(n1252), .C(n1299), .Y(n2285) );
  NAND2X1 U853 ( .A(\mem<30><11> ), .B(n87), .Y(n1300) );
  OAI21X1 U854 ( .A(n86), .B(n1254), .C(n1300), .Y(n2284) );
  NAND2X1 U855 ( .A(\mem<30><12> ), .B(n87), .Y(n1301) );
  OAI21X1 U856 ( .A(n86), .B(n1256), .C(n1301), .Y(n2283) );
  NAND2X1 U857 ( .A(\mem<30><13> ), .B(n87), .Y(n1302) );
  OAI21X1 U858 ( .A(n86), .B(n1258), .C(n1302), .Y(n2282) );
  NAND2X1 U859 ( .A(\mem<30><14> ), .B(n87), .Y(n1303) );
  OAI21X1 U860 ( .A(n86), .B(n1260), .C(n1303), .Y(n2281) );
  NAND2X1 U861 ( .A(\mem<30><15> ), .B(n87), .Y(n1304) );
  OAI21X1 U862 ( .A(n86), .B(n1262), .C(n1304), .Y(n2280) );
  NAND3X1 U863 ( .A(n1263), .B(n1184), .C(n1266), .Y(n1305) );
  NAND2X1 U864 ( .A(\mem<29><0> ), .B(n90), .Y(n1306) );
  OAI21X1 U865 ( .A(n89), .B(n1232), .C(n1306), .Y(n2279) );
  NAND2X1 U866 ( .A(\mem<29><1> ), .B(n90), .Y(n1307) );
  OAI21X1 U867 ( .A(n89), .B(n1234), .C(n1307), .Y(n2278) );
  NAND2X1 U868 ( .A(\mem<29><2> ), .B(n90), .Y(n1308) );
  OAI21X1 U869 ( .A(n89), .B(n1236), .C(n1308), .Y(n2277) );
  NAND2X1 U870 ( .A(\mem<29><3> ), .B(n90), .Y(n1309) );
  OAI21X1 U871 ( .A(n89), .B(n1238), .C(n1309), .Y(n2276) );
  NAND2X1 U872 ( .A(\mem<29><4> ), .B(n90), .Y(n1310) );
  OAI21X1 U873 ( .A(n89), .B(n1240), .C(n1310), .Y(n2275) );
  NAND2X1 U874 ( .A(\mem<29><5> ), .B(n90), .Y(n1311) );
  OAI21X1 U875 ( .A(n89), .B(n1242), .C(n1311), .Y(n2274) );
  NAND2X1 U876 ( .A(\mem<29><6> ), .B(n90), .Y(n1312) );
  OAI21X1 U877 ( .A(n89), .B(n1244), .C(n1312), .Y(n2273) );
  NAND2X1 U878 ( .A(\mem<29><7> ), .B(n90), .Y(n1313) );
  OAI21X1 U879 ( .A(n89), .B(n1246), .C(n1313), .Y(n2272) );
  NAND2X1 U880 ( .A(\mem<29><8> ), .B(n90), .Y(n1314) );
  OAI21X1 U881 ( .A(n89), .B(n1249), .C(n1314), .Y(n2271) );
  NAND2X1 U882 ( .A(\mem<29><9> ), .B(n90), .Y(n1315) );
  OAI21X1 U883 ( .A(n89), .B(n1251), .C(n1315), .Y(n2270) );
  NAND2X1 U884 ( .A(\mem<29><10> ), .B(n90), .Y(n1316) );
  OAI21X1 U885 ( .A(n89), .B(n1253), .C(n1316), .Y(n2269) );
  NAND2X1 U886 ( .A(\mem<29><11> ), .B(n90), .Y(n1317) );
  OAI21X1 U887 ( .A(n89), .B(n1254), .C(n1317), .Y(n2268) );
  NAND2X1 U888 ( .A(\mem<29><12> ), .B(n90), .Y(n1318) );
  OAI21X1 U889 ( .A(n89), .B(n1255), .C(n1318), .Y(n2267) );
  NAND2X1 U890 ( .A(\mem<29><13> ), .B(n90), .Y(n1319) );
  OAI21X1 U891 ( .A(n89), .B(n1257), .C(n1319), .Y(n2266) );
  NAND2X1 U892 ( .A(\mem<29><14> ), .B(n90), .Y(n1320) );
  OAI21X1 U893 ( .A(n89), .B(n1259), .C(n1320), .Y(n2265) );
  NAND2X1 U894 ( .A(\mem<29><15> ), .B(n90), .Y(n1321) );
  OAI21X1 U895 ( .A(n89), .B(n1261), .C(n1321), .Y(n2264) );
  NAND3X1 U896 ( .A(n1185), .B(n1266), .C(n1264), .Y(n1322) );
  NAND2X1 U897 ( .A(\mem<28><0> ), .B(n93), .Y(n1323) );
  OAI21X1 U898 ( .A(n92), .B(n1232), .C(n1323), .Y(n2263) );
  NAND2X1 U899 ( .A(\mem<28><1> ), .B(n93), .Y(n1324) );
  OAI21X1 U900 ( .A(n92), .B(n1235), .C(n1324), .Y(n2262) );
  NAND2X1 U901 ( .A(\mem<28><2> ), .B(n93), .Y(n1325) );
  OAI21X1 U902 ( .A(n92), .B(n1237), .C(n1325), .Y(n2261) );
  NAND2X1 U903 ( .A(\mem<28><3> ), .B(n93), .Y(n1326) );
  OAI21X1 U904 ( .A(n92), .B(n1239), .C(n1326), .Y(n2260) );
  NAND2X1 U905 ( .A(\mem<28><4> ), .B(n93), .Y(n1327) );
  OAI21X1 U906 ( .A(n92), .B(n1241), .C(n1327), .Y(n2259) );
  NAND2X1 U907 ( .A(\mem<28><5> ), .B(n93), .Y(n1328) );
  OAI21X1 U908 ( .A(n92), .B(n1243), .C(n1328), .Y(n2258) );
  NAND2X1 U909 ( .A(\mem<28><6> ), .B(n93), .Y(n1329) );
  OAI21X1 U910 ( .A(n92), .B(n1245), .C(n1329), .Y(n2257) );
  NAND2X1 U911 ( .A(\mem<28><7> ), .B(n93), .Y(n1330) );
  OAI21X1 U912 ( .A(n92), .B(n1247), .C(n1330), .Y(n2256) );
  NAND2X1 U913 ( .A(\mem<28><8> ), .B(n93), .Y(n1331) );
  OAI21X1 U914 ( .A(n92), .B(n1248), .C(n1331), .Y(n2255) );
  NAND2X1 U915 ( .A(\mem<28><9> ), .B(n93), .Y(n1332) );
  OAI21X1 U916 ( .A(n92), .B(n1250), .C(n1332), .Y(n2254) );
  NAND2X1 U917 ( .A(\mem<28><10> ), .B(n93), .Y(n1333) );
  OAI21X1 U918 ( .A(n92), .B(n1252), .C(n1333), .Y(n2253) );
  NAND2X1 U919 ( .A(\mem<28><11> ), .B(n93), .Y(n1334) );
  OAI21X1 U920 ( .A(n92), .B(n1254), .C(n1334), .Y(n2252) );
  NAND2X1 U921 ( .A(\mem<28><12> ), .B(n93), .Y(n1335) );
  OAI21X1 U922 ( .A(n92), .B(n1256), .C(n1335), .Y(n2251) );
  NAND2X1 U923 ( .A(\mem<28><13> ), .B(n93), .Y(n1336) );
  OAI21X1 U924 ( .A(n92), .B(n1258), .C(n1336), .Y(n2250) );
  NAND2X1 U925 ( .A(\mem<28><14> ), .B(n93), .Y(n1337) );
  OAI21X1 U926 ( .A(n92), .B(n1260), .C(n1337), .Y(n2249) );
  NAND2X1 U927 ( .A(\mem<28><15> ), .B(n93), .Y(n1338) );
  OAI21X1 U928 ( .A(n92), .B(n1262), .C(n1338), .Y(n2248) );
  NAND3X1 U929 ( .A(n1263), .B(n1265), .C(n1267), .Y(n1339) );
  NAND2X1 U930 ( .A(\mem<27><0> ), .B(n96), .Y(n1340) );
  OAI21X1 U931 ( .A(n95), .B(n1232), .C(n1340), .Y(n2247) );
  NAND2X1 U932 ( .A(\mem<27><1> ), .B(n96), .Y(n1341) );
  OAI21X1 U933 ( .A(n95), .B(n1234), .C(n1341), .Y(n2246) );
  NAND2X1 U934 ( .A(\mem<27><2> ), .B(n96), .Y(n1342) );
  OAI21X1 U935 ( .A(n95), .B(n1236), .C(n1342), .Y(n2245) );
  NAND2X1 U936 ( .A(\mem<27><3> ), .B(n96), .Y(n1343) );
  OAI21X1 U937 ( .A(n95), .B(n1238), .C(n1343), .Y(n2244) );
  NAND2X1 U938 ( .A(\mem<27><4> ), .B(n96), .Y(n1344) );
  OAI21X1 U939 ( .A(n95), .B(n1240), .C(n1344), .Y(n2243) );
  NAND2X1 U940 ( .A(\mem<27><5> ), .B(n96), .Y(n1345) );
  OAI21X1 U941 ( .A(n95), .B(n1242), .C(n1345), .Y(n2242) );
  NAND2X1 U942 ( .A(\mem<27><6> ), .B(n96), .Y(n1346) );
  OAI21X1 U943 ( .A(n95), .B(n1244), .C(n1346), .Y(n2241) );
  NAND2X1 U944 ( .A(\mem<27><7> ), .B(n96), .Y(n1347) );
  OAI21X1 U945 ( .A(n95), .B(n1246), .C(n1347), .Y(n2240) );
  NAND2X1 U946 ( .A(\mem<27><8> ), .B(n96), .Y(n1348) );
  OAI21X1 U947 ( .A(n95), .B(n1249), .C(n1348), .Y(n2239) );
  NAND2X1 U948 ( .A(\mem<27><9> ), .B(n96), .Y(n1349) );
  OAI21X1 U949 ( .A(n95), .B(n1251), .C(n1349), .Y(n2238) );
  NAND2X1 U950 ( .A(\mem<27><10> ), .B(n96), .Y(n1350) );
  OAI21X1 U951 ( .A(n95), .B(n1253), .C(n1350), .Y(n2237) );
  NAND2X1 U952 ( .A(\mem<27><11> ), .B(n96), .Y(n1351) );
  OAI21X1 U953 ( .A(n95), .B(n1254), .C(n1351), .Y(n2236) );
  NAND2X1 U954 ( .A(\mem<27><12> ), .B(n96), .Y(n1352) );
  OAI21X1 U955 ( .A(n95), .B(n1255), .C(n1352), .Y(n2235) );
  NAND2X1 U956 ( .A(\mem<27><13> ), .B(n96), .Y(n1353) );
  OAI21X1 U957 ( .A(n95), .B(n1257), .C(n1353), .Y(n2234) );
  NAND2X1 U958 ( .A(\mem<27><14> ), .B(n96), .Y(n1354) );
  OAI21X1 U959 ( .A(n95), .B(n1259), .C(n1354), .Y(n2233) );
  NAND2X1 U960 ( .A(\mem<27><15> ), .B(n96), .Y(n1355) );
  OAI21X1 U961 ( .A(n95), .B(n1261), .C(n1355), .Y(n2232) );
  NAND3X1 U962 ( .A(n1267), .B(n1265), .C(n1264), .Y(n1356) );
  NAND2X1 U963 ( .A(\mem<26><0> ), .B(n99), .Y(n1357) );
  OAI21X1 U964 ( .A(n98), .B(n1232), .C(n1357), .Y(n2231) );
  NAND2X1 U965 ( .A(\mem<26><1> ), .B(n99), .Y(n1358) );
  OAI21X1 U966 ( .A(n98), .B(n1235), .C(n1358), .Y(n2230) );
  NAND2X1 U967 ( .A(\mem<26><2> ), .B(n99), .Y(n1359) );
  OAI21X1 U968 ( .A(n98), .B(n1237), .C(n1359), .Y(n2229) );
  NAND2X1 U969 ( .A(\mem<26><3> ), .B(n99), .Y(n1360) );
  OAI21X1 U970 ( .A(n98), .B(n1239), .C(n1360), .Y(n2228) );
  NAND2X1 U971 ( .A(\mem<26><4> ), .B(n99), .Y(n1361) );
  OAI21X1 U972 ( .A(n98), .B(n1241), .C(n1361), .Y(n2227) );
  NAND2X1 U973 ( .A(\mem<26><5> ), .B(n99), .Y(n1362) );
  OAI21X1 U974 ( .A(n98), .B(n1243), .C(n1362), .Y(n2226) );
  NAND2X1 U975 ( .A(\mem<26><6> ), .B(n99), .Y(n1363) );
  OAI21X1 U976 ( .A(n98), .B(n1245), .C(n1363), .Y(n2225) );
  NAND2X1 U977 ( .A(\mem<26><7> ), .B(n99), .Y(n1364) );
  OAI21X1 U978 ( .A(n98), .B(n1247), .C(n1364), .Y(n2224) );
  NAND2X1 U979 ( .A(\mem<26><8> ), .B(n99), .Y(n1365) );
  OAI21X1 U980 ( .A(n98), .B(n1248), .C(n1365), .Y(n2223) );
  NAND2X1 U981 ( .A(\mem<26><9> ), .B(n99), .Y(n1366) );
  OAI21X1 U982 ( .A(n98), .B(n1250), .C(n1366), .Y(n2222) );
  NAND2X1 U983 ( .A(\mem<26><10> ), .B(n99), .Y(n1367) );
  OAI21X1 U984 ( .A(n98), .B(n1252), .C(n1367), .Y(n2221) );
  NAND2X1 U985 ( .A(\mem<26><11> ), .B(n99), .Y(n1368) );
  OAI21X1 U986 ( .A(n98), .B(n1254), .C(n1368), .Y(n2220) );
  NAND2X1 U987 ( .A(\mem<26><12> ), .B(n99), .Y(n1369) );
  OAI21X1 U988 ( .A(n98), .B(n1256), .C(n1369), .Y(n2219) );
  NAND2X1 U989 ( .A(\mem<26><13> ), .B(n99), .Y(n1370) );
  OAI21X1 U990 ( .A(n98), .B(n1258), .C(n1370), .Y(n2218) );
  NAND2X1 U991 ( .A(\mem<26><14> ), .B(n99), .Y(n1371) );
  OAI21X1 U992 ( .A(n98), .B(n1260), .C(n1371), .Y(n2217) );
  NAND2X1 U993 ( .A(\mem<26><15> ), .B(n99), .Y(n1372) );
  OAI21X1 U994 ( .A(n98), .B(n1262), .C(n1372), .Y(n2216) );
  NAND3X1 U995 ( .A(n1263), .B(n1267), .C(n1266), .Y(n1373) );
  NAND2X1 U996 ( .A(\mem<25><0> ), .B(n102), .Y(n1374) );
  OAI21X1 U997 ( .A(n101), .B(n1232), .C(n1374), .Y(n2215) );
  NAND2X1 U998 ( .A(\mem<25><1> ), .B(n102), .Y(n1375) );
  OAI21X1 U999 ( .A(n101), .B(n1234), .C(n1375), .Y(n2214) );
  NAND2X1 U1000 ( .A(\mem<25><2> ), .B(n102), .Y(n1376) );
  OAI21X1 U1001 ( .A(n101), .B(n1236), .C(n1376), .Y(n2213) );
  NAND2X1 U1002 ( .A(\mem<25><3> ), .B(n102), .Y(n1377) );
  OAI21X1 U1003 ( .A(n101), .B(n1238), .C(n1377), .Y(n2212) );
  NAND2X1 U1004 ( .A(\mem<25><4> ), .B(n102), .Y(n1378) );
  OAI21X1 U1005 ( .A(n101), .B(n1240), .C(n1378), .Y(n2211) );
  NAND2X1 U1006 ( .A(\mem<25><5> ), .B(n102), .Y(n1379) );
  OAI21X1 U1007 ( .A(n101), .B(n1242), .C(n1379), .Y(n2210) );
  NAND2X1 U1008 ( .A(\mem<25><6> ), .B(n102), .Y(n1380) );
  OAI21X1 U1009 ( .A(n101), .B(n1244), .C(n1380), .Y(n2209) );
  NAND2X1 U1010 ( .A(\mem<25><7> ), .B(n102), .Y(n1381) );
  OAI21X1 U1011 ( .A(n101), .B(n1246), .C(n1381), .Y(n2208) );
  NAND2X1 U1012 ( .A(\mem<25><8> ), .B(n102), .Y(n1382) );
  OAI21X1 U1013 ( .A(n101), .B(n1249), .C(n1382), .Y(n2207) );
  NAND2X1 U1014 ( .A(\mem<25><9> ), .B(n102), .Y(n1383) );
  OAI21X1 U1015 ( .A(n101), .B(n1251), .C(n1383), .Y(n2206) );
  NAND2X1 U1016 ( .A(\mem<25><10> ), .B(n102), .Y(n1384) );
  OAI21X1 U1017 ( .A(n101), .B(n1253), .C(n1384), .Y(n2205) );
  NAND2X1 U1018 ( .A(\mem<25><11> ), .B(n102), .Y(n1385) );
  OAI21X1 U1019 ( .A(n101), .B(n1254), .C(n1385), .Y(n2204) );
  NAND2X1 U1020 ( .A(\mem<25><12> ), .B(n102), .Y(n1386) );
  OAI21X1 U1021 ( .A(n101), .B(n1255), .C(n1386), .Y(n2203) );
  NAND2X1 U1022 ( .A(\mem<25><13> ), .B(n102), .Y(n1387) );
  OAI21X1 U1023 ( .A(n101), .B(n1257), .C(n1387), .Y(n2202) );
  NAND2X1 U1024 ( .A(\mem<25><14> ), .B(n102), .Y(n1388) );
  OAI21X1 U1025 ( .A(n101), .B(n1259), .C(n1388), .Y(n2201) );
  NAND2X1 U1026 ( .A(\mem<25><15> ), .B(n102), .Y(n1389) );
  OAI21X1 U1027 ( .A(n101), .B(n1261), .C(n1389), .Y(n2200) );
  NOR3X1 U1028 ( .A(n1263), .B(n1265), .C(n1184), .Y(n1783) );
  NAND2X1 U1029 ( .A(\mem<24><0> ), .B(n103), .Y(n1390) );
  OAI21X1 U1030 ( .A(n1216), .B(n1232), .C(n1390), .Y(n2199) );
  NAND2X1 U1031 ( .A(\mem<24><1> ), .B(n103), .Y(n1391) );
  OAI21X1 U1032 ( .A(n1216), .B(n1234), .C(n1391), .Y(n2198) );
  NAND2X1 U1033 ( .A(\mem<24><2> ), .B(n103), .Y(n1392) );
  OAI21X1 U1034 ( .A(n1216), .B(n1236), .C(n1392), .Y(n2197) );
  NAND2X1 U1035 ( .A(\mem<24><3> ), .B(n103), .Y(n1393) );
  OAI21X1 U1036 ( .A(n1216), .B(n1238), .C(n1393), .Y(n2196) );
  NAND2X1 U1037 ( .A(\mem<24><4> ), .B(n103), .Y(n1394) );
  OAI21X1 U1038 ( .A(n1216), .B(n1240), .C(n1394), .Y(n2195) );
  NAND2X1 U1039 ( .A(\mem<24><5> ), .B(n103), .Y(n1395) );
  OAI21X1 U1040 ( .A(n1216), .B(n1242), .C(n1395), .Y(n2194) );
  NAND2X1 U1041 ( .A(\mem<24><6> ), .B(n103), .Y(n1396) );
  OAI21X1 U1042 ( .A(n1216), .B(n1244), .C(n1396), .Y(n2193) );
  NAND2X1 U1043 ( .A(\mem<24><7> ), .B(n103), .Y(n1397) );
  OAI21X1 U1044 ( .A(n1216), .B(n1246), .C(n1397), .Y(n2192) );
  NAND2X1 U1045 ( .A(\mem<24><8> ), .B(n103), .Y(n1398) );
  OAI21X1 U1046 ( .A(n1216), .B(n1248), .C(n1398), .Y(n2191) );
  NAND2X1 U1047 ( .A(\mem<24><9> ), .B(n103), .Y(n1399) );
  OAI21X1 U1048 ( .A(n1216), .B(n1250), .C(n1399), .Y(n2190) );
  NAND2X1 U1049 ( .A(\mem<24><10> ), .B(n103), .Y(n1400) );
  OAI21X1 U1050 ( .A(n1216), .B(n1252), .C(n1400), .Y(n2189) );
  NAND2X1 U1051 ( .A(\mem<24><11> ), .B(n103), .Y(n1401) );
  OAI21X1 U1052 ( .A(n1216), .B(n1254), .C(n1401), .Y(n2188) );
  NAND2X1 U1053 ( .A(\mem<24><12> ), .B(n103), .Y(n1402) );
  OAI21X1 U1054 ( .A(n1216), .B(n1256), .C(n1402), .Y(n2187) );
  NAND2X1 U1055 ( .A(\mem<24><13> ), .B(n103), .Y(n1403) );
  OAI21X1 U1056 ( .A(n1216), .B(n1258), .C(n1403), .Y(n2186) );
  NAND2X1 U1057 ( .A(\mem<24><14> ), .B(n103), .Y(n1404) );
  OAI21X1 U1058 ( .A(n1216), .B(n1260), .C(n1404), .Y(n2185) );
  NAND2X1 U1059 ( .A(\mem<24><15> ), .B(n103), .Y(n1405) );
  OAI21X1 U1060 ( .A(n1216), .B(n1262), .C(n1405), .Y(n2184) );
  NAND2X1 U1061 ( .A(\mem<23><0> ), .B(n106), .Y(n1406) );
  OAI21X1 U1062 ( .A(n105), .B(n1232), .C(n1406), .Y(n2183) );
  NAND2X1 U1063 ( .A(\mem<23><1> ), .B(n106), .Y(n1407) );
  OAI21X1 U1064 ( .A(n105), .B(n1235), .C(n1407), .Y(n2182) );
  NAND2X1 U1065 ( .A(\mem<23><2> ), .B(n106), .Y(n1408) );
  OAI21X1 U1066 ( .A(n105), .B(n1237), .C(n1408), .Y(n2181) );
  NAND2X1 U1067 ( .A(\mem<23><3> ), .B(n106), .Y(n1409) );
  OAI21X1 U1068 ( .A(n105), .B(n1239), .C(n1409), .Y(n2180) );
  NAND2X1 U1069 ( .A(\mem<23><4> ), .B(n106), .Y(n1410) );
  OAI21X1 U1070 ( .A(n105), .B(n1241), .C(n1410), .Y(n2179) );
  NAND2X1 U1071 ( .A(\mem<23><5> ), .B(n106), .Y(n1411) );
  OAI21X1 U1072 ( .A(n105), .B(n1243), .C(n1411), .Y(n2178) );
  NAND2X1 U1073 ( .A(\mem<23><6> ), .B(n106), .Y(n1412) );
  OAI21X1 U1074 ( .A(n105), .B(n1245), .C(n1412), .Y(n2177) );
  NAND2X1 U1075 ( .A(\mem<23><7> ), .B(n106), .Y(n1413) );
  OAI21X1 U1076 ( .A(n105), .B(n1247), .C(n1413), .Y(n2176) );
  NAND2X1 U1077 ( .A(\mem<23><8> ), .B(n106), .Y(n1414) );
  OAI21X1 U1078 ( .A(n105), .B(n1249), .C(n1414), .Y(n2175) );
  NAND2X1 U1079 ( .A(\mem<23><9> ), .B(n106), .Y(n1415) );
  OAI21X1 U1080 ( .A(n105), .B(n1251), .C(n1415), .Y(n2174) );
  NAND2X1 U1081 ( .A(\mem<23><10> ), .B(n106), .Y(n1416) );
  OAI21X1 U1082 ( .A(n105), .B(n1253), .C(n1416), .Y(n2173) );
  NAND2X1 U1083 ( .A(\mem<23><11> ), .B(n106), .Y(n1417) );
  OAI21X1 U1084 ( .A(n105), .B(n1254), .C(n1417), .Y(n2172) );
  NAND2X1 U1085 ( .A(\mem<23><12> ), .B(n106), .Y(n1418) );
  OAI21X1 U1086 ( .A(n105), .B(n1256), .C(n1418), .Y(n2171) );
  NAND2X1 U1087 ( .A(\mem<23><13> ), .B(n106), .Y(n1419) );
  OAI21X1 U1088 ( .A(n105), .B(n1258), .C(n1419), .Y(n2170) );
  NAND2X1 U1089 ( .A(\mem<23><14> ), .B(n106), .Y(n1420) );
  OAI21X1 U1090 ( .A(n105), .B(n1260), .C(n1420), .Y(n2169) );
  NAND2X1 U1091 ( .A(\mem<23><15> ), .B(n106), .Y(n1421) );
  OAI21X1 U1092 ( .A(n105), .B(n1262), .C(n1421), .Y(n2168) );
  NAND2X1 U1093 ( .A(\mem<22><0> ), .B(n109), .Y(n1422) );
  OAI21X1 U1094 ( .A(n108), .B(n1232), .C(n1422), .Y(n2167) );
  NAND2X1 U1095 ( .A(\mem<22><1> ), .B(n109), .Y(n1423) );
  OAI21X1 U1096 ( .A(n108), .B(n1235), .C(n1423), .Y(n2166) );
  NAND2X1 U1097 ( .A(\mem<22><2> ), .B(n109), .Y(n1424) );
  OAI21X1 U1098 ( .A(n108), .B(n1237), .C(n1424), .Y(n2165) );
  NAND2X1 U1099 ( .A(\mem<22><3> ), .B(n109), .Y(n1425) );
  OAI21X1 U1100 ( .A(n108), .B(n1239), .C(n1425), .Y(n2164) );
  NAND2X1 U1101 ( .A(\mem<22><4> ), .B(n109), .Y(n1426) );
  OAI21X1 U1102 ( .A(n108), .B(n1241), .C(n1426), .Y(n2163) );
  NAND2X1 U1103 ( .A(\mem<22><5> ), .B(n109), .Y(n1427) );
  OAI21X1 U1104 ( .A(n108), .B(n1243), .C(n1427), .Y(n2162) );
  NAND2X1 U1105 ( .A(\mem<22><6> ), .B(n109), .Y(n1428) );
  OAI21X1 U1106 ( .A(n108), .B(n1245), .C(n1428), .Y(n2161) );
  NAND2X1 U1107 ( .A(\mem<22><7> ), .B(n109), .Y(n1429) );
  OAI21X1 U1108 ( .A(n108), .B(n1247), .C(n1429), .Y(n2160) );
  NAND2X1 U1109 ( .A(\mem<22><8> ), .B(n109), .Y(n1430) );
  OAI21X1 U1110 ( .A(n108), .B(n1249), .C(n1430), .Y(n2159) );
  NAND2X1 U1111 ( .A(\mem<22><9> ), .B(n109), .Y(n1431) );
  OAI21X1 U1112 ( .A(n108), .B(n1251), .C(n1431), .Y(n2158) );
  NAND2X1 U1113 ( .A(\mem<22><10> ), .B(n109), .Y(n1432) );
  OAI21X1 U1114 ( .A(n108), .B(n1253), .C(n1432), .Y(n2157) );
  NAND2X1 U1115 ( .A(\mem<22><11> ), .B(n109), .Y(n1433) );
  OAI21X1 U1116 ( .A(n108), .B(n1254), .C(n1433), .Y(n2156) );
  NAND2X1 U1117 ( .A(\mem<22><12> ), .B(n109), .Y(n1434) );
  OAI21X1 U1118 ( .A(n108), .B(n1256), .C(n1434), .Y(n2155) );
  NAND2X1 U1119 ( .A(\mem<22><13> ), .B(n109), .Y(n1435) );
  OAI21X1 U1120 ( .A(n108), .B(n1258), .C(n1435), .Y(n2154) );
  NAND2X1 U1121 ( .A(\mem<22><14> ), .B(n109), .Y(n1436) );
  OAI21X1 U1122 ( .A(n108), .B(n1260), .C(n1436), .Y(n2153) );
  NAND2X1 U1123 ( .A(\mem<22><15> ), .B(n109), .Y(n1437) );
  OAI21X1 U1124 ( .A(n108), .B(n1262), .C(n1437), .Y(n2152) );
  NAND2X1 U1125 ( .A(\mem<21><0> ), .B(n112), .Y(n1438) );
  OAI21X1 U1126 ( .A(n111), .B(n1232), .C(n1438), .Y(n2151) );
  NAND2X1 U1127 ( .A(\mem<21><1> ), .B(n112), .Y(n1439) );
  OAI21X1 U1128 ( .A(n111), .B(n1235), .C(n1439), .Y(n2150) );
  NAND2X1 U1129 ( .A(\mem<21><2> ), .B(n112), .Y(n1440) );
  OAI21X1 U1130 ( .A(n111), .B(n1237), .C(n1440), .Y(n2149) );
  NAND2X1 U1131 ( .A(\mem<21><3> ), .B(n112), .Y(n1441) );
  OAI21X1 U1132 ( .A(n111), .B(n1239), .C(n1441), .Y(n2148) );
  NAND2X1 U1133 ( .A(\mem<21><4> ), .B(n112), .Y(n1442) );
  OAI21X1 U1134 ( .A(n111), .B(n1241), .C(n1442), .Y(n2147) );
  NAND2X1 U1135 ( .A(\mem<21><5> ), .B(n112), .Y(n1443) );
  OAI21X1 U1136 ( .A(n111), .B(n1243), .C(n1443), .Y(n2146) );
  NAND2X1 U1137 ( .A(\mem<21><6> ), .B(n112), .Y(n1444) );
  OAI21X1 U1138 ( .A(n111), .B(n1245), .C(n1444), .Y(n2145) );
  NAND2X1 U1139 ( .A(\mem<21><7> ), .B(n112), .Y(n1445) );
  OAI21X1 U1140 ( .A(n111), .B(n1247), .C(n1445), .Y(n2144) );
  NAND2X1 U1141 ( .A(\mem<21><8> ), .B(n112), .Y(n1446) );
  OAI21X1 U1142 ( .A(n111), .B(n1249), .C(n1446), .Y(n2143) );
  NAND2X1 U1143 ( .A(\mem<21><9> ), .B(n112), .Y(n1447) );
  OAI21X1 U1144 ( .A(n111), .B(n1251), .C(n1447), .Y(n2142) );
  NAND2X1 U1145 ( .A(\mem<21><10> ), .B(n112), .Y(n1448) );
  OAI21X1 U1146 ( .A(n111), .B(n1253), .C(n1448), .Y(n2141) );
  NAND2X1 U1147 ( .A(\mem<21><11> ), .B(n112), .Y(n1449) );
  OAI21X1 U1148 ( .A(n111), .B(n1254), .C(n1449), .Y(n2140) );
  NAND2X1 U1149 ( .A(\mem<21><12> ), .B(n112), .Y(n1450) );
  OAI21X1 U1150 ( .A(n111), .B(n1256), .C(n1450), .Y(n2139) );
  NAND2X1 U1151 ( .A(\mem<21><13> ), .B(n112), .Y(n1451) );
  OAI21X1 U1152 ( .A(n111), .B(n1258), .C(n1451), .Y(n2138) );
  NAND2X1 U1153 ( .A(\mem<21><14> ), .B(n112), .Y(n1452) );
  OAI21X1 U1154 ( .A(n111), .B(n1260), .C(n1452), .Y(n2137) );
  NAND2X1 U1155 ( .A(\mem<21><15> ), .B(n112), .Y(n1453) );
  OAI21X1 U1156 ( .A(n111), .B(n1262), .C(n1453), .Y(n2136) );
  NAND2X1 U1157 ( .A(\mem<20><0> ), .B(n115), .Y(n1454) );
  OAI21X1 U1158 ( .A(n114), .B(n1232), .C(n1454), .Y(n2135) );
  NAND2X1 U1159 ( .A(\mem<20><1> ), .B(n115), .Y(n1455) );
  OAI21X1 U1160 ( .A(n114), .B(n1235), .C(n1455), .Y(n2134) );
  NAND2X1 U1161 ( .A(\mem<20><2> ), .B(n115), .Y(n1456) );
  OAI21X1 U1162 ( .A(n114), .B(n1237), .C(n1456), .Y(n2133) );
  NAND2X1 U1163 ( .A(\mem<20><3> ), .B(n115), .Y(n1457) );
  OAI21X1 U1164 ( .A(n114), .B(n1239), .C(n1457), .Y(n2132) );
  NAND2X1 U1165 ( .A(\mem<20><4> ), .B(n115), .Y(n1458) );
  OAI21X1 U1166 ( .A(n114), .B(n1241), .C(n1458), .Y(n2131) );
  NAND2X1 U1167 ( .A(\mem<20><5> ), .B(n115), .Y(n1459) );
  OAI21X1 U1168 ( .A(n114), .B(n1243), .C(n1459), .Y(n2130) );
  NAND2X1 U1169 ( .A(\mem<20><6> ), .B(n115), .Y(n1460) );
  OAI21X1 U1170 ( .A(n114), .B(n1245), .C(n1460), .Y(n2129) );
  NAND2X1 U1171 ( .A(\mem<20><7> ), .B(n115), .Y(n1461) );
  OAI21X1 U1172 ( .A(n114), .B(n1247), .C(n1461), .Y(n2128) );
  NAND2X1 U1173 ( .A(\mem<20><8> ), .B(n115), .Y(n1462) );
  OAI21X1 U1174 ( .A(n114), .B(n1249), .C(n1462), .Y(n2127) );
  NAND2X1 U1175 ( .A(\mem<20><9> ), .B(n115), .Y(n1463) );
  OAI21X1 U1177 ( .A(n114), .B(n1251), .C(n1463), .Y(n2126) );
  NAND2X1 U1178 ( .A(\mem<20><10> ), .B(n115), .Y(n1464) );
  OAI21X1 U1179 ( .A(n114), .B(n1253), .C(n1464), .Y(n2125) );
  NAND2X1 U1180 ( .A(\mem<20><11> ), .B(n115), .Y(n1465) );
  OAI21X1 U1181 ( .A(n114), .B(n1254), .C(n1465), .Y(n2124) );
  NAND2X1 U1182 ( .A(\mem<20><12> ), .B(n115), .Y(n1466) );
  OAI21X1 U1183 ( .A(n114), .B(n1256), .C(n1466), .Y(n2123) );
  NAND2X1 U1184 ( .A(\mem<20><13> ), .B(n115), .Y(n1467) );
  OAI21X1 U1185 ( .A(n114), .B(n1258), .C(n1467), .Y(n2122) );
  NAND2X1 U1186 ( .A(\mem<20><14> ), .B(n115), .Y(n1468) );
  OAI21X1 U1187 ( .A(n114), .B(n1260), .C(n1468), .Y(n2121) );
  NAND2X1 U1188 ( .A(\mem<20><15> ), .B(n115), .Y(n1469) );
  OAI21X1 U1189 ( .A(n114), .B(n1262), .C(n1469), .Y(n2120) );
  NAND2X1 U1190 ( .A(\mem<19><0> ), .B(n1217), .Y(n1470) );
  OAI21X1 U1191 ( .A(n117), .B(n1233), .C(n1470), .Y(n2119) );
  NAND2X1 U1192 ( .A(\mem<19><1> ), .B(n2), .Y(n1471) );
  OAI21X1 U1193 ( .A(n117), .B(n1235), .C(n1471), .Y(n2118) );
  NAND2X1 U1194 ( .A(\mem<19><2> ), .B(n1218), .Y(n1472) );
  OAI21X1 U1195 ( .A(n117), .B(n1237), .C(n1472), .Y(n2117) );
  NAND2X1 U1196 ( .A(\mem<19><3> ), .B(n1217), .Y(n1473) );
  OAI21X1 U1197 ( .A(n117), .B(n1239), .C(n1473), .Y(n2116) );
  NAND2X1 U1198 ( .A(\mem<19><4> ), .B(n2), .Y(n1474) );
  OAI21X1 U1199 ( .A(n117), .B(n1241), .C(n1474), .Y(n2115) );
  NAND2X1 U1200 ( .A(\mem<19><5> ), .B(n1218), .Y(n1475) );
  OAI21X1 U1201 ( .A(n117), .B(n1243), .C(n1475), .Y(n2114) );
  NAND2X1 U1202 ( .A(\mem<19><6> ), .B(n1217), .Y(n1476) );
  OAI21X1 U1203 ( .A(n117), .B(n1245), .C(n1476), .Y(n2113) );
  NAND2X1 U1204 ( .A(\mem<19><7> ), .B(n2), .Y(n1477) );
  OAI21X1 U1205 ( .A(n117), .B(n1247), .C(n1477), .Y(n2112) );
  NAND2X1 U1206 ( .A(\mem<19><8> ), .B(n1218), .Y(n1478) );
  OAI21X1 U1207 ( .A(n117), .B(n1249), .C(n1478), .Y(n2111) );
  NAND2X1 U1208 ( .A(\mem<19><9> ), .B(n1217), .Y(n1479) );
  OAI21X1 U1209 ( .A(n117), .B(n1251), .C(n1479), .Y(n2110) );
  NAND2X1 U1210 ( .A(\mem<19><10> ), .B(n2), .Y(n1480) );
  OAI21X1 U1211 ( .A(n117), .B(n1253), .C(n1480), .Y(n2109) );
  NAND2X1 U1212 ( .A(\mem<19><11> ), .B(n1218), .Y(n1481) );
  OAI21X1 U1213 ( .A(n117), .B(n1254), .C(n1481), .Y(n2108) );
  NAND2X1 U1214 ( .A(\mem<19><12> ), .B(n1217), .Y(n1482) );
  OAI21X1 U1215 ( .A(n117), .B(n1256), .C(n1482), .Y(n2107) );
  NAND2X1 U1216 ( .A(\mem<19><13> ), .B(n2), .Y(n1483) );
  OAI21X1 U1217 ( .A(n117), .B(n1258), .C(n1483), .Y(n2106) );
  NAND2X1 U1218 ( .A(\mem<19><14> ), .B(n1218), .Y(n1484) );
  OAI21X1 U1219 ( .A(n117), .B(n1260), .C(n1484), .Y(n2105) );
  NAND2X1 U1220 ( .A(\mem<19><15> ), .B(n1217), .Y(n1485) );
  OAI21X1 U1221 ( .A(n117), .B(n1262), .C(n1485), .Y(n2104) );
  NAND2X1 U1222 ( .A(\mem<18><0> ), .B(n120), .Y(n1486) );
  OAI21X1 U1223 ( .A(n119), .B(n1233), .C(n1486), .Y(n2103) );
  NAND2X1 U1224 ( .A(\mem<18><1> ), .B(n120), .Y(n1487) );
  OAI21X1 U1225 ( .A(n119), .B(n1235), .C(n1487), .Y(n2102) );
  NAND2X1 U1226 ( .A(\mem<18><2> ), .B(n120), .Y(n1488) );
  OAI21X1 U1227 ( .A(n119), .B(n1237), .C(n1488), .Y(n2101) );
  NAND2X1 U1228 ( .A(\mem<18><3> ), .B(n120), .Y(n1489) );
  OAI21X1 U1229 ( .A(n119), .B(n1239), .C(n1489), .Y(n2100) );
  NAND2X1 U1230 ( .A(\mem<18><4> ), .B(n120), .Y(n1490) );
  OAI21X1 U1231 ( .A(n119), .B(n1241), .C(n1490), .Y(n2099) );
  NAND2X1 U1232 ( .A(\mem<18><5> ), .B(n120), .Y(n1491) );
  OAI21X1 U1233 ( .A(n119), .B(n1243), .C(n1491), .Y(n2098) );
  NAND2X1 U1234 ( .A(\mem<18><6> ), .B(n120), .Y(n1492) );
  OAI21X1 U1235 ( .A(n119), .B(n1245), .C(n1492), .Y(n2097) );
  NAND2X1 U1236 ( .A(\mem<18><7> ), .B(n120), .Y(n1493) );
  OAI21X1 U1237 ( .A(n119), .B(n1247), .C(n1493), .Y(n2096) );
  NAND2X1 U1238 ( .A(\mem<18><8> ), .B(n120), .Y(n1494) );
  OAI21X1 U1239 ( .A(n119), .B(n1249), .C(n1494), .Y(n2095) );
  NAND2X1 U1240 ( .A(\mem<18><9> ), .B(n120), .Y(n1495) );
  OAI21X1 U1241 ( .A(n119), .B(n1251), .C(n1495), .Y(n2094) );
  NAND2X1 U1242 ( .A(\mem<18><10> ), .B(n120), .Y(n1496) );
  OAI21X1 U1243 ( .A(n119), .B(n1253), .C(n1496), .Y(n2093) );
  NAND2X1 U1244 ( .A(\mem<18><11> ), .B(n120), .Y(n1497) );
  OAI21X1 U1245 ( .A(n119), .B(n1254), .C(n1497), .Y(n2092) );
  NAND2X1 U1246 ( .A(\mem<18><12> ), .B(n120), .Y(n1498) );
  OAI21X1 U1247 ( .A(n119), .B(n1256), .C(n1498), .Y(n2091) );
  NAND2X1 U1248 ( .A(\mem<18><13> ), .B(n120), .Y(n1499) );
  OAI21X1 U1249 ( .A(n119), .B(n1258), .C(n1499), .Y(n2090) );
  NAND2X1 U1250 ( .A(\mem<18><14> ), .B(n120), .Y(n1500) );
  OAI21X1 U1251 ( .A(n119), .B(n1260), .C(n1500), .Y(n2089) );
  NAND2X1 U1252 ( .A(\mem<18><15> ), .B(n120), .Y(n1501) );
  OAI21X1 U1253 ( .A(n119), .B(n1262), .C(n1501), .Y(n2088) );
  NAND2X1 U1254 ( .A(\mem<17><0> ), .B(n123), .Y(n1502) );
  OAI21X1 U1255 ( .A(n122), .B(n1233), .C(n1502), .Y(n2087) );
  NAND2X1 U1256 ( .A(\mem<17><1> ), .B(n123), .Y(n1503) );
  OAI21X1 U1257 ( .A(n122), .B(n1235), .C(n1503), .Y(n2086) );
  NAND2X1 U1258 ( .A(\mem<17><2> ), .B(n123), .Y(n1504) );
  OAI21X1 U1259 ( .A(n122), .B(n1237), .C(n1504), .Y(n2085) );
  NAND2X1 U1260 ( .A(\mem<17><3> ), .B(n123), .Y(n1505) );
  OAI21X1 U1261 ( .A(n122), .B(n1239), .C(n1505), .Y(n2084) );
  NAND2X1 U1262 ( .A(\mem<17><4> ), .B(n123), .Y(n1506) );
  OAI21X1 U1263 ( .A(n122), .B(n1241), .C(n1506), .Y(n2083) );
  NAND2X1 U1264 ( .A(\mem<17><5> ), .B(n123), .Y(n1507) );
  OAI21X1 U1265 ( .A(n122), .B(n1243), .C(n1507), .Y(n2082) );
  NAND2X1 U1266 ( .A(\mem<17><6> ), .B(n123), .Y(n1508) );
  OAI21X1 U1267 ( .A(n122), .B(n1245), .C(n1508), .Y(n2081) );
  NAND2X1 U1268 ( .A(\mem<17><7> ), .B(n123), .Y(n1509) );
  OAI21X1 U1269 ( .A(n122), .B(n1247), .C(n1509), .Y(n2080) );
  NAND2X1 U1270 ( .A(\mem<17><8> ), .B(n123), .Y(n1510) );
  OAI21X1 U1271 ( .A(n122), .B(n1249), .C(n1510), .Y(n2079) );
  NAND2X1 U1272 ( .A(\mem<17><9> ), .B(n123), .Y(n1511) );
  OAI21X1 U1273 ( .A(n122), .B(n1251), .C(n1511), .Y(n2078) );
  NAND2X1 U1274 ( .A(\mem<17><10> ), .B(n123), .Y(n1512) );
  OAI21X1 U1275 ( .A(n122), .B(n1253), .C(n1512), .Y(n2077) );
  NAND2X1 U1276 ( .A(\mem<17><11> ), .B(n123), .Y(n1513) );
  OAI21X1 U1277 ( .A(n122), .B(n1254), .C(n1513), .Y(n2076) );
  NAND2X1 U1278 ( .A(\mem<17><12> ), .B(n123), .Y(n1514) );
  OAI21X1 U1279 ( .A(n122), .B(n1256), .C(n1514), .Y(n2075) );
  NAND2X1 U1280 ( .A(\mem<17><13> ), .B(n123), .Y(n1515) );
  OAI21X1 U1281 ( .A(n122), .B(n1258), .C(n1515), .Y(n2074) );
  NAND2X1 U1282 ( .A(\mem<17><14> ), .B(n123), .Y(n1516) );
  OAI21X1 U1283 ( .A(n122), .B(n1260), .C(n1516), .Y(n2073) );
  NAND2X1 U1284 ( .A(\mem<17><15> ), .B(n123), .Y(n1517) );
  OAI21X1 U1285 ( .A(n122), .B(n1262), .C(n1517), .Y(n2072) );
  NAND2X1 U1286 ( .A(\mem<16><0> ), .B(n124), .Y(n1518) );
  OAI21X1 U1287 ( .A(n1219), .B(n1233), .C(n1518), .Y(n2071) );
  NAND2X1 U1288 ( .A(\mem<16><1> ), .B(n124), .Y(n1519) );
  OAI21X1 U1289 ( .A(n1219), .B(n1235), .C(n1519), .Y(n2070) );
  NAND2X1 U1290 ( .A(\mem<16><2> ), .B(n124), .Y(n1520) );
  OAI21X1 U1291 ( .A(n1219), .B(n1237), .C(n1520), .Y(n2069) );
  NAND2X1 U1292 ( .A(\mem<16><3> ), .B(n124), .Y(n1521) );
  OAI21X1 U1293 ( .A(n1219), .B(n1239), .C(n1521), .Y(n2068) );
  NAND2X1 U1294 ( .A(\mem<16><4> ), .B(n124), .Y(n1522) );
  OAI21X1 U1295 ( .A(n1219), .B(n1241), .C(n1522), .Y(n2067) );
  NAND2X1 U1296 ( .A(\mem<16><5> ), .B(n124), .Y(n1523) );
  OAI21X1 U1297 ( .A(n1219), .B(n1243), .C(n1523), .Y(n2066) );
  NAND2X1 U1298 ( .A(\mem<16><6> ), .B(n124), .Y(n1524) );
  OAI21X1 U1299 ( .A(n1219), .B(n1245), .C(n1524), .Y(n2065) );
  NAND2X1 U1300 ( .A(\mem<16><7> ), .B(n124), .Y(n1525) );
  OAI21X1 U1301 ( .A(n1219), .B(n1247), .C(n1525), .Y(n2064) );
  NAND2X1 U1302 ( .A(\mem<16><8> ), .B(n124), .Y(n1526) );
  OAI21X1 U1303 ( .A(n1219), .B(n1249), .C(n1526), .Y(n2063) );
  NAND2X1 U1304 ( .A(\mem<16><9> ), .B(n124), .Y(n1527) );
  OAI21X1 U1305 ( .A(n1219), .B(n1251), .C(n1527), .Y(n2062) );
  NAND2X1 U1306 ( .A(\mem<16><10> ), .B(n124), .Y(n1528) );
  OAI21X1 U1307 ( .A(n1219), .B(n1253), .C(n1528), .Y(n2061) );
  NAND2X1 U1308 ( .A(\mem<16><11> ), .B(n124), .Y(n1529) );
  OAI21X1 U1309 ( .A(n1219), .B(n1254), .C(n1529), .Y(n2060) );
  NAND2X1 U1310 ( .A(\mem<16><12> ), .B(n124), .Y(n1530) );
  OAI21X1 U1311 ( .A(n1219), .B(n1256), .C(n1530), .Y(n2059) );
  NAND2X1 U1312 ( .A(\mem<16><13> ), .B(n124), .Y(n1531) );
  OAI21X1 U1313 ( .A(n1219), .B(n1258), .C(n1531), .Y(n2058) );
  NAND2X1 U1314 ( .A(\mem<16><14> ), .B(n124), .Y(n1532) );
  OAI21X1 U1315 ( .A(n1219), .B(n1260), .C(n1532), .Y(n2057) );
  NAND2X1 U1316 ( .A(\mem<16><15> ), .B(n124), .Y(n1533) );
  OAI21X1 U1317 ( .A(n1219), .B(n1262), .C(n1533), .Y(n2056) );
  NAND3X1 U1318 ( .A(n1180), .B(n2312), .C(n1270), .Y(n1534) );
  NAND2X1 U1319 ( .A(\mem<15><0> ), .B(n1220), .Y(n1535) );
  OAI21X1 U1320 ( .A(n126), .B(n1233), .C(n1535), .Y(n2055) );
  NAND2X1 U1321 ( .A(\mem<15><1> ), .B(n1), .Y(n1536) );
  OAI21X1 U1322 ( .A(n126), .B(n1235), .C(n1536), .Y(n2054) );
  NAND2X1 U1323 ( .A(\mem<15><2> ), .B(n1221), .Y(n1537) );
  OAI21X1 U1324 ( .A(n126), .B(n1237), .C(n1537), .Y(n2053) );
  NAND2X1 U1325 ( .A(\mem<15><3> ), .B(n1220), .Y(n1538) );
  OAI21X1 U1326 ( .A(n126), .B(n1239), .C(n1538), .Y(n2052) );
  NAND2X1 U1327 ( .A(\mem<15><4> ), .B(n1), .Y(n1539) );
  OAI21X1 U1328 ( .A(n126), .B(n1241), .C(n1539), .Y(n2051) );
  NAND2X1 U1329 ( .A(\mem<15><5> ), .B(n1221), .Y(n1540) );
  OAI21X1 U1330 ( .A(n126), .B(n1243), .C(n1540), .Y(n2050) );
  NAND2X1 U1331 ( .A(\mem<15><6> ), .B(n1220), .Y(n1541) );
  OAI21X1 U1332 ( .A(n126), .B(n1245), .C(n1541), .Y(n2049) );
  NAND2X1 U1333 ( .A(\mem<15><7> ), .B(n1), .Y(n1542) );
  OAI21X1 U1334 ( .A(n126), .B(n1247), .C(n1542), .Y(n2048) );
  NAND2X1 U1335 ( .A(\mem<15><8> ), .B(n1221), .Y(n1543) );
  OAI21X1 U1336 ( .A(n126), .B(n1249), .C(n1543), .Y(n2047) );
  NAND2X1 U1337 ( .A(\mem<15><9> ), .B(n1220), .Y(n1544) );
  OAI21X1 U1338 ( .A(n126), .B(n1251), .C(n1544), .Y(n2046) );
  NAND2X1 U1339 ( .A(\mem<15><10> ), .B(n1), .Y(n1545) );
  OAI21X1 U1340 ( .A(n126), .B(n1253), .C(n1545), .Y(n2045) );
  NAND2X1 U1341 ( .A(\mem<15><11> ), .B(n1221), .Y(n1546) );
  OAI21X1 U1342 ( .A(n126), .B(n1254), .C(n1546), .Y(n2044) );
  NAND2X1 U1343 ( .A(\mem<15><12> ), .B(n1220), .Y(n1547) );
  OAI21X1 U1344 ( .A(n126), .B(n1256), .C(n1547), .Y(n2043) );
  NAND2X1 U1345 ( .A(\mem<15><13> ), .B(n1), .Y(n1548) );
  OAI21X1 U1346 ( .A(n126), .B(n1258), .C(n1548), .Y(n2042) );
  NAND2X1 U1347 ( .A(\mem<15><14> ), .B(n1221), .Y(n1549) );
  OAI21X1 U1348 ( .A(n126), .B(n1260), .C(n1549), .Y(n2041) );
  NAND2X1 U1349 ( .A(\mem<15><15> ), .B(n1220), .Y(n1550) );
  OAI21X1 U1350 ( .A(n126), .B(n1262), .C(n1550), .Y(n2040) );
  NAND2X1 U1351 ( .A(\mem<14><0> ), .B(n129), .Y(n1551) );
  OAI21X1 U1352 ( .A(n128), .B(n1233), .C(n1551), .Y(n2039) );
  NAND2X1 U1353 ( .A(\mem<14><1> ), .B(n129), .Y(n1552) );
  OAI21X1 U1354 ( .A(n128), .B(n1235), .C(n1552), .Y(n2038) );
  NAND2X1 U1355 ( .A(\mem<14><2> ), .B(n129), .Y(n1553) );
  OAI21X1 U1356 ( .A(n128), .B(n1237), .C(n1553), .Y(n2037) );
  NAND2X1 U1357 ( .A(\mem<14><3> ), .B(n129), .Y(n1554) );
  OAI21X1 U1358 ( .A(n128), .B(n1239), .C(n1554), .Y(n2036) );
  NAND2X1 U1359 ( .A(\mem<14><4> ), .B(n129), .Y(n1555) );
  OAI21X1 U1360 ( .A(n128), .B(n1241), .C(n1555), .Y(n2035) );
  NAND2X1 U1361 ( .A(\mem<14><5> ), .B(n129), .Y(n1556) );
  OAI21X1 U1362 ( .A(n128), .B(n1243), .C(n1556), .Y(n2034) );
  NAND2X1 U1363 ( .A(\mem<14><6> ), .B(n129), .Y(n1557) );
  OAI21X1 U1364 ( .A(n128), .B(n1245), .C(n1557), .Y(n2033) );
  NAND2X1 U1365 ( .A(\mem<14><7> ), .B(n129), .Y(n1558) );
  OAI21X1 U1366 ( .A(n128), .B(n1247), .C(n1558), .Y(n2032) );
  NAND2X1 U1367 ( .A(\mem<14><8> ), .B(n129), .Y(n1559) );
  OAI21X1 U1368 ( .A(n128), .B(n1249), .C(n1559), .Y(n2031) );
  NAND2X1 U1369 ( .A(\mem<14><9> ), .B(n129), .Y(n1560) );
  OAI21X1 U1370 ( .A(n128), .B(n1251), .C(n1560), .Y(n2030) );
  NAND2X1 U1371 ( .A(\mem<14><10> ), .B(n129), .Y(n1561) );
  OAI21X1 U1372 ( .A(n128), .B(n1253), .C(n1561), .Y(n2029) );
  NAND2X1 U1373 ( .A(\mem<14><11> ), .B(n129), .Y(n1562) );
  OAI21X1 U1374 ( .A(n128), .B(n1254), .C(n1562), .Y(n2028) );
  NAND2X1 U1375 ( .A(\mem<14><12> ), .B(n129), .Y(n1563) );
  OAI21X1 U1376 ( .A(n128), .B(n1256), .C(n1563), .Y(n2027) );
  NAND2X1 U1377 ( .A(\mem<14><13> ), .B(n129), .Y(n1564) );
  OAI21X1 U1378 ( .A(n128), .B(n1258), .C(n1564), .Y(n2026) );
  NAND2X1 U1379 ( .A(\mem<14><14> ), .B(n129), .Y(n1565) );
  OAI21X1 U1380 ( .A(n128), .B(n1260), .C(n1565), .Y(n2025) );
  NAND2X1 U1381 ( .A(\mem<14><15> ), .B(n129), .Y(n1566) );
  OAI21X1 U1382 ( .A(n128), .B(n1262), .C(n1566), .Y(n2024) );
  NAND2X1 U1383 ( .A(\mem<13><0> ), .B(n132), .Y(n1567) );
  OAI21X1 U1384 ( .A(n131), .B(n1233), .C(n1567), .Y(n2023) );
  NAND2X1 U1385 ( .A(\mem<13><1> ), .B(n132), .Y(n1568) );
  OAI21X1 U1386 ( .A(n131), .B(n1235), .C(n1568), .Y(n2022) );
  NAND2X1 U1387 ( .A(\mem<13><2> ), .B(n132), .Y(n1569) );
  OAI21X1 U1388 ( .A(n131), .B(n1237), .C(n1569), .Y(n2021) );
  NAND2X1 U1389 ( .A(\mem<13><3> ), .B(n132), .Y(n1570) );
  OAI21X1 U1390 ( .A(n131), .B(n1239), .C(n1570), .Y(n2020) );
  NAND2X1 U1391 ( .A(\mem<13><4> ), .B(n132), .Y(n1571) );
  OAI21X1 U1392 ( .A(n131), .B(n1241), .C(n1571), .Y(n2019) );
  NAND2X1 U1393 ( .A(\mem<13><5> ), .B(n132), .Y(n1572) );
  OAI21X1 U1394 ( .A(n131), .B(n1243), .C(n1572), .Y(n2018) );
  NAND2X1 U1395 ( .A(\mem<13><6> ), .B(n132), .Y(n1573) );
  OAI21X1 U1396 ( .A(n131), .B(n1245), .C(n1573), .Y(n2017) );
  NAND2X1 U1397 ( .A(\mem<13><7> ), .B(n132), .Y(n1574) );
  OAI21X1 U1398 ( .A(n131), .B(n1247), .C(n1574), .Y(n2016) );
  NAND2X1 U1399 ( .A(\mem<13><8> ), .B(n132), .Y(n1575) );
  OAI21X1 U1400 ( .A(n131), .B(n1249), .C(n1575), .Y(n2015) );
  NAND2X1 U1401 ( .A(\mem<13><9> ), .B(n132), .Y(n1576) );
  OAI21X1 U1402 ( .A(n131), .B(n1251), .C(n1576), .Y(n2014) );
  NAND2X1 U1403 ( .A(\mem<13><10> ), .B(n132), .Y(n1577) );
  OAI21X1 U1404 ( .A(n131), .B(n1253), .C(n1577), .Y(n2013) );
  NAND2X1 U1405 ( .A(\mem<13><11> ), .B(n132), .Y(n1578) );
  OAI21X1 U1406 ( .A(n131), .B(n1254), .C(n1578), .Y(n2012) );
  NAND2X1 U1407 ( .A(\mem<13><12> ), .B(n132), .Y(n1579) );
  OAI21X1 U1408 ( .A(n131), .B(n1256), .C(n1579), .Y(n2011) );
  NAND2X1 U1409 ( .A(\mem<13><13> ), .B(n132), .Y(n1580) );
  OAI21X1 U1410 ( .A(n131), .B(n1258), .C(n1580), .Y(n2010) );
  NAND2X1 U1411 ( .A(\mem<13><14> ), .B(n132), .Y(n1581) );
  OAI21X1 U1412 ( .A(n131), .B(n1260), .C(n1581), .Y(n2009) );
  NAND2X1 U1413 ( .A(\mem<13><15> ), .B(n132), .Y(n1582) );
  OAI21X1 U1414 ( .A(n131), .B(n1262), .C(n1582), .Y(n2008) );
  NAND2X1 U1415 ( .A(\mem<12><0> ), .B(n135), .Y(n1583) );
  OAI21X1 U1416 ( .A(n134), .B(n1233), .C(n1583), .Y(n2007) );
  NAND2X1 U1417 ( .A(\mem<12><1> ), .B(n135), .Y(n1584) );
  OAI21X1 U1418 ( .A(n134), .B(n1235), .C(n1584), .Y(n2006) );
  NAND2X1 U1419 ( .A(\mem<12><2> ), .B(n135), .Y(n1585) );
  OAI21X1 U1420 ( .A(n134), .B(n1237), .C(n1585), .Y(n2005) );
  NAND2X1 U1421 ( .A(\mem<12><3> ), .B(n135), .Y(n1586) );
  OAI21X1 U1422 ( .A(n134), .B(n1239), .C(n1586), .Y(n2004) );
  NAND2X1 U1423 ( .A(\mem<12><4> ), .B(n135), .Y(n1587) );
  OAI21X1 U1424 ( .A(n134), .B(n1241), .C(n1587), .Y(n2003) );
  NAND2X1 U1425 ( .A(\mem<12><5> ), .B(n135), .Y(n1588) );
  OAI21X1 U1426 ( .A(n134), .B(n1243), .C(n1588), .Y(n2002) );
  NAND2X1 U1427 ( .A(\mem<12><6> ), .B(n135), .Y(n1589) );
  OAI21X1 U1428 ( .A(n134), .B(n1245), .C(n1589), .Y(n2001) );
  NAND2X1 U1429 ( .A(\mem<12><7> ), .B(n135), .Y(n1590) );
  OAI21X1 U1430 ( .A(n134), .B(n1247), .C(n1590), .Y(n2000) );
  NAND2X1 U1431 ( .A(\mem<12><8> ), .B(n135), .Y(n1591) );
  OAI21X1 U1432 ( .A(n134), .B(n1249), .C(n1591), .Y(n1999) );
  NAND2X1 U1433 ( .A(\mem<12><9> ), .B(n135), .Y(n1592) );
  OAI21X1 U1434 ( .A(n134), .B(n1251), .C(n1592), .Y(n1998) );
  NAND2X1 U1435 ( .A(\mem<12><10> ), .B(n135), .Y(n1593) );
  OAI21X1 U1436 ( .A(n134), .B(n1253), .C(n1593), .Y(n1997) );
  NAND2X1 U1437 ( .A(\mem<12><11> ), .B(n135), .Y(n1594) );
  OAI21X1 U1438 ( .A(n134), .B(n1254), .C(n1594), .Y(n1996) );
  NAND2X1 U1439 ( .A(\mem<12><12> ), .B(n135), .Y(n1595) );
  OAI21X1 U1440 ( .A(n134), .B(n1256), .C(n1595), .Y(n1995) );
  NAND2X1 U1441 ( .A(\mem<12><13> ), .B(n135), .Y(n1596) );
  OAI21X1 U1442 ( .A(n134), .B(n1258), .C(n1596), .Y(n1994) );
  NAND2X1 U1443 ( .A(\mem<12><14> ), .B(n135), .Y(n1597) );
  OAI21X1 U1444 ( .A(n134), .B(n1260), .C(n1597), .Y(n1993) );
  NAND2X1 U1445 ( .A(\mem<12><15> ), .B(n135), .Y(n1598) );
  OAI21X1 U1446 ( .A(n134), .B(n1262), .C(n1598), .Y(n1992) );
  NAND2X1 U1447 ( .A(\mem<11><0> ), .B(n138), .Y(n1599) );
  OAI21X1 U1448 ( .A(n137), .B(n1233), .C(n1599), .Y(n1991) );
  NAND2X1 U1449 ( .A(\mem<11><1> ), .B(n138), .Y(n1600) );
  OAI21X1 U1450 ( .A(n137), .B(n1234), .C(n1600), .Y(n1990) );
  NAND2X1 U1451 ( .A(\mem<11><2> ), .B(n138), .Y(n1601) );
  OAI21X1 U1452 ( .A(n137), .B(n1236), .C(n1601), .Y(n1989) );
  NAND2X1 U1453 ( .A(\mem<11><3> ), .B(n138), .Y(n1602) );
  OAI21X1 U1454 ( .A(n137), .B(n1238), .C(n1602), .Y(n1988) );
  NAND2X1 U1455 ( .A(\mem<11><4> ), .B(n138), .Y(n1603) );
  OAI21X1 U1456 ( .A(n137), .B(n1240), .C(n1603), .Y(n1987) );
  NAND2X1 U1457 ( .A(\mem<11><5> ), .B(n138), .Y(n1604) );
  OAI21X1 U1458 ( .A(n137), .B(n1242), .C(n1604), .Y(n1986) );
  NAND2X1 U1459 ( .A(\mem<11><6> ), .B(n138), .Y(n1605) );
  OAI21X1 U1460 ( .A(n137), .B(n1244), .C(n1605), .Y(n1985) );
  NAND2X1 U1461 ( .A(\mem<11><7> ), .B(n138), .Y(n1606) );
  OAI21X1 U1462 ( .A(n137), .B(n1246), .C(n1606), .Y(n1984) );
  NAND2X1 U1463 ( .A(\mem<11><8> ), .B(n138), .Y(n1607) );
  OAI21X1 U1464 ( .A(n137), .B(n1248), .C(n1607), .Y(n1983) );
  NAND2X1 U1465 ( .A(\mem<11><9> ), .B(n138), .Y(n1608) );
  OAI21X1 U1466 ( .A(n137), .B(n1250), .C(n1608), .Y(n1982) );
  NAND2X1 U1467 ( .A(\mem<11><10> ), .B(n138), .Y(n1609) );
  OAI21X1 U1468 ( .A(n137), .B(n1252), .C(n1609), .Y(n1981) );
  NAND2X1 U1469 ( .A(\mem<11><11> ), .B(n138), .Y(n1610) );
  OAI21X1 U1470 ( .A(n137), .B(n1254), .C(n1610), .Y(n1980) );
  NAND2X1 U1471 ( .A(\mem<11><12> ), .B(n138), .Y(n1611) );
  OAI21X1 U1472 ( .A(n137), .B(n1255), .C(n1611), .Y(n1979) );
  NAND2X1 U1473 ( .A(\mem<11><13> ), .B(n138), .Y(n1612) );
  OAI21X1 U1474 ( .A(n137), .B(n1257), .C(n1612), .Y(n1978) );
  NAND2X1 U1475 ( .A(\mem<11><14> ), .B(n138), .Y(n1613) );
  OAI21X1 U1476 ( .A(n137), .B(n1259), .C(n1613), .Y(n1977) );
  NAND2X1 U1477 ( .A(\mem<11><15> ), .B(n138), .Y(n1614) );
  OAI21X1 U1478 ( .A(n137), .B(n1261), .C(n1614), .Y(n1976) );
  NAND2X1 U1479 ( .A(\mem<10><0> ), .B(n141), .Y(n1615) );
  OAI21X1 U1480 ( .A(n140), .B(n1233), .C(n1615), .Y(n1975) );
  NAND2X1 U1481 ( .A(\mem<10><1> ), .B(n141), .Y(n1616) );
  OAI21X1 U1482 ( .A(n140), .B(n1234), .C(n1616), .Y(n1974) );
  NAND2X1 U1483 ( .A(\mem<10><2> ), .B(n141), .Y(n1617) );
  OAI21X1 U1484 ( .A(n140), .B(n1236), .C(n1617), .Y(n1973) );
  NAND2X1 U1485 ( .A(\mem<10><3> ), .B(n141), .Y(n1618) );
  OAI21X1 U1486 ( .A(n140), .B(n1238), .C(n1618), .Y(n1972) );
  NAND2X1 U1487 ( .A(\mem<10><4> ), .B(n141), .Y(n1619) );
  OAI21X1 U1488 ( .A(n140), .B(n1240), .C(n1619), .Y(n1971) );
  NAND2X1 U1489 ( .A(\mem<10><5> ), .B(n141), .Y(n1620) );
  OAI21X1 U1490 ( .A(n140), .B(n1242), .C(n1620), .Y(n1970) );
  NAND2X1 U1491 ( .A(\mem<10><6> ), .B(n141), .Y(n1621) );
  OAI21X1 U1492 ( .A(n140), .B(n1244), .C(n1621), .Y(n1969) );
  NAND2X1 U1493 ( .A(\mem<10><7> ), .B(n141), .Y(n1622) );
  OAI21X1 U1494 ( .A(n140), .B(n1246), .C(n1622), .Y(n1968) );
  NAND2X1 U1495 ( .A(\mem<10><8> ), .B(n141), .Y(n1623) );
  OAI21X1 U1496 ( .A(n140), .B(n1248), .C(n1623), .Y(n1967) );
  NAND2X1 U1497 ( .A(\mem<10><9> ), .B(n141), .Y(n1624) );
  OAI21X1 U1498 ( .A(n140), .B(n1250), .C(n1624), .Y(n1966) );
  NAND2X1 U1499 ( .A(\mem<10><10> ), .B(n141), .Y(n1625) );
  OAI21X1 U1500 ( .A(n140), .B(n1252), .C(n1625), .Y(n1965) );
  NAND2X1 U1501 ( .A(\mem<10><11> ), .B(n141), .Y(n1626) );
  OAI21X1 U1502 ( .A(n140), .B(n1254), .C(n1626), .Y(n1964) );
  NAND2X1 U1503 ( .A(\mem<10><12> ), .B(n141), .Y(n1627) );
  OAI21X1 U1504 ( .A(n140), .B(n1255), .C(n1627), .Y(n1963) );
  NAND2X1 U1505 ( .A(\mem<10><13> ), .B(n141), .Y(n1628) );
  OAI21X1 U1506 ( .A(n140), .B(n1257), .C(n1628), .Y(n1962) );
  NAND2X1 U1507 ( .A(\mem<10><14> ), .B(n141), .Y(n1629) );
  OAI21X1 U1508 ( .A(n140), .B(n1259), .C(n1629), .Y(n1961) );
  NAND2X1 U1509 ( .A(\mem<10><15> ), .B(n141), .Y(n1630) );
  OAI21X1 U1510 ( .A(n140), .B(n1261), .C(n1630), .Y(n1960) );
  NAND2X1 U1511 ( .A(\mem<9><0> ), .B(n144), .Y(n1631) );
  OAI21X1 U1512 ( .A(n143), .B(n1233), .C(n1631), .Y(n1959) );
  NAND2X1 U1513 ( .A(\mem<9><1> ), .B(n144), .Y(n1632) );
  OAI21X1 U1514 ( .A(n143), .B(n1234), .C(n1632), .Y(n1958) );
  NAND2X1 U1515 ( .A(\mem<9><2> ), .B(n144), .Y(n1633) );
  OAI21X1 U1516 ( .A(n143), .B(n1236), .C(n1633), .Y(n1957) );
  NAND2X1 U1517 ( .A(\mem<9><3> ), .B(n144), .Y(n1634) );
  OAI21X1 U1518 ( .A(n143), .B(n1238), .C(n1634), .Y(n1956) );
  NAND2X1 U1519 ( .A(\mem<9><4> ), .B(n144), .Y(n1635) );
  OAI21X1 U1520 ( .A(n143), .B(n1240), .C(n1635), .Y(n1955) );
  NAND2X1 U1521 ( .A(\mem<9><5> ), .B(n144), .Y(n1636) );
  OAI21X1 U1522 ( .A(n143), .B(n1242), .C(n1636), .Y(n1954) );
  NAND2X1 U1523 ( .A(\mem<9><6> ), .B(n144), .Y(n1637) );
  OAI21X1 U1524 ( .A(n143), .B(n1244), .C(n1637), .Y(n1953) );
  NAND2X1 U1525 ( .A(\mem<9><7> ), .B(n144), .Y(n1638) );
  OAI21X1 U1526 ( .A(n143), .B(n1246), .C(n1638), .Y(n1952) );
  NAND2X1 U1527 ( .A(\mem<9><8> ), .B(n144), .Y(n1639) );
  OAI21X1 U1528 ( .A(n143), .B(n1248), .C(n1639), .Y(n1951) );
  NAND2X1 U1529 ( .A(\mem<9><9> ), .B(n144), .Y(n1640) );
  OAI21X1 U1530 ( .A(n143), .B(n1250), .C(n1640), .Y(n1950) );
  NAND2X1 U1531 ( .A(\mem<9><10> ), .B(n144), .Y(n1641) );
  OAI21X1 U1532 ( .A(n143), .B(n1252), .C(n1641), .Y(n1949) );
  NAND2X1 U1533 ( .A(\mem<9><11> ), .B(n144), .Y(n1642) );
  OAI21X1 U1534 ( .A(n143), .B(n1254), .C(n1642), .Y(n1948) );
  NAND2X1 U1535 ( .A(\mem<9><12> ), .B(n144), .Y(n1643) );
  OAI21X1 U1536 ( .A(n143), .B(n1255), .C(n1643), .Y(n1947) );
  NAND2X1 U1537 ( .A(\mem<9><13> ), .B(n144), .Y(n1644) );
  OAI21X1 U1538 ( .A(n143), .B(n1257), .C(n1644), .Y(n1946) );
  NAND2X1 U1539 ( .A(\mem<9><14> ), .B(n144), .Y(n1645) );
  OAI21X1 U1540 ( .A(n143), .B(n1259), .C(n1645), .Y(n1945) );
  NAND2X1 U1541 ( .A(\mem<9><15> ), .B(n144), .Y(n1646) );
  OAI21X1 U1542 ( .A(n143), .B(n1261), .C(n1646), .Y(n1944) );
  NAND2X1 U1543 ( .A(\mem<8><0> ), .B(n1223), .Y(n1648) );
  OAI21X1 U1544 ( .A(n1222), .B(n1233), .C(n1648), .Y(n1943) );
  NAND2X1 U1545 ( .A(\mem<8><1> ), .B(n4), .Y(n1649) );
  OAI21X1 U1546 ( .A(n1222), .B(n1234), .C(n1649), .Y(n1942) );
  NAND2X1 U1547 ( .A(\mem<8><2> ), .B(n4), .Y(n1650) );
  OAI21X1 U1548 ( .A(n1222), .B(n1236), .C(n1650), .Y(n1941) );
  NAND2X1 U1549 ( .A(\mem<8><3> ), .B(n1224), .Y(n1651) );
  OAI21X1 U1550 ( .A(n1222), .B(n1238), .C(n1651), .Y(n1940) );
  NAND2X1 U1551 ( .A(\mem<8><4> ), .B(n1224), .Y(n1652) );
  OAI21X1 U1552 ( .A(n1222), .B(n1240), .C(n1652), .Y(n1939) );
  NAND2X1 U1553 ( .A(\mem<8><5> ), .B(n1223), .Y(n1653) );
  OAI21X1 U1554 ( .A(n1222), .B(n1242), .C(n1653), .Y(n1938) );
  NAND2X1 U1555 ( .A(\mem<8><6> ), .B(n1223), .Y(n1654) );
  OAI21X1 U1556 ( .A(n1222), .B(n1244), .C(n1654), .Y(n1937) );
  NAND2X1 U1557 ( .A(\mem<8><7> ), .B(n4), .Y(n1655) );
  OAI21X1 U1558 ( .A(n1222), .B(n1246), .C(n1655), .Y(n1936) );
  NAND2X1 U1559 ( .A(\mem<8><8> ), .B(n1224), .Y(n1656) );
  OAI21X1 U1560 ( .A(n1222), .B(n1248), .C(n1656), .Y(n1935) );
  NAND2X1 U1561 ( .A(\mem<8><9> ), .B(n1223), .Y(n1657) );
  OAI21X1 U1562 ( .A(n1222), .B(n1250), .C(n1657), .Y(n1934) );
  NAND2X1 U1563 ( .A(\mem<8><10> ), .B(n1223), .Y(n1658) );
  OAI21X1 U1564 ( .A(n1222), .B(n1252), .C(n1658), .Y(n1933) );
  NAND2X1 U1565 ( .A(\mem<8><11> ), .B(n4), .Y(n1659) );
  OAI21X1 U1566 ( .A(n1222), .B(n1254), .C(n1659), .Y(n1932) );
  NAND2X1 U1567 ( .A(\mem<8><12> ), .B(n4), .Y(n1660) );
  OAI21X1 U1568 ( .A(n1222), .B(n1255), .C(n1660), .Y(n1931) );
  NAND2X1 U1569 ( .A(\mem<8><13> ), .B(n1224), .Y(n1661) );
  OAI21X1 U1570 ( .A(n1222), .B(n1257), .C(n1661), .Y(n1930) );
  NAND2X1 U1571 ( .A(\mem<8><14> ), .B(n1224), .Y(n1662) );
  OAI21X1 U1572 ( .A(n1222), .B(n1259), .C(n1662), .Y(n1929) );
  NAND2X1 U1573 ( .A(\mem<8><15> ), .B(n1223), .Y(n1663) );
  OAI21X1 U1574 ( .A(n1222), .B(n1261), .C(n1663), .Y(n1928) );
  NAND3X1 U1575 ( .A(n1268), .B(n2312), .C(n1270), .Y(n1664) );
  NAND2X1 U1576 ( .A(\mem<7><0> ), .B(n147), .Y(n1665) );
  OAI21X1 U1577 ( .A(n146), .B(n1232), .C(n1665), .Y(n1927) );
  NAND2X1 U1578 ( .A(\mem<7><1> ), .B(n147), .Y(n1666) );
  OAI21X1 U1579 ( .A(n146), .B(n1234), .C(n1666), .Y(n1926) );
  NAND2X1 U1580 ( .A(\mem<7><2> ), .B(n147), .Y(n1667) );
  OAI21X1 U1581 ( .A(n146), .B(n1236), .C(n1667), .Y(n1925) );
  NAND2X1 U1582 ( .A(\mem<7><3> ), .B(n147), .Y(n1668) );
  OAI21X1 U1583 ( .A(n146), .B(n1238), .C(n1668), .Y(n1924) );
  NAND2X1 U1584 ( .A(\mem<7><4> ), .B(n147), .Y(n1669) );
  OAI21X1 U1585 ( .A(n146), .B(n1240), .C(n1669), .Y(n1923) );
  NAND2X1 U1586 ( .A(\mem<7><5> ), .B(n147), .Y(n1670) );
  OAI21X1 U1587 ( .A(n146), .B(n1242), .C(n1670), .Y(n1922) );
  NAND2X1 U1588 ( .A(\mem<7><6> ), .B(n147), .Y(n1671) );
  OAI21X1 U1589 ( .A(n146), .B(n1244), .C(n1671), .Y(n1921) );
  NAND2X1 U1590 ( .A(\mem<7><7> ), .B(n147), .Y(n1672) );
  OAI21X1 U1591 ( .A(n146), .B(n1246), .C(n1672), .Y(n1920) );
  NAND2X1 U1592 ( .A(\mem<7><8> ), .B(n147), .Y(n1673) );
  OAI21X1 U1593 ( .A(n146), .B(n1248), .C(n1673), .Y(n1919) );
  NAND2X1 U1594 ( .A(\mem<7><9> ), .B(n147), .Y(n1674) );
  OAI21X1 U1595 ( .A(n146), .B(n1250), .C(n1674), .Y(n1918) );
  NAND2X1 U1596 ( .A(\mem<7><10> ), .B(n147), .Y(n1675) );
  OAI21X1 U1597 ( .A(n146), .B(n1252), .C(n1675), .Y(n1917) );
  NAND2X1 U1598 ( .A(\mem<7><11> ), .B(n147), .Y(n1676) );
  OAI21X1 U1599 ( .A(n146), .B(n1254), .C(n1676), .Y(n1916) );
  NAND2X1 U1600 ( .A(\mem<7><12> ), .B(n147), .Y(n1677) );
  OAI21X1 U1601 ( .A(n146), .B(n1255), .C(n1677), .Y(n1915) );
  NAND2X1 U1602 ( .A(\mem<7><13> ), .B(n147), .Y(n1678) );
  OAI21X1 U1603 ( .A(n146), .B(n1257), .C(n1678), .Y(n1914) );
  NAND2X1 U1604 ( .A(\mem<7><14> ), .B(n147), .Y(n1679) );
  OAI21X1 U1605 ( .A(n146), .B(n1259), .C(n1679), .Y(n1913) );
  NAND2X1 U1606 ( .A(\mem<7><15> ), .B(n147), .Y(n1680) );
  OAI21X1 U1607 ( .A(n146), .B(n1261), .C(n1680), .Y(n1912) );
  NAND2X1 U1608 ( .A(\mem<6><0> ), .B(n150), .Y(n1681) );
  OAI21X1 U1609 ( .A(n149), .B(n1233), .C(n1681), .Y(n1911) );
  NAND2X1 U1610 ( .A(\mem<6><1> ), .B(n150), .Y(n1682) );
  OAI21X1 U1611 ( .A(n149), .B(n1234), .C(n1682), .Y(n1910) );
  NAND2X1 U1612 ( .A(\mem<6><2> ), .B(n150), .Y(n1683) );
  OAI21X1 U1613 ( .A(n149), .B(n1236), .C(n1683), .Y(n1909) );
  NAND2X1 U1614 ( .A(\mem<6><3> ), .B(n150), .Y(n1684) );
  OAI21X1 U1615 ( .A(n149), .B(n1238), .C(n1684), .Y(n1908) );
  NAND2X1 U1616 ( .A(\mem<6><4> ), .B(n150), .Y(n1685) );
  OAI21X1 U1617 ( .A(n149), .B(n1240), .C(n1685), .Y(n1907) );
  NAND2X1 U1618 ( .A(\mem<6><5> ), .B(n150), .Y(n1686) );
  OAI21X1 U1619 ( .A(n149), .B(n1242), .C(n1686), .Y(n1906) );
  NAND2X1 U1620 ( .A(\mem<6><6> ), .B(n150), .Y(n1687) );
  OAI21X1 U1621 ( .A(n149), .B(n1244), .C(n1687), .Y(n1905) );
  NAND2X1 U1622 ( .A(\mem<6><7> ), .B(n150), .Y(n1688) );
  OAI21X1 U1623 ( .A(n149), .B(n1246), .C(n1688), .Y(n1904) );
  NAND2X1 U1624 ( .A(\mem<6><8> ), .B(n150), .Y(n1689) );
  OAI21X1 U1625 ( .A(n149), .B(n1248), .C(n1689), .Y(n1903) );
  NAND2X1 U1626 ( .A(\mem<6><9> ), .B(n150), .Y(n1690) );
  OAI21X1 U1627 ( .A(n149), .B(n1250), .C(n1690), .Y(n1902) );
  NAND2X1 U1628 ( .A(\mem<6><10> ), .B(n150), .Y(n1691) );
  OAI21X1 U1629 ( .A(n149), .B(n1252), .C(n1691), .Y(n1901) );
  NAND2X1 U1630 ( .A(\mem<6><11> ), .B(n150), .Y(n1692) );
  OAI21X1 U1631 ( .A(n149), .B(n1254), .C(n1692), .Y(n1900) );
  NAND2X1 U1632 ( .A(\mem<6><12> ), .B(n150), .Y(n1693) );
  OAI21X1 U1633 ( .A(n149), .B(n1255), .C(n1693), .Y(n1899) );
  NAND2X1 U1634 ( .A(\mem<6><13> ), .B(n150), .Y(n1694) );
  OAI21X1 U1635 ( .A(n149), .B(n1257), .C(n1694), .Y(n1898) );
  NAND2X1 U1636 ( .A(\mem<6><14> ), .B(n150), .Y(n1695) );
  OAI21X1 U1637 ( .A(n149), .B(n1259), .C(n1695), .Y(n1897) );
  NAND2X1 U1638 ( .A(\mem<6><15> ), .B(n150), .Y(n1696) );
  OAI21X1 U1639 ( .A(n149), .B(n1261), .C(n1696), .Y(n1896) );
  NAND2X1 U1640 ( .A(\mem<5><0> ), .B(n153), .Y(n1698) );
  OAI21X1 U1641 ( .A(n152), .B(n1232), .C(n1698), .Y(n1895) );
  NAND2X1 U1642 ( .A(\mem<5><1> ), .B(n153), .Y(n1699) );
  OAI21X1 U1643 ( .A(n152), .B(n1234), .C(n1699), .Y(n1894) );
  NAND2X1 U1644 ( .A(\mem<5><2> ), .B(n153), .Y(n1700) );
  OAI21X1 U1645 ( .A(n152), .B(n1236), .C(n1700), .Y(n1893) );
  NAND2X1 U1646 ( .A(\mem<5><3> ), .B(n153), .Y(n1701) );
  OAI21X1 U1647 ( .A(n152), .B(n1238), .C(n1701), .Y(n1892) );
  NAND2X1 U1648 ( .A(\mem<5><4> ), .B(n153), .Y(n1702) );
  OAI21X1 U1649 ( .A(n152), .B(n1240), .C(n1702), .Y(n1891) );
  NAND2X1 U1650 ( .A(\mem<5><5> ), .B(n153), .Y(n1703) );
  OAI21X1 U1651 ( .A(n152), .B(n1242), .C(n1703), .Y(n1890) );
  NAND2X1 U1652 ( .A(\mem<5><6> ), .B(n153), .Y(n1704) );
  OAI21X1 U1653 ( .A(n152), .B(n1244), .C(n1704), .Y(n1889) );
  NAND2X1 U1654 ( .A(\mem<5><7> ), .B(n153), .Y(n1705) );
  OAI21X1 U1655 ( .A(n152), .B(n1246), .C(n1705), .Y(n1888) );
  NAND2X1 U1656 ( .A(\mem<5><8> ), .B(n153), .Y(n1706) );
  OAI21X1 U1657 ( .A(n152), .B(n1248), .C(n1706), .Y(n1887) );
  NAND2X1 U1658 ( .A(\mem<5><9> ), .B(n153), .Y(n1707) );
  OAI21X1 U1659 ( .A(n152), .B(n1250), .C(n1707), .Y(n1886) );
  NAND2X1 U1660 ( .A(\mem<5><10> ), .B(n153), .Y(n1708) );
  OAI21X1 U1661 ( .A(n152), .B(n1252), .C(n1708), .Y(n1885) );
  NAND2X1 U1662 ( .A(\mem<5><11> ), .B(n153), .Y(n1709) );
  OAI21X1 U1663 ( .A(n152), .B(n1254), .C(n1709), .Y(n1884) );
  NAND2X1 U1664 ( .A(\mem<5><12> ), .B(n153), .Y(n1710) );
  OAI21X1 U1665 ( .A(n152), .B(n1255), .C(n1710), .Y(n1883) );
  NAND2X1 U1666 ( .A(\mem<5><13> ), .B(n153), .Y(n1711) );
  OAI21X1 U1667 ( .A(n152), .B(n1257), .C(n1711), .Y(n1882) );
  NAND2X1 U1668 ( .A(\mem<5><14> ), .B(n153), .Y(n1712) );
  OAI21X1 U1669 ( .A(n152), .B(n1259), .C(n1712), .Y(n1881) );
  NAND2X1 U1670 ( .A(\mem<5><15> ), .B(n153), .Y(n1713) );
  OAI21X1 U1671 ( .A(n152), .B(n1261), .C(n1713), .Y(n1880) );
  NAND2X1 U1672 ( .A(\mem<4><0> ), .B(n156), .Y(n1715) );
  OAI21X1 U1673 ( .A(n155), .B(n1233), .C(n1715), .Y(n1879) );
  NAND2X1 U1674 ( .A(\mem<4><1> ), .B(n156), .Y(n1716) );
  OAI21X1 U1675 ( .A(n155), .B(n1234), .C(n1716), .Y(n1878) );
  NAND2X1 U1676 ( .A(\mem<4><2> ), .B(n156), .Y(n1717) );
  OAI21X1 U1677 ( .A(n155), .B(n1236), .C(n1717), .Y(n1877) );
  NAND2X1 U1678 ( .A(\mem<4><3> ), .B(n156), .Y(n1718) );
  OAI21X1 U1679 ( .A(n155), .B(n1238), .C(n1718), .Y(n1876) );
  NAND2X1 U1680 ( .A(\mem<4><4> ), .B(n156), .Y(n1719) );
  OAI21X1 U1681 ( .A(n155), .B(n1240), .C(n1719), .Y(n1875) );
  NAND2X1 U1682 ( .A(\mem<4><5> ), .B(n156), .Y(n1720) );
  OAI21X1 U1683 ( .A(n155), .B(n1242), .C(n1720), .Y(n1874) );
  NAND2X1 U1684 ( .A(\mem<4><6> ), .B(n156), .Y(n1721) );
  OAI21X1 U1685 ( .A(n155), .B(n1244), .C(n1721), .Y(n1873) );
  NAND2X1 U1686 ( .A(\mem<4><7> ), .B(n156), .Y(n1722) );
  OAI21X1 U1687 ( .A(n155), .B(n1246), .C(n1722), .Y(n1872) );
  NAND2X1 U1688 ( .A(\mem<4><8> ), .B(n156), .Y(n1723) );
  OAI21X1 U1689 ( .A(n155), .B(n1248), .C(n1723), .Y(n1871) );
  NAND2X1 U1690 ( .A(\mem<4><9> ), .B(n156), .Y(n1724) );
  OAI21X1 U1691 ( .A(n155), .B(n1250), .C(n1724), .Y(n1870) );
  NAND2X1 U1692 ( .A(\mem<4><10> ), .B(n156), .Y(n1725) );
  OAI21X1 U1693 ( .A(n155), .B(n1252), .C(n1725), .Y(n1869) );
  NAND2X1 U1694 ( .A(\mem<4><11> ), .B(n156), .Y(n1726) );
  OAI21X1 U1695 ( .A(n155), .B(n1254), .C(n1726), .Y(n1868) );
  NAND2X1 U1696 ( .A(\mem<4><12> ), .B(n156), .Y(n1727) );
  OAI21X1 U1697 ( .A(n155), .B(n1255), .C(n1727), .Y(n1867) );
  NAND2X1 U1698 ( .A(\mem<4><13> ), .B(n156), .Y(n1728) );
  OAI21X1 U1699 ( .A(n155), .B(n1257), .C(n1728), .Y(n1866) );
  NAND2X1 U1700 ( .A(\mem<4><14> ), .B(n156), .Y(n1729) );
  OAI21X1 U1701 ( .A(n155), .B(n1259), .C(n1729), .Y(n1865) );
  NAND2X1 U1702 ( .A(\mem<4><15> ), .B(n156), .Y(n1730) );
  OAI21X1 U1703 ( .A(n155), .B(n1261), .C(n1730), .Y(n1864) );
  NAND2X1 U1704 ( .A(\mem<3><0> ), .B(n159), .Y(n1732) );
  OAI21X1 U1705 ( .A(n158), .B(n1232), .C(n1732), .Y(n1863) );
  NAND2X1 U1706 ( .A(\mem<3><1> ), .B(n159), .Y(n1733) );
  OAI21X1 U1707 ( .A(n158), .B(n1234), .C(n1733), .Y(n1862) );
  NAND2X1 U1708 ( .A(\mem<3><2> ), .B(n159), .Y(n1734) );
  OAI21X1 U1709 ( .A(n158), .B(n1236), .C(n1734), .Y(n1861) );
  NAND2X1 U1710 ( .A(\mem<3><3> ), .B(n159), .Y(n1735) );
  OAI21X1 U1711 ( .A(n158), .B(n1238), .C(n1735), .Y(n1860) );
  NAND2X1 U1712 ( .A(\mem<3><4> ), .B(n159), .Y(n1736) );
  OAI21X1 U1713 ( .A(n158), .B(n1240), .C(n1736), .Y(n1859) );
  NAND2X1 U1714 ( .A(\mem<3><5> ), .B(n159), .Y(n1737) );
  OAI21X1 U1715 ( .A(n158), .B(n1242), .C(n1737), .Y(n1858) );
  NAND2X1 U1716 ( .A(\mem<3><6> ), .B(n159), .Y(n1738) );
  OAI21X1 U1717 ( .A(n158), .B(n1244), .C(n1738), .Y(n1857) );
  NAND2X1 U1718 ( .A(\mem<3><7> ), .B(n159), .Y(n1739) );
  OAI21X1 U1719 ( .A(n158), .B(n1246), .C(n1739), .Y(n1856) );
  NAND2X1 U1720 ( .A(\mem<3><8> ), .B(n159), .Y(n1740) );
  OAI21X1 U1721 ( .A(n158), .B(n1248), .C(n1740), .Y(n1855) );
  NAND2X1 U1722 ( .A(\mem<3><9> ), .B(n159), .Y(n1741) );
  OAI21X1 U1723 ( .A(n158), .B(n1250), .C(n1741), .Y(n1854) );
  NAND2X1 U1724 ( .A(\mem<3><10> ), .B(n159), .Y(n1742) );
  OAI21X1 U1725 ( .A(n158), .B(n1252), .C(n1742), .Y(n1853) );
  NAND2X1 U1726 ( .A(\mem<3><11> ), .B(n159), .Y(n1743) );
  OAI21X1 U1727 ( .A(n158), .B(n1254), .C(n1743), .Y(n1852) );
  NAND2X1 U1728 ( .A(\mem<3><12> ), .B(n159), .Y(n1744) );
  OAI21X1 U1729 ( .A(n158), .B(n1255), .C(n1744), .Y(n1851) );
  NAND2X1 U1730 ( .A(\mem<3><13> ), .B(n159), .Y(n1745) );
  OAI21X1 U1731 ( .A(n158), .B(n1257), .C(n1745), .Y(n1850) );
  NAND2X1 U1732 ( .A(\mem<3><14> ), .B(n159), .Y(n1746) );
  OAI21X1 U1733 ( .A(n158), .B(n1259), .C(n1746), .Y(n1849) );
  NAND2X1 U1734 ( .A(\mem<3><15> ), .B(n159), .Y(n1747) );
  OAI21X1 U1735 ( .A(n158), .B(n1261), .C(n1747), .Y(n1848) );
  NAND2X1 U1736 ( .A(\mem<2><0> ), .B(n162), .Y(n1749) );
  OAI21X1 U1737 ( .A(n161), .B(n1233), .C(n1749), .Y(n1847) );
  NAND2X1 U1738 ( .A(\mem<2><1> ), .B(n162), .Y(n1750) );
  OAI21X1 U1739 ( .A(n161), .B(n1234), .C(n1750), .Y(n1846) );
  NAND2X1 U1740 ( .A(\mem<2><2> ), .B(n162), .Y(n1751) );
  OAI21X1 U1741 ( .A(n161), .B(n1236), .C(n1751), .Y(n1845) );
  NAND2X1 U1742 ( .A(\mem<2><3> ), .B(n162), .Y(n1752) );
  OAI21X1 U1743 ( .A(n161), .B(n1238), .C(n1752), .Y(n1844) );
  NAND2X1 U1744 ( .A(\mem<2><4> ), .B(n162), .Y(n1753) );
  OAI21X1 U1745 ( .A(n161), .B(n1240), .C(n1753), .Y(n1843) );
  NAND2X1 U1746 ( .A(\mem<2><5> ), .B(n162), .Y(n1754) );
  OAI21X1 U1747 ( .A(n161), .B(n1242), .C(n1754), .Y(n1842) );
  NAND2X1 U1748 ( .A(\mem<2><6> ), .B(n162), .Y(n1755) );
  OAI21X1 U1749 ( .A(n161), .B(n1244), .C(n1755), .Y(n1841) );
  NAND2X1 U1750 ( .A(\mem<2><7> ), .B(n162), .Y(n1756) );
  OAI21X1 U1751 ( .A(n161), .B(n1246), .C(n1756), .Y(n1840) );
  NAND2X1 U1752 ( .A(\mem<2><8> ), .B(n162), .Y(n1757) );
  OAI21X1 U1753 ( .A(n161), .B(n1248), .C(n1757), .Y(n1839) );
  NAND2X1 U1754 ( .A(\mem<2><9> ), .B(n162), .Y(n1758) );
  OAI21X1 U1755 ( .A(n161), .B(n1250), .C(n1758), .Y(n1838) );
  NAND2X1 U1756 ( .A(\mem<2><10> ), .B(n162), .Y(n1759) );
  OAI21X1 U1757 ( .A(n161), .B(n1252), .C(n1759), .Y(n1837) );
  NAND2X1 U1758 ( .A(\mem<2><11> ), .B(n162), .Y(n1760) );
  OAI21X1 U1759 ( .A(n161), .B(n1254), .C(n1760), .Y(n1836) );
  NAND2X1 U1760 ( .A(\mem<2><12> ), .B(n162), .Y(n1761) );
  OAI21X1 U1761 ( .A(n161), .B(n1255), .C(n1761), .Y(n1835) );
  NAND2X1 U1762 ( .A(\mem<2><13> ), .B(n162), .Y(n1762) );
  OAI21X1 U1763 ( .A(n161), .B(n1257), .C(n1762), .Y(n1834) );
  NAND2X1 U1764 ( .A(\mem<2><14> ), .B(n162), .Y(n1763) );
  OAI21X1 U1765 ( .A(n161), .B(n1259), .C(n1763), .Y(n1833) );
  NAND2X1 U1766 ( .A(\mem<2><15> ), .B(n162), .Y(n1764) );
  OAI21X1 U1767 ( .A(n161), .B(n1261), .C(n1764), .Y(n1832) );
  NAND2X1 U1768 ( .A(\mem<1><0> ), .B(n165), .Y(n1766) );
  OAI21X1 U1769 ( .A(n164), .B(n1232), .C(n1766), .Y(n1831) );
  NAND2X1 U1770 ( .A(\mem<1><1> ), .B(n165), .Y(n1767) );
  OAI21X1 U1771 ( .A(n164), .B(n1234), .C(n1767), .Y(n1830) );
  NAND2X1 U1772 ( .A(\mem<1><2> ), .B(n165), .Y(n1768) );
  OAI21X1 U1773 ( .A(n164), .B(n1236), .C(n1768), .Y(n1829) );
  NAND2X1 U1774 ( .A(\mem<1><3> ), .B(n165), .Y(n1769) );
  OAI21X1 U1775 ( .A(n164), .B(n1238), .C(n1769), .Y(n1828) );
  NAND2X1 U1776 ( .A(\mem<1><4> ), .B(n165), .Y(n1770) );
  OAI21X1 U1777 ( .A(n164), .B(n1240), .C(n1770), .Y(n1827) );
  NAND2X1 U1778 ( .A(\mem<1><5> ), .B(n165), .Y(n1771) );
  OAI21X1 U1779 ( .A(n164), .B(n1242), .C(n1771), .Y(n1826) );
  NAND2X1 U1780 ( .A(\mem<1><6> ), .B(n165), .Y(n1772) );
  OAI21X1 U1781 ( .A(n164), .B(n1244), .C(n1772), .Y(n1825) );
  NAND2X1 U1782 ( .A(\mem<1><7> ), .B(n165), .Y(n1773) );
  OAI21X1 U1783 ( .A(n164), .B(n1246), .C(n1773), .Y(n1824) );
  NAND2X1 U1784 ( .A(\mem<1><8> ), .B(n165), .Y(n1774) );
  OAI21X1 U1785 ( .A(n164), .B(n1248), .C(n1774), .Y(n1823) );
  NAND2X1 U1786 ( .A(\mem<1><9> ), .B(n165), .Y(n1775) );
  OAI21X1 U1787 ( .A(n164), .B(n1250), .C(n1775), .Y(n1822) );
  NAND2X1 U1788 ( .A(\mem<1><10> ), .B(n165), .Y(n1776) );
  OAI21X1 U1789 ( .A(n164), .B(n1252), .C(n1776), .Y(n1821) );
  NAND2X1 U1790 ( .A(\mem<1><11> ), .B(n165), .Y(n1777) );
  OAI21X1 U1791 ( .A(n164), .B(n1254), .C(n1777), .Y(n1820) );
  NAND2X1 U1792 ( .A(\mem<1><12> ), .B(n165), .Y(n1778) );
  OAI21X1 U1793 ( .A(n164), .B(n1255), .C(n1778), .Y(n1819) );
  NAND2X1 U1794 ( .A(\mem<1><13> ), .B(n165), .Y(n1779) );
  OAI21X1 U1795 ( .A(n164), .B(n1257), .C(n1779), .Y(n1818) );
  NAND2X1 U1796 ( .A(\mem<1><14> ), .B(n165), .Y(n1780) );
  OAI21X1 U1797 ( .A(n164), .B(n1259), .C(n1780), .Y(n1817) );
  NAND2X1 U1798 ( .A(\mem<1><15> ), .B(n165), .Y(n1781) );
  OAI21X1 U1799 ( .A(n164), .B(n1261), .C(n1781), .Y(n1816) );
  NAND2X1 U1800 ( .A(\mem<0><0> ), .B(n1226), .Y(n1784) );
  OAI21X1 U1801 ( .A(n1225), .B(n1233), .C(n1784), .Y(n1815) );
  NAND2X1 U1802 ( .A(\mem<0><1> ), .B(n3), .Y(n1785) );
  OAI21X1 U1803 ( .A(n1225), .B(n1234), .C(n1785), .Y(n1814) );
  NAND2X1 U1804 ( .A(\mem<0><2> ), .B(n3), .Y(n1786) );
  OAI21X1 U1805 ( .A(n1225), .B(n1236), .C(n1786), .Y(n1813) );
  NAND2X1 U1806 ( .A(\mem<0><3> ), .B(n1227), .Y(n1787) );
  OAI21X1 U1807 ( .A(n1225), .B(n1238), .C(n1787), .Y(n1812) );
  NAND2X1 U1808 ( .A(\mem<0><4> ), .B(n1227), .Y(n1788) );
  OAI21X1 U1809 ( .A(n1225), .B(n1240), .C(n1788), .Y(n1811) );
  NAND2X1 U1810 ( .A(\mem<0><5> ), .B(n1226), .Y(n1789) );
  OAI21X1 U1811 ( .A(n1225), .B(n1242), .C(n1789), .Y(n1810) );
  NAND2X1 U1812 ( .A(\mem<0><6> ), .B(n1226), .Y(n1790) );
  OAI21X1 U1813 ( .A(n1225), .B(n1244), .C(n1790), .Y(n1809) );
  NAND2X1 U1814 ( .A(\mem<0><7> ), .B(n3), .Y(n1791) );
  OAI21X1 U1815 ( .A(n1225), .B(n1246), .C(n1791), .Y(n1808) );
  NAND2X1 U1816 ( .A(\mem<0><8> ), .B(n1227), .Y(n1792) );
  OAI21X1 U1817 ( .A(n1225), .B(n1248), .C(n1792), .Y(n1807) );
  NAND2X1 U1818 ( .A(\mem<0><9> ), .B(n1226), .Y(n1793) );
  OAI21X1 U1819 ( .A(n1225), .B(n1250), .C(n1793), .Y(n1806) );
  NAND2X1 U1820 ( .A(\mem<0><10> ), .B(n1226), .Y(n1794) );
  OAI21X1 U1821 ( .A(n1225), .B(n1252), .C(n1794), .Y(n1805) );
  NAND2X1 U1822 ( .A(\mem<0><11> ), .B(n3), .Y(n1795) );
  OAI21X1 U1823 ( .A(n1225), .B(n1254), .C(n1795), .Y(n1804) );
  NAND2X1 U1824 ( .A(\mem<0><12> ), .B(n3), .Y(n1796) );
  OAI21X1 U1825 ( .A(n1225), .B(n1255), .C(n1796), .Y(n1803) );
  NAND2X1 U1826 ( .A(\mem<0><13> ), .B(n1227), .Y(n1797) );
  OAI21X1 U1827 ( .A(n1225), .B(n1257), .C(n1797), .Y(n1802) );
  NAND2X1 U1828 ( .A(\mem<0><14> ), .B(n1227), .Y(n1798) );
  OAI21X1 U1829 ( .A(n1225), .B(n1259), .C(n1798), .Y(n1801) );
  NAND2X1 U1830 ( .A(\mem<0><15> ), .B(n1226), .Y(n1799) );
  OAI21X1 U1831 ( .A(n1225), .B(n1261), .C(n1799), .Y(n1800) );
endmodule


module memc_Size5_1 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , n56, n57, n65, n73, n81, n89, n97, n105,
         n113, n114, n115, n172, n229, n286, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, net57308, net58992, net59300, net59298, net59428, net59426,
         net59578, net59576, net59846, net59844, net59842, net59840, net59838,
         net59836, net60300, net60296, net60292, net60288, net60286, net60284,
         net60282, net66027, net72395, net72480, net72479, net100826,
         net101283, net101551, net101667, net101707, net101711, net101734,
         net101796, net57403, net57401, net101794, net60298, net60290,
         net57431, net57426, net101672, net101670, net101709, net60860,
         net60858, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n31, n33, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n58, n59, n60, n61, n62,
         n63, n64, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n106, n107, n108,
         n109, n110, n111, n112, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n287, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;
  assign \data_out<1>  = net100826;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n447), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n446), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n445), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n444), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n443), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n442), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n441), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n440), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n439), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n438), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n437), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n436), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n435), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n434), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n433), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n432), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n431), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n430), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n429), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n428), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n427), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n426), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n425), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n424), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n423), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n422), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n421), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n420), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n419), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n418), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n417), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n416), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n415), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n414), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n413), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n412), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n411), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n410), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n409), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n408), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n407), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n406), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n405), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n404), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n403), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n402), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n401), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n400), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n399), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n398), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n397), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n396), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n395), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n394), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n393), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n392), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n391), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n390), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n389), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n388), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n387), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n386), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n385), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n384), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n383), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n382), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n381), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n380), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n379), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n378), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n377), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n376), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n375), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n374), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n373), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n372), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n371), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n370), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n369), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n368), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n367), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n366), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n365), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n364), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n363), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n362), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n361), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n360), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n359), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n358), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n357), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n356), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n355), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n354), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n353), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n352), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n351), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n350), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n349), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n348), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n347), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n346), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n345), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n344), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n343), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n342), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n341), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n340), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n339), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n338), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n337), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n336), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n335), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n334), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n333), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n332), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n331), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n330), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n329), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n328), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n327), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n326), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n325), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n324), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n323), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n322), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n321), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n320), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n319), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n318), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n317), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n316), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n315), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n314), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n313), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n312), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n311), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n310), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n309), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n308), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n307), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n306), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n305), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n304), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n303), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n302), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n301), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n300), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n299), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n298), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n297), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n296), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n292), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n291), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n290), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n289), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n288), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(write), .B(net58992), .Y(n56) );
  OAI21X1 U50 ( .A(n610), .B(n677), .C(n531), .Y(n288) );
  OAI21X1 U52 ( .A(n610), .B(n676), .C(n529), .Y(n289) );
  OAI21X1 U54 ( .A(n610), .B(n675), .C(n527), .Y(n290) );
  OAI21X1 U56 ( .A(n610), .B(n674), .C(n525), .Y(n291) );
  OAI21X1 U58 ( .A(n610), .B(n673), .C(n523), .Y(n292) );
  OAI21X1 U62 ( .A(n677), .B(n672), .C(n521), .Y(n293) );
  OAI21X1 U64 ( .A(n676), .B(n672), .C(n519), .Y(n294) );
  OAI21X1 U66 ( .A(n675), .B(n672), .C(n517), .Y(n295) );
  OAI21X1 U68 ( .A(n674), .B(n672), .C(n515), .Y(n296) );
  OAI21X1 U70 ( .A(n673), .B(n672), .C(n513), .Y(n297) );
  OAI21X1 U74 ( .A(n677), .B(n670), .C(n511), .Y(n298) );
  OAI21X1 U76 ( .A(n676), .B(n670), .C(n509), .Y(n299) );
  OAI21X1 U78 ( .A(n675), .B(n670), .C(n507), .Y(n300) );
  OAI21X1 U80 ( .A(n674), .B(n670), .C(n505), .Y(n301) );
  OAI21X1 U82 ( .A(n673), .B(n670), .C(n503), .Y(n302) );
  OAI21X1 U86 ( .A(n677), .B(n668), .C(n501), .Y(n303) );
  OAI21X1 U88 ( .A(n676), .B(n668), .C(n499), .Y(n304) );
  OAI21X1 U90 ( .A(n675), .B(n668), .C(n497), .Y(n305) );
  OAI21X1 U92 ( .A(n674), .B(n668), .C(n495), .Y(n306) );
  OAI21X1 U94 ( .A(n673), .B(n668), .C(n493), .Y(n307) );
  OAI21X1 U98 ( .A(n677), .B(n666), .C(n491), .Y(n308) );
  OAI21X1 U100 ( .A(n676), .B(n666), .C(n489), .Y(n309) );
  OAI21X1 U102 ( .A(n675), .B(n666), .C(n487), .Y(n310) );
  OAI21X1 U104 ( .A(n674), .B(n666), .C(n485), .Y(n311) );
  OAI21X1 U106 ( .A(n673), .B(n666), .C(n483), .Y(n312) );
  OAI21X1 U110 ( .A(n677), .B(n664), .C(n481), .Y(n313) );
  OAI21X1 U112 ( .A(n676), .B(n664), .C(n479), .Y(n314) );
  OAI21X1 U114 ( .A(n675), .B(n664), .C(n477), .Y(n315) );
  OAI21X1 U116 ( .A(n674), .B(n664), .C(n475), .Y(n316) );
  OAI21X1 U118 ( .A(n673), .B(n664), .C(n473), .Y(n317) );
  OAI21X1 U122 ( .A(n677), .B(n662), .C(n471), .Y(n318) );
  OAI21X1 U124 ( .A(n676), .B(n662), .C(n469), .Y(n319) );
  OAI21X1 U126 ( .A(n675), .B(n662), .C(n467), .Y(n320) );
  OAI21X1 U128 ( .A(n674), .B(n662), .C(n465), .Y(n321) );
  OAI21X1 U130 ( .A(n673), .B(n662), .C(n463), .Y(n322) );
  OAI21X1 U134 ( .A(n677), .B(n660), .C(n461), .Y(n323) );
  OAI21X1 U136 ( .A(n676), .B(n660), .C(n459), .Y(n324) );
  OAI21X1 U138 ( .A(n675), .B(n660), .C(n457), .Y(n325) );
  OAI21X1 U140 ( .A(n674), .B(n660), .C(n455), .Y(n326) );
  OAI21X1 U142 ( .A(n673), .B(n660), .C(n453), .Y(n327) );
  NAND3X1 U146 ( .A(net59426), .B(n115), .C(net59298), .Y(n114) );
  OAI21X1 U147 ( .A(n677), .B(n658), .C(n451), .Y(n328) );
  OAI21X1 U149 ( .A(n676), .B(n658), .C(n449), .Y(n329) );
  OAI21X1 U151 ( .A(n675), .B(n658), .C(n287), .Y(n330) );
  OAI21X1 U153 ( .A(n674), .B(n658), .C(n284), .Y(n331) );
  OAI21X1 U155 ( .A(n673), .B(n658), .C(n282), .Y(n332) );
  OAI21X1 U159 ( .A(n677), .B(n656), .C(n280), .Y(n333) );
  OAI21X1 U161 ( .A(n676), .B(n656), .C(n278), .Y(n334) );
  OAI21X1 U163 ( .A(n675), .B(n656), .C(n276), .Y(n335) );
  OAI21X1 U165 ( .A(n674), .B(n656), .C(n274), .Y(n336) );
  OAI21X1 U167 ( .A(n673), .B(n656), .C(n272), .Y(n337) );
  OAI21X1 U171 ( .A(n677), .B(n654), .C(n270), .Y(n338) );
  OAI21X1 U173 ( .A(n676), .B(n654), .C(n268), .Y(n339) );
  OAI21X1 U175 ( .A(n675), .B(n654), .C(n266), .Y(n340) );
  OAI21X1 U177 ( .A(n674), .B(n654), .C(n264), .Y(n341) );
  OAI21X1 U179 ( .A(n673), .B(n654), .C(n262), .Y(n342) );
  OAI21X1 U183 ( .A(n677), .B(n652), .C(n260), .Y(n343) );
  OAI21X1 U185 ( .A(n676), .B(n652), .C(n258), .Y(n344) );
  OAI21X1 U187 ( .A(n675), .B(n652), .C(n256), .Y(n345) );
  OAI21X1 U189 ( .A(n674), .B(n652), .C(n254), .Y(n346) );
  OAI21X1 U191 ( .A(n673), .B(n652), .C(n252), .Y(n347) );
  OAI21X1 U195 ( .A(n677), .B(n650), .C(n250), .Y(n348) );
  OAI21X1 U197 ( .A(n676), .B(n650), .C(n248), .Y(n349) );
  OAI21X1 U199 ( .A(n675), .B(n650), .C(n246), .Y(n350) );
  OAI21X1 U201 ( .A(n674), .B(n650), .C(n244), .Y(n351) );
  OAI21X1 U203 ( .A(n673), .B(n650), .C(n242), .Y(n352) );
  OAI21X1 U207 ( .A(n677), .B(n648), .C(n240), .Y(n353) );
  OAI21X1 U209 ( .A(n676), .B(n648), .C(n238), .Y(n354) );
  OAI21X1 U211 ( .A(n675), .B(n648), .C(n236), .Y(n355) );
  OAI21X1 U213 ( .A(n674), .B(n648), .C(n234), .Y(n356) );
  OAI21X1 U215 ( .A(n673), .B(n648), .C(n232), .Y(n357) );
  OAI21X1 U219 ( .A(n677), .B(n645), .C(n230), .Y(n358) );
  OAI21X1 U221 ( .A(n676), .B(n645), .C(n227), .Y(n359) );
  OAI21X1 U223 ( .A(n675), .B(n645), .C(n225), .Y(n360) );
  OAI21X1 U225 ( .A(n674), .B(n645), .C(n223), .Y(n361) );
  OAI21X1 U227 ( .A(n673), .B(n645), .C(n221), .Y(n362) );
  OAI21X1 U231 ( .A(n677), .B(n643), .C(n219), .Y(n363) );
  OAI21X1 U233 ( .A(n676), .B(n643), .C(n217), .Y(n364) );
  OAI21X1 U235 ( .A(n675), .B(n643), .C(n215), .Y(n365) );
  OAI21X1 U237 ( .A(n674), .B(n643), .C(n213), .Y(n366) );
  OAI21X1 U239 ( .A(n673), .B(n643), .C(n211), .Y(n367) );
  NAND3X1 U243 ( .A(n115), .B(net59428), .C(net59298), .Y(n172) );
  OAI21X1 U244 ( .A(n677), .B(n642), .C(n209), .Y(n368) );
  OAI21X1 U246 ( .A(n676), .B(n642), .C(n207), .Y(n369) );
  OAI21X1 U248 ( .A(n675), .B(n642), .C(n205), .Y(n370) );
  OAI21X1 U250 ( .A(n674), .B(n642), .C(n203), .Y(n371) );
  OAI21X1 U252 ( .A(n673), .B(n642), .C(n201), .Y(n372) );
  OAI21X1 U256 ( .A(n677), .B(n640), .C(n199), .Y(n373) );
  OAI21X1 U258 ( .A(n676), .B(n640), .C(n197), .Y(n374) );
  OAI21X1 U260 ( .A(n675), .B(n640), .C(n195), .Y(n375) );
  OAI21X1 U262 ( .A(n674), .B(n640), .C(n193), .Y(n376) );
  OAI21X1 U264 ( .A(n673), .B(n640), .C(n191), .Y(n377) );
  OAI21X1 U268 ( .A(n677), .B(n638), .C(n189), .Y(n378) );
  OAI21X1 U270 ( .A(n676), .B(n638), .C(n187), .Y(n379) );
  OAI21X1 U272 ( .A(n675), .B(n638), .C(n185), .Y(n380) );
  OAI21X1 U274 ( .A(n674), .B(n638), .C(n183), .Y(n381) );
  OAI21X1 U276 ( .A(n673), .B(n638), .C(n181), .Y(n382) );
  OAI21X1 U280 ( .A(n677), .B(n636), .C(n179), .Y(n383) );
  OAI21X1 U282 ( .A(n676), .B(n636), .C(n177), .Y(n384) );
  OAI21X1 U284 ( .A(n675), .B(n636), .C(n175), .Y(n385) );
  OAI21X1 U286 ( .A(n674), .B(n636), .C(n173), .Y(n386) );
  OAI21X1 U288 ( .A(n673), .B(n636), .C(n170), .Y(n387) );
  OAI21X1 U292 ( .A(n677), .B(n634), .C(n168), .Y(n388) );
  OAI21X1 U294 ( .A(n676), .B(n634), .C(n166), .Y(n389) );
  OAI21X1 U296 ( .A(n675), .B(n634), .C(n164), .Y(n390) );
  OAI21X1 U298 ( .A(n674), .B(n634), .C(n162), .Y(n391) );
  OAI21X1 U300 ( .A(n673), .B(n634), .C(n160), .Y(n392) );
  OAI21X1 U304 ( .A(n677), .B(n632), .C(n158), .Y(n393) );
  OAI21X1 U306 ( .A(n676), .B(n632), .C(n156), .Y(n394) );
  OAI21X1 U308 ( .A(n675), .B(n632), .C(n154), .Y(n395) );
  OAI21X1 U310 ( .A(n674), .B(n632), .C(n152), .Y(n396) );
  OAI21X1 U312 ( .A(n673), .B(n632), .C(n150), .Y(n397) );
  OAI21X1 U316 ( .A(n677), .B(n629), .C(n148), .Y(n398) );
  OAI21X1 U318 ( .A(n676), .B(n629), .C(n146), .Y(n399) );
  OAI21X1 U320 ( .A(n675), .B(n629), .C(n144), .Y(n400) );
  OAI21X1 U322 ( .A(n674), .B(n629), .C(n142), .Y(n401) );
  OAI21X1 U324 ( .A(n673), .B(n629), .C(n140), .Y(n402) );
  OAI21X1 U328 ( .A(n677), .B(n627), .C(n138), .Y(n403) );
  OAI21X1 U330 ( .A(n676), .B(n627), .C(n136), .Y(n404) );
  OAI21X1 U332 ( .A(n675), .B(n627), .C(n134), .Y(n405) );
  OAI21X1 U334 ( .A(n674), .B(n627), .C(n132), .Y(n406) );
  OAI21X1 U336 ( .A(n673), .B(n627), .C(n130), .Y(n407) );
  NAND3X1 U340 ( .A(n115), .B(net59300), .C(net59426), .Y(n229) );
  OAI21X1 U341 ( .A(n677), .B(n626), .C(n128), .Y(n408) );
  OAI21X1 U343 ( .A(n676), .B(n626), .C(n126), .Y(n409) );
  OAI21X1 U345 ( .A(n675), .B(n626), .C(n124), .Y(n410) );
  OAI21X1 U347 ( .A(n674), .B(n626), .C(n122), .Y(n411) );
  OAI21X1 U349 ( .A(n673), .B(n626), .C(n120), .Y(n412) );
  NOR3X1 U353 ( .A(net59844), .B(net66027), .C(net59578), .Y(n57) );
  OAI21X1 U354 ( .A(n677), .B(n624), .C(n118), .Y(n413) );
  OAI21X1 U356 ( .A(n676), .B(n624), .C(n116), .Y(n414) );
  OAI21X1 U358 ( .A(n675), .B(n624), .C(n111), .Y(n415) );
  OAI21X1 U360 ( .A(n674), .B(n624), .C(n109), .Y(n416) );
  OAI21X1 U362 ( .A(n673), .B(n624), .C(n107), .Y(n417) );
  NOR3X1 U366 ( .A(net59846), .B(net101551), .C(net59578), .Y(n65) );
  OAI21X1 U367 ( .A(n677), .B(n622), .C(n104), .Y(n418) );
  OAI21X1 U369 ( .A(n676), .B(n622), .C(n102), .Y(n419) );
  OAI21X1 U371 ( .A(n675), .B(n622), .C(n100), .Y(n420) );
  OAI21X1 U373 ( .A(n674), .B(n622), .C(n98), .Y(n421) );
  OAI21X1 U375 ( .A(n673), .B(n622), .C(n95), .Y(n422) );
  NOR3X1 U379 ( .A(net60296), .B(net59842), .C(net59578), .Y(n73) );
  OAI21X1 U380 ( .A(n677), .B(n620), .C(n93), .Y(n423) );
  OAI21X1 U382 ( .A(n676), .B(n620), .C(n91), .Y(n424) );
  OAI21X1 U384 ( .A(n675), .B(n620), .C(n88), .Y(n425) );
  OAI21X1 U386 ( .A(n674), .B(n620), .C(n86), .Y(n426) );
  OAI21X1 U388 ( .A(n673), .B(n620), .C(n84), .Y(n427) );
  NOR3X1 U392 ( .A(net101667), .B(net59838), .C(net101707), .Y(n81) );
  OAI21X1 U393 ( .A(n677), .B(n618), .C(n82), .Y(n428) );
  OAI21X1 U395 ( .A(n676), .B(n618), .C(n79), .Y(n429) );
  OAI21X1 U397 ( .A(n675), .B(n618), .C(n77), .Y(n430) );
  OAI21X1 U399 ( .A(n674), .B(n618), .C(n75), .Y(n431) );
  OAI21X1 U401 ( .A(n673), .B(n618), .C(n72), .Y(n432) );
  NOR3X1 U405 ( .A(net66027), .B(net59576), .C(net59846), .Y(n89) );
  OAI21X1 U406 ( .A(n677), .B(n616), .C(n70), .Y(n433) );
  OAI21X1 U408 ( .A(n676), .B(n616), .C(n68), .Y(n434) );
  OAI21X1 U410 ( .A(n675), .B(n616), .C(n66), .Y(n435) );
  OAI21X1 U412 ( .A(n674), .B(n616), .C(n63), .Y(n436) );
  OAI21X1 U414 ( .A(n673), .B(n616), .C(n61), .Y(n437) );
  NOR3X1 U418 ( .A(net101551), .B(net59576), .C(net59846), .Y(n97) );
  OAI21X1 U419 ( .A(n677), .B(n613), .C(n59), .Y(n438) );
  OAI21X1 U421 ( .A(n676), .B(n613), .C(n55), .Y(n439) );
  OAI21X1 U423 ( .A(n675), .B(n613), .C(n53), .Y(n440) );
  OAI21X1 U425 ( .A(n674), .B(n613), .C(n51), .Y(n441) );
  OAI21X1 U427 ( .A(n673), .B(n613), .C(n49), .Y(n442) );
  NOR3X1 U431 ( .A(net59838), .B(net59576), .C(net66027), .Y(n105) );
  OAI21X1 U432 ( .A(n677), .B(n611), .C(n47), .Y(n443) );
  OAI21X1 U435 ( .A(n676), .B(n611), .C(n45), .Y(n444) );
  OAI21X1 U438 ( .A(n675), .B(n611), .C(n43), .Y(n445) );
  OAI21X1 U441 ( .A(n674), .B(n611), .C(n41), .Y(n446) );
  OAI21X1 U444 ( .A(n673), .B(n611), .C(n39), .Y(n447) );
  NOR3X1 U448 ( .A(net59838), .B(net59576), .C(net101667), .Y(n113) );
  NAND3X1 U449 ( .A(net59428), .B(net59300), .C(n115), .Y(n286) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n115) );
  OR2X2 U3 ( .A(n708), .B(net57308), .Y(n29) );
  INVX2 U4 ( .A(n29), .Y(\data_out<0> ) );
  OR2X2 U5 ( .A(n739), .B(net57308), .Y(n31) );
  INVX2 U6 ( .A(n31), .Y(\data_out<2> ) );
  INVX4 U7 ( .A(net60298), .Y(net60290) );
  INVX1 U8 ( .A(N12), .Y(net101734) );
  AND2X1 U9 ( .A(n794), .B(net72395), .Y(n532) );
  INVX1 U10 ( .A(N12), .Y(net101283) );
  AND2X1 U11 ( .A(\mem<29><4> ), .B(n604), .Y(n502) );
  AND2X1 U12 ( .A(\mem<27><4> ), .B(n600), .Y(n482) );
  AND2X1 U13 ( .A(\mem<26><4> ), .B(n598), .Y(n472) );
  AND2X1 U14 ( .A(\mem<25><4> ), .B(n596), .Y(n462) );
  AND2X1 U15 ( .A(\mem<24><4> ), .B(n594), .Y(n452) );
  AND2X1 U16 ( .A(\mem<23><4> ), .B(n592), .Y(n281) );
  AND2X1 U17 ( .A(\mem<22><4> ), .B(n590), .Y(n271) );
  AND2X1 U18 ( .A(\mem<21><4> ), .B(n588), .Y(n261) );
  AND2X1 U19 ( .A(\mem<20><4> ), .B(n586), .Y(n251) );
  AND2X1 U20 ( .A(\mem<19><4> ), .B(n584), .Y(n241) );
  AND2X1 U21 ( .A(\mem<18><4> ), .B(n582), .Y(n231) );
  AND2X1 U22 ( .A(\mem<17><4> ), .B(n580), .Y(n220) );
  AND2X1 U23 ( .A(\mem<16><4> ), .B(n578), .Y(n210) );
  AND2X1 U24 ( .A(\mem<15><4> ), .B(n576), .Y(n200) );
  AND2X1 U25 ( .A(\mem<14><4> ), .B(n574), .Y(n190) );
  AND2X1 U26 ( .A(\mem<13><4> ), .B(n572), .Y(n180) );
  AND2X1 U27 ( .A(\mem<12><4> ), .B(n570), .Y(n169) );
  AND2X1 U28 ( .A(\mem<11><4> ), .B(n568), .Y(n159) );
  AND2X1 U29 ( .A(\mem<10><4> ), .B(n566), .Y(n149) );
  AND2X1 U30 ( .A(\mem<9><4> ), .B(n564), .Y(n139) );
  AND2X1 U31 ( .A(\mem<8><4> ), .B(n562), .Y(n129) );
  AND2X1 U32 ( .A(\mem<7><4> ), .B(n560), .Y(n119) );
  AND2X1 U33 ( .A(\mem<6><4> ), .B(n558), .Y(n106) );
  AND2X1 U34 ( .A(\mem<5><4> ), .B(n556), .Y(n94) );
  AND2X1 U35 ( .A(\mem<4><4> ), .B(n554), .Y(n83) );
  AND2X1 U36 ( .A(\mem<3><4> ), .B(n552), .Y(n71) );
  AND2X1 U37 ( .A(\mem<2><4> ), .B(n550), .Y(n60) );
  AND2X1 U38 ( .A(\mem<1><4> ), .B(n548), .Y(n48) );
  AND2X1 U39 ( .A(\mem<0><4> ), .B(n546), .Y(n38) );
  INVX8 U40 ( .A(net60858), .Y(net60298) );
  INVX4 U41 ( .A(net60860), .Y(net60858) );
  INVX1 U42 ( .A(N10), .Y(net60860) );
  INVX8 U43 ( .A(net60858), .Y(net60296) );
  INVX8 U44 ( .A(net60858), .Y(net60300) );
  MUX2X1 U45 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(net101709), .Y(n1) );
  INVX1 U46 ( .A(net60298), .Y(net101709) );
  MUX2X1 U47 ( .B(net57431), .A(n1), .S(net59844), .Y(net57426) );
  MUX2X1 U48 ( .B(n4), .A(n3), .S(net59428), .Y(n2) );
  MUX2X1 U49 ( .B(n5), .A(n6), .S(N12), .Y(n4) );
  MUX2X1 U51 ( .B(n9), .A(n10), .S(net59836), .Y(n5) );
  MUX2X1 U53 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(net60290), .Y(n9) );
  MUX2X1 U55 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(net101672), .Y(n10) );
  INVX1 U57 ( .A(net60298), .Y(net101672) );
  INVX4 U59 ( .A(net59844), .Y(net59836) );
  MUX2X1 U60 ( .B(n7), .A(n8), .S(net59838), .Y(n6) );
  MUX2X1 U61 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(net60288), .Y(n7) );
  INVX8 U63 ( .A(net60298), .Y(net60288) );
  MUX2X1 U65 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(net101796), .Y(n8) );
  INVX1 U67 ( .A(net60298), .Y(net101796) );
  INVX8 U69 ( .A(net59844), .Y(net59838) );
  MUX2X1 U71 ( .B(net57426), .A(n11), .S(N12), .Y(n3) );
  MUX2X1 U72 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(net101670), .Y(net57431)
         );
  INVX1 U73 ( .A(net60300), .Y(net101670) );
  INVX8 U75 ( .A(N11), .Y(net59844) );
  MUX2X1 U77 ( .B(n12), .A(n13), .S(net59842), .Y(n11) );
  MUX2X1 U79 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(net60288), .Y(n12) );
  MUX2X1 U81 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(net60290), .Y(n13) );
  INVX2 U83 ( .A(net59844), .Y(net59842) );
  INVX8 U84 ( .A(N13), .Y(net59428) );
  MUX2X1 U85 ( .B(n2), .A(net57403), .S(net59298), .Y(net57401) );
  INVX1 U87 ( .A(n14), .Y(net100826) );
  OR2X1 U89 ( .A(net57401), .B(net57308), .Y(n14) );
  MUX2X1 U91 ( .B(n15), .A(n16), .S(N13), .Y(net57403) );
  MUX2X1 U93 ( .B(n23), .A(n24), .S(N12), .Y(n15) );
  MUX2X1 U95 ( .B(n27), .A(n28), .S(net59838), .Y(n23) );
  MUX2X1 U96 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(net60288), .Y(n27) );
  MUX2X1 U97 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(net60288), .Y(n28) );
  MUX2X1 U99 ( .B(n25), .A(n26), .S(net59838), .Y(n24) );
  MUX2X1 U101 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(net60286), .Y(n25) );
  INVX8 U103 ( .A(net60296), .Y(net60286) );
  MUX2X1 U105 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(net60288), .Y(n26) );
  MUX2X1 U107 ( .B(n17), .A(n18), .S(N12), .Y(n16) );
  MUX2X1 U108 ( .B(n21), .A(n22), .S(net59838), .Y(n17) );
  MUX2X1 U109 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(net60288), .Y(n21) );
  MUX2X1 U111 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(net101794), .Y(n22) );
  INVX1 U113 ( .A(net60296), .Y(net101794) );
  MUX2X1 U115 ( .B(n19), .A(n20), .S(net59842), .Y(n18) );
  MUX2X1 U117 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(net60288), .Y(n19) );
  MUX2X1 U119 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(net60286), .Y(n20) );
  INVX8 U120 ( .A(net59300), .Y(net59298) );
  OR2X2 U121 ( .A(write), .B(rst), .Y(net57308) );
  INVX1 U123 ( .A(N12), .Y(net101707) );
  INVX1 U125 ( .A(rst), .Y(net58992) );
  OR2X1 U127 ( .A(n770), .B(net57308), .Y(n33) );
  MUX2X1 U129 ( .B(n697), .A(n696), .S(N12), .Y(n705) );
  MUX2X1 U131 ( .B(n713), .A(n714), .S(net101734), .Y(n722) );
  MUX2X1 U132 ( .B(n799), .A(n798), .S(N14), .Y(n800) );
  INVX1 U133 ( .A(net60300), .Y(net101711) );
  MUX2X1 U135 ( .B(n727), .A(n728), .S(net101707), .Y(n736) );
  INVX2 U137 ( .A(net60300), .Y(net101551) );
  INVX1 U139 ( .A(n33), .Y(\data_out<3> ) );
  INVX4 U141 ( .A(net60300), .Y(net101667) );
  INVX4 U143 ( .A(net59578), .Y(net59576) );
  MUX2X1 U144 ( .B(n768), .A(n769), .S(net59300), .Y(n770) );
  MUX2X1 U145 ( .B(\mem<1><2> ), .A(\mem<0><2> ), .S(net72480), .Y(n710) );
  MUX2X1 U148 ( .B(n719), .A(n720), .S(net101283), .Y(n721) );
  INVX8 U150 ( .A(net59428), .Y(net59426) );
  OR2X2 U152 ( .A(net57308), .B(n800), .Y(n35) );
  INVX1 U154 ( .A(n35), .Y(\data_out<4> ) );
  AND2X2 U156 ( .A(n533), .B(n540), .Y(n37) );
  INVX1 U157 ( .A(n38), .Y(n39) );
  AND2X2 U158 ( .A(\mem<0><3> ), .B(n546), .Y(n40) );
  INVX1 U160 ( .A(n40), .Y(n41) );
  AND2X2 U162 ( .A(\mem<0><2> ), .B(n546), .Y(n42) );
  INVX1 U164 ( .A(n42), .Y(n43) );
  AND2X2 U166 ( .A(\mem<0><1> ), .B(n546), .Y(n44) );
  INVX1 U168 ( .A(n44), .Y(n45) );
  AND2X2 U169 ( .A(\mem<0><0> ), .B(n546), .Y(n46) );
  INVX1 U170 ( .A(n46), .Y(n47) );
  INVX1 U172 ( .A(n48), .Y(n49) );
  AND2X2 U174 ( .A(\mem<1><3> ), .B(n548), .Y(n50) );
  INVX1 U176 ( .A(n50), .Y(n51) );
  AND2X2 U178 ( .A(\mem<1><2> ), .B(n548), .Y(n52) );
  INVX1 U180 ( .A(n52), .Y(n53) );
  AND2X2 U181 ( .A(\mem<1><1> ), .B(n548), .Y(n54) );
  INVX1 U182 ( .A(n54), .Y(n55) );
  AND2X2 U184 ( .A(\mem<1><0> ), .B(n548), .Y(n58) );
  INVX1 U186 ( .A(n58), .Y(n59) );
  INVX1 U188 ( .A(n60), .Y(n61) );
  AND2X2 U190 ( .A(\mem<2><3> ), .B(n550), .Y(n62) );
  INVX1 U192 ( .A(n62), .Y(n63) );
  AND2X2 U193 ( .A(\mem<2><2> ), .B(n550), .Y(n64) );
  INVX1 U194 ( .A(n64), .Y(n66) );
  AND2X2 U196 ( .A(\mem<2><1> ), .B(n550), .Y(n67) );
  INVX1 U198 ( .A(n67), .Y(n68) );
  AND2X2 U200 ( .A(\mem<2><0> ), .B(n550), .Y(n69) );
  INVX1 U202 ( .A(n69), .Y(n70) );
  INVX1 U204 ( .A(n71), .Y(n72) );
  AND2X2 U205 ( .A(\mem<3><3> ), .B(n552), .Y(n74) );
  INVX1 U206 ( .A(n74), .Y(n75) );
  AND2X2 U208 ( .A(\mem<3><2> ), .B(n552), .Y(n76) );
  INVX1 U210 ( .A(n76), .Y(n77) );
  AND2X2 U212 ( .A(\mem<3><1> ), .B(n552), .Y(n78) );
  INVX1 U214 ( .A(n78), .Y(n79) );
  AND2X2 U216 ( .A(\mem<3><0> ), .B(n552), .Y(n80) );
  INVX1 U217 ( .A(n80), .Y(n82) );
  INVX1 U218 ( .A(n83), .Y(n84) );
  AND2X2 U220 ( .A(\mem<4><3> ), .B(n554), .Y(n85) );
  INVX1 U222 ( .A(n85), .Y(n86) );
  AND2X2 U224 ( .A(\mem<4><2> ), .B(n554), .Y(n87) );
  INVX1 U226 ( .A(n87), .Y(n88) );
  AND2X2 U228 ( .A(\mem<4><1> ), .B(n554), .Y(n90) );
  INVX1 U229 ( .A(n90), .Y(n91) );
  AND2X2 U230 ( .A(\mem<4><0> ), .B(n554), .Y(n92) );
  INVX1 U232 ( .A(n92), .Y(n93) );
  INVX1 U234 ( .A(n94), .Y(n95) );
  AND2X2 U236 ( .A(\mem<5><3> ), .B(n556), .Y(n96) );
  INVX1 U238 ( .A(n96), .Y(n98) );
  AND2X2 U240 ( .A(\mem<5><2> ), .B(n556), .Y(n99) );
  INVX1 U241 ( .A(n99), .Y(n100) );
  AND2X2 U242 ( .A(\mem<5><1> ), .B(n556), .Y(n101) );
  INVX1 U245 ( .A(n101), .Y(n102) );
  AND2X2 U247 ( .A(\mem<5><0> ), .B(n556), .Y(n103) );
  INVX1 U249 ( .A(n103), .Y(n104) );
  INVX1 U251 ( .A(n106), .Y(n107) );
  AND2X2 U253 ( .A(\mem<6><3> ), .B(n558), .Y(n108) );
  INVX1 U254 ( .A(n108), .Y(n109) );
  AND2X2 U255 ( .A(\mem<6><2> ), .B(n558), .Y(n110) );
  INVX1 U257 ( .A(n110), .Y(n111) );
  AND2X2 U259 ( .A(\mem<6><1> ), .B(n558), .Y(n112) );
  INVX1 U261 ( .A(n112), .Y(n116) );
  AND2X2 U263 ( .A(\mem<6><0> ), .B(n558), .Y(n117) );
  INVX1 U265 ( .A(n117), .Y(n118) );
  INVX1 U266 ( .A(n119), .Y(n120) );
  AND2X2 U267 ( .A(\mem<7><3> ), .B(n560), .Y(n121) );
  INVX1 U269 ( .A(n121), .Y(n122) );
  AND2X2 U271 ( .A(\mem<7><2> ), .B(n560), .Y(n123) );
  INVX1 U273 ( .A(n123), .Y(n124) );
  AND2X2 U275 ( .A(\mem<7><1> ), .B(n560), .Y(n125) );
  INVX1 U277 ( .A(n125), .Y(n126) );
  AND2X2 U278 ( .A(\mem<7><0> ), .B(n560), .Y(n127) );
  INVX1 U279 ( .A(n127), .Y(n128) );
  INVX1 U281 ( .A(n129), .Y(n130) );
  AND2X2 U283 ( .A(\mem<8><3> ), .B(n562), .Y(n131) );
  INVX1 U285 ( .A(n131), .Y(n132) );
  AND2X2 U287 ( .A(\mem<8><2> ), .B(n562), .Y(n133) );
  INVX1 U289 ( .A(n133), .Y(n134) );
  AND2X2 U290 ( .A(\mem<8><1> ), .B(n562), .Y(n135) );
  INVX1 U291 ( .A(n135), .Y(n136) );
  AND2X2 U293 ( .A(\mem<8><0> ), .B(n562), .Y(n137) );
  INVX1 U295 ( .A(n137), .Y(n138) );
  INVX1 U297 ( .A(n139), .Y(n140) );
  AND2X2 U299 ( .A(\mem<9><3> ), .B(n564), .Y(n141) );
  INVX1 U301 ( .A(n141), .Y(n142) );
  AND2X2 U302 ( .A(\mem<9><2> ), .B(n564), .Y(n143) );
  INVX1 U303 ( .A(n143), .Y(n144) );
  AND2X2 U305 ( .A(\mem<9><1> ), .B(n564), .Y(n145) );
  INVX1 U307 ( .A(n145), .Y(n146) );
  AND2X2 U309 ( .A(\mem<9><0> ), .B(n564), .Y(n147) );
  INVX1 U311 ( .A(n147), .Y(n148) );
  INVX1 U313 ( .A(n149), .Y(n150) );
  AND2X2 U314 ( .A(\mem<10><3> ), .B(n566), .Y(n151) );
  INVX1 U315 ( .A(n151), .Y(n152) );
  AND2X2 U317 ( .A(\mem<10><2> ), .B(n566), .Y(n153) );
  INVX1 U319 ( .A(n153), .Y(n154) );
  AND2X2 U321 ( .A(\mem<10><1> ), .B(n566), .Y(n155) );
  INVX1 U323 ( .A(n155), .Y(n156) );
  AND2X2 U325 ( .A(\mem<10><0> ), .B(n566), .Y(n157) );
  INVX1 U326 ( .A(n157), .Y(n158) );
  INVX1 U327 ( .A(n159), .Y(n160) );
  AND2X2 U329 ( .A(\mem<11><3> ), .B(n568), .Y(n161) );
  INVX1 U331 ( .A(n161), .Y(n162) );
  AND2X2 U333 ( .A(\mem<11><2> ), .B(n568), .Y(n163) );
  INVX1 U335 ( .A(n163), .Y(n164) );
  AND2X2 U337 ( .A(\mem<11><1> ), .B(n568), .Y(n165) );
  INVX1 U338 ( .A(n165), .Y(n166) );
  AND2X2 U339 ( .A(\mem<11><0> ), .B(n568), .Y(n167) );
  INVX1 U342 ( .A(n167), .Y(n168) );
  INVX1 U344 ( .A(n169), .Y(n170) );
  AND2X2 U346 ( .A(\mem<12><3> ), .B(n570), .Y(n171) );
  INVX1 U348 ( .A(n171), .Y(n173) );
  AND2X2 U350 ( .A(\mem<12><2> ), .B(n570), .Y(n174) );
  INVX1 U351 ( .A(n174), .Y(n175) );
  AND2X2 U352 ( .A(\mem<12><1> ), .B(n570), .Y(n176) );
  INVX1 U355 ( .A(n176), .Y(n177) );
  AND2X2 U357 ( .A(\mem<12><0> ), .B(n570), .Y(n178) );
  INVX1 U359 ( .A(n178), .Y(n179) );
  INVX1 U361 ( .A(n180), .Y(n181) );
  AND2X2 U363 ( .A(\mem<13><3> ), .B(n572), .Y(n182) );
  INVX1 U364 ( .A(n182), .Y(n183) );
  AND2X2 U365 ( .A(\mem<13><2> ), .B(n572), .Y(n184) );
  INVX1 U368 ( .A(n184), .Y(n185) );
  AND2X2 U370 ( .A(\mem<13><1> ), .B(n572), .Y(n186) );
  INVX1 U372 ( .A(n186), .Y(n187) );
  AND2X2 U374 ( .A(\mem<13><0> ), .B(n572), .Y(n188) );
  INVX1 U376 ( .A(n188), .Y(n189) );
  INVX1 U377 ( .A(n190), .Y(n191) );
  AND2X2 U378 ( .A(\mem<14><3> ), .B(n574), .Y(n192) );
  INVX1 U381 ( .A(n192), .Y(n193) );
  AND2X2 U383 ( .A(\mem<14><2> ), .B(n574), .Y(n194) );
  INVX1 U385 ( .A(n194), .Y(n195) );
  AND2X2 U387 ( .A(\mem<14><1> ), .B(n574), .Y(n196) );
  INVX1 U389 ( .A(n196), .Y(n197) );
  AND2X2 U390 ( .A(\mem<14><0> ), .B(n574), .Y(n198) );
  INVX1 U391 ( .A(n198), .Y(n199) );
  INVX1 U394 ( .A(n200), .Y(n201) );
  AND2X2 U396 ( .A(\mem<15><3> ), .B(n576), .Y(n202) );
  INVX1 U398 ( .A(n202), .Y(n203) );
  AND2X2 U400 ( .A(\mem<15><2> ), .B(n576), .Y(n204) );
  INVX1 U402 ( .A(n204), .Y(n205) );
  AND2X2 U403 ( .A(\mem<15><1> ), .B(n576), .Y(n206) );
  INVX1 U404 ( .A(n206), .Y(n207) );
  AND2X2 U407 ( .A(\mem<15><0> ), .B(n576), .Y(n208) );
  INVX1 U409 ( .A(n208), .Y(n209) );
  INVX1 U411 ( .A(n210), .Y(n211) );
  AND2X2 U413 ( .A(\mem<16><3> ), .B(n578), .Y(n212) );
  INVX1 U415 ( .A(n212), .Y(n213) );
  AND2X2 U416 ( .A(\mem<16><2> ), .B(n578), .Y(n214) );
  INVX1 U417 ( .A(n214), .Y(n215) );
  AND2X2 U420 ( .A(\mem<16><1> ), .B(n578), .Y(n216) );
  INVX1 U422 ( .A(n216), .Y(n217) );
  AND2X2 U424 ( .A(\mem<16><0> ), .B(n578), .Y(n218) );
  INVX1 U426 ( .A(n218), .Y(n219) );
  INVX1 U428 ( .A(n220), .Y(n221) );
  AND2X2 U429 ( .A(\mem<17><3> ), .B(n580), .Y(n222) );
  INVX1 U430 ( .A(n222), .Y(n223) );
  AND2X2 U433 ( .A(\mem<17><2> ), .B(n580), .Y(n224) );
  INVX1 U434 ( .A(n224), .Y(n225) );
  AND2X2 U436 ( .A(\mem<17><1> ), .B(n580), .Y(n226) );
  INVX1 U437 ( .A(n226), .Y(n227) );
  AND2X2 U439 ( .A(\mem<17><0> ), .B(n580), .Y(n228) );
  INVX1 U440 ( .A(n228), .Y(n230) );
  INVX1 U442 ( .A(n231), .Y(n232) );
  AND2X2 U443 ( .A(\mem<18><3> ), .B(n582), .Y(n233) );
  INVX1 U445 ( .A(n233), .Y(n234) );
  AND2X2 U446 ( .A(\mem<18><2> ), .B(n582), .Y(n235) );
  INVX1 U447 ( .A(n235), .Y(n236) );
  AND2X2 U451 ( .A(\mem<18><1> ), .B(n582), .Y(n237) );
  INVX1 U452 ( .A(n237), .Y(n238) );
  AND2X2 U453 ( .A(\mem<18><0> ), .B(n582), .Y(n239) );
  INVX1 U454 ( .A(n239), .Y(n240) );
  INVX1 U455 ( .A(n241), .Y(n242) );
  AND2X2 U456 ( .A(\mem<19><3> ), .B(n584), .Y(n243) );
  INVX1 U457 ( .A(n243), .Y(n244) );
  AND2X2 U458 ( .A(\mem<19><2> ), .B(n584), .Y(n245) );
  INVX1 U459 ( .A(n245), .Y(n246) );
  AND2X2 U460 ( .A(\mem<19><1> ), .B(n584), .Y(n247) );
  INVX1 U461 ( .A(n247), .Y(n248) );
  AND2X2 U462 ( .A(\mem<19><0> ), .B(n584), .Y(n249) );
  INVX1 U463 ( .A(n249), .Y(n250) );
  INVX1 U464 ( .A(n251), .Y(n252) );
  AND2X2 U465 ( .A(\mem<20><3> ), .B(n586), .Y(n253) );
  INVX1 U466 ( .A(n253), .Y(n254) );
  AND2X2 U467 ( .A(\mem<20><2> ), .B(n586), .Y(n255) );
  INVX1 U468 ( .A(n255), .Y(n256) );
  AND2X2 U469 ( .A(\mem<20><1> ), .B(n586), .Y(n257) );
  INVX1 U470 ( .A(n257), .Y(n258) );
  AND2X2 U471 ( .A(\mem<20><0> ), .B(n586), .Y(n259) );
  INVX1 U472 ( .A(n259), .Y(n260) );
  INVX1 U473 ( .A(n261), .Y(n262) );
  AND2X2 U474 ( .A(\mem<21><3> ), .B(n588), .Y(n263) );
  INVX1 U475 ( .A(n263), .Y(n264) );
  AND2X2 U476 ( .A(\mem<21><2> ), .B(n588), .Y(n265) );
  INVX1 U477 ( .A(n265), .Y(n266) );
  AND2X2 U478 ( .A(\mem<21><1> ), .B(n588), .Y(n267) );
  INVX1 U479 ( .A(n267), .Y(n268) );
  AND2X2 U480 ( .A(\mem<21><0> ), .B(n588), .Y(n269) );
  INVX1 U481 ( .A(n269), .Y(n270) );
  INVX1 U482 ( .A(n271), .Y(n272) );
  AND2X2 U483 ( .A(\mem<22><3> ), .B(n590), .Y(n273) );
  INVX1 U484 ( .A(n273), .Y(n274) );
  AND2X2 U485 ( .A(\mem<22><2> ), .B(n590), .Y(n275) );
  INVX1 U486 ( .A(n275), .Y(n276) );
  AND2X2 U487 ( .A(\mem<22><1> ), .B(n590), .Y(n277) );
  INVX1 U488 ( .A(n277), .Y(n278) );
  AND2X2 U489 ( .A(\mem<22><0> ), .B(n590), .Y(n279) );
  INVX1 U490 ( .A(n279), .Y(n280) );
  INVX1 U491 ( .A(n281), .Y(n282) );
  AND2X2 U492 ( .A(\mem<23><3> ), .B(n592), .Y(n283) );
  INVX1 U493 ( .A(n283), .Y(n284) );
  AND2X2 U494 ( .A(\mem<23><2> ), .B(n592), .Y(n285) );
  INVX1 U495 ( .A(n285), .Y(n287) );
  AND2X2 U496 ( .A(\mem<23><1> ), .B(n592), .Y(n448) );
  INVX1 U497 ( .A(n448), .Y(n449) );
  AND2X2 U498 ( .A(\mem<23><0> ), .B(n592), .Y(n450) );
  INVX1 U499 ( .A(n450), .Y(n451) );
  INVX1 U500 ( .A(n452), .Y(n453) );
  AND2X2 U501 ( .A(\mem<24><3> ), .B(n594), .Y(n454) );
  INVX1 U502 ( .A(n454), .Y(n455) );
  AND2X2 U503 ( .A(\mem<24><2> ), .B(n594), .Y(n456) );
  INVX1 U504 ( .A(n456), .Y(n457) );
  AND2X2 U505 ( .A(\mem<24><1> ), .B(n594), .Y(n458) );
  INVX1 U506 ( .A(n458), .Y(n459) );
  AND2X2 U507 ( .A(\mem<24><0> ), .B(n594), .Y(n460) );
  INVX1 U508 ( .A(n460), .Y(n461) );
  INVX1 U509 ( .A(n462), .Y(n463) );
  AND2X2 U510 ( .A(\mem<25><3> ), .B(n596), .Y(n464) );
  INVX1 U511 ( .A(n464), .Y(n465) );
  AND2X2 U512 ( .A(\mem<25><2> ), .B(n596), .Y(n466) );
  INVX1 U513 ( .A(n466), .Y(n467) );
  AND2X2 U514 ( .A(\mem<25><1> ), .B(n596), .Y(n468) );
  INVX1 U515 ( .A(n468), .Y(n469) );
  AND2X2 U516 ( .A(\mem<25><0> ), .B(n596), .Y(n470) );
  INVX1 U517 ( .A(n470), .Y(n471) );
  INVX1 U518 ( .A(n472), .Y(n473) );
  AND2X2 U519 ( .A(\mem<26><3> ), .B(n598), .Y(n474) );
  INVX1 U520 ( .A(n474), .Y(n475) );
  AND2X2 U521 ( .A(\mem<26><2> ), .B(n598), .Y(n476) );
  INVX1 U522 ( .A(n476), .Y(n477) );
  AND2X2 U523 ( .A(\mem<26><1> ), .B(n598), .Y(n478) );
  INVX1 U524 ( .A(n478), .Y(n479) );
  AND2X2 U525 ( .A(\mem<26><0> ), .B(n598), .Y(n480) );
  INVX1 U526 ( .A(n480), .Y(n481) );
  INVX1 U527 ( .A(n482), .Y(n483) );
  AND2X2 U528 ( .A(\mem<27><3> ), .B(n600), .Y(n484) );
  INVX1 U529 ( .A(n484), .Y(n485) );
  AND2X2 U530 ( .A(\mem<27><2> ), .B(n600), .Y(n486) );
  INVX1 U531 ( .A(n486), .Y(n487) );
  AND2X2 U532 ( .A(\mem<27><1> ), .B(n600), .Y(n488) );
  INVX1 U533 ( .A(n488), .Y(n489) );
  AND2X2 U534 ( .A(\mem<27><0> ), .B(n600), .Y(n490) );
  INVX1 U535 ( .A(n490), .Y(n491) );
  AND2X2 U536 ( .A(\mem<28><4> ), .B(n602), .Y(n492) );
  INVX1 U537 ( .A(n492), .Y(n493) );
  AND2X2 U538 ( .A(\mem<28><3> ), .B(n602), .Y(n494) );
  INVX1 U539 ( .A(n494), .Y(n495) );
  AND2X2 U540 ( .A(\mem<28><2> ), .B(n602), .Y(n496) );
  INVX1 U541 ( .A(n496), .Y(n497) );
  AND2X2 U542 ( .A(\mem<28><1> ), .B(n602), .Y(n498) );
  INVX1 U543 ( .A(n498), .Y(n499) );
  AND2X2 U544 ( .A(\mem<28><0> ), .B(n602), .Y(n500) );
  INVX1 U545 ( .A(n500), .Y(n501) );
  INVX1 U546 ( .A(n502), .Y(n503) );
  AND2X2 U547 ( .A(\mem<29><3> ), .B(n604), .Y(n504) );
  INVX1 U548 ( .A(n504), .Y(n505) );
  AND2X2 U549 ( .A(\mem<29><2> ), .B(n604), .Y(n506) );
  INVX1 U550 ( .A(n506), .Y(n507) );
  AND2X2 U551 ( .A(\mem<29><1> ), .B(n604), .Y(n508) );
  INVX1 U552 ( .A(n508), .Y(n509) );
  AND2X2 U553 ( .A(\mem<29><0> ), .B(n604), .Y(n510) );
  INVX1 U554 ( .A(n510), .Y(n511) );
  AND2X2 U555 ( .A(\mem<30><4> ), .B(n606), .Y(n512) );
  INVX1 U556 ( .A(n512), .Y(n513) );
  AND2X2 U557 ( .A(\mem<30><3> ), .B(n606), .Y(n514) );
  INVX1 U558 ( .A(n514), .Y(n515) );
  AND2X2 U559 ( .A(\mem<30><2> ), .B(n606), .Y(n516) );
  INVX1 U560 ( .A(n516), .Y(n517) );
  AND2X2 U561 ( .A(\mem<30><1> ), .B(n606), .Y(n518) );
  INVX1 U562 ( .A(n518), .Y(n519) );
  AND2X2 U563 ( .A(\mem<30><0> ), .B(n606), .Y(n520) );
  INVX1 U564 ( .A(n520), .Y(n521) );
  AND2X2 U565 ( .A(\mem<31><4> ), .B(n608), .Y(n522) );
  INVX1 U566 ( .A(n522), .Y(n523) );
  AND2X2 U567 ( .A(\mem<31><3> ), .B(n608), .Y(n524) );
  INVX1 U568 ( .A(n524), .Y(n525) );
  AND2X2 U569 ( .A(\mem<31><2> ), .B(n608), .Y(n526) );
  INVX1 U570 ( .A(n526), .Y(n527) );
  AND2X2 U571 ( .A(\mem<31><1> ), .B(n608), .Y(n528) );
  INVX1 U572 ( .A(n528), .Y(n529) );
  AND2X2 U573 ( .A(\mem<31><0> ), .B(n608), .Y(n530) );
  INVX1 U574 ( .A(n530), .Y(n531) );
  INVX1 U575 ( .A(n532), .Y(n533) );
  AND2X1 U576 ( .A(\data_in<4> ), .B(n56), .Y(n534) );
  AND2X1 U577 ( .A(\data_in<3> ), .B(n56), .Y(n535) );
  AND2X1 U578 ( .A(\data_in<2> ), .B(n56), .Y(n536) );
  AND2X1 U579 ( .A(\data_in<1> ), .B(n56), .Y(n537) );
  AND2X1 U580 ( .A(\data_in<0> ), .B(n56), .Y(n538) );
  AND2X2 U581 ( .A(n793), .B(net59838), .Y(n539) );
  INVX1 U582 ( .A(n539), .Y(n540) );
  BUFX2 U583 ( .A(n286), .Y(n541) );
  INVX1 U584 ( .A(n541), .Y(n801) );
  BUFX2 U585 ( .A(n229), .Y(n542) );
  INVX1 U586 ( .A(n542), .Y(n804) );
  BUFX2 U587 ( .A(n172), .Y(n543) );
  INVX1 U588 ( .A(n543), .Y(n802) );
  BUFX2 U589 ( .A(n114), .Y(n544) );
  INVX1 U590 ( .A(n544), .Y(n803) );
  INVX1 U591 ( .A(n534), .Y(n673) );
  INVX1 U592 ( .A(n535), .Y(n674) );
  INVX1 U593 ( .A(n536), .Y(n675) );
  INVX1 U594 ( .A(n537), .Y(n676) );
  INVX1 U595 ( .A(n538), .Y(n677) );
  AND2X1 U596 ( .A(n612), .B(n56), .Y(n545) );
  INVX1 U597 ( .A(n545), .Y(n546) );
  AND2X1 U598 ( .A(n614), .B(n56), .Y(n547) );
  INVX1 U599 ( .A(n547), .Y(n548) );
  AND2X1 U600 ( .A(n615), .B(n56), .Y(n549) );
  INVX1 U601 ( .A(n549), .Y(n550) );
  AND2X1 U602 ( .A(n617), .B(n56), .Y(n551) );
  INVX1 U603 ( .A(n551), .Y(n552) );
  AND2X1 U604 ( .A(n619), .B(n56), .Y(n553) );
  INVX1 U605 ( .A(n553), .Y(n554) );
  AND2X1 U606 ( .A(n621), .B(n56), .Y(n555) );
  INVX1 U607 ( .A(n555), .Y(n556) );
  AND2X1 U608 ( .A(n623), .B(n56), .Y(n557) );
  INVX1 U609 ( .A(n557), .Y(n558) );
  AND2X1 U610 ( .A(n625), .B(n56), .Y(n559) );
  INVX1 U611 ( .A(n559), .Y(n560) );
  AND2X1 U612 ( .A(n628), .B(n56), .Y(n561) );
  INVX1 U613 ( .A(n561), .Y(n562) );
  AND2X1 U614 ( .A(n630), .B(n56), .Y(n563) );
  INVX1 U615 ( .A(n563), .Y(n564) );
  AND2X1 U616 ( .A(n631), .B(n56), .Y(n565) );
  INVX1 U617 ( .A(n565), .Y(n566) );
  AND2X1 U618 ( .A(n633), .B(n56), .Y(n567) );
  INVX1 U619 ( .A(n567), .Y(n568) );
  AND2X1 U620 ( .A(n635), .B(n56), .Y(n569) );
  INVX1 U621 ( .A(n569), .Y(n570) );
  AND2X1 U622 ( .A(n637), .B(n56), .Y(n571) );
  INVX1 U623 ( .A(n571), .Y(n572) );
  AND2X1 U624 ( .A(n639), .B(n56), .Y(n573) );
  INVX1 U625 ( .A(n573), .Y(n574) );
  AND2X1 U626 ( .A(n641), .B(n56), .Y(n575) );
  INVX1 U627 ( .A(n575), .Y(n576) );
  AND2X1 U628 ( .A(n644), .B(n56), .Y(n577) );
  INVX1 U629 ( .A(n577), .Y(n578) );
  AND2X1 U630 ( .A(n646), .B(n56), .Y(n579) );
  INVX1 U631 ( .A(n579), .Y(n580) );
  AND2X1 U632 ( .A(n647), .B(n56), .Y(n581) );
  INVX1 U633 ( .A(n581), .Y(n582) );
  AND2X1 U634 ( .A(n649), .B(n56), .Y(n583) );
  INVX1 U635 ( .A(n583), .Y(n584) );
  AND2X1 U636 ( .A(n651), .B(n56), .Y(n585) );
  INVX1 U637 ( .A(n585), .Y(n586) );
  AND2X1 U638 ( .A(n653), .B(n56), .Y(n587) );
  INVX1 U639 ( .A(n587), .Y(n588) );
  AND2X1 U640 ( .A(n655), .B(n56), .Y(n589) );
  INVX1 U641 ( .A(n589), .Y(n590) );
  AND2X1 U642 ( .A(n657), .B(n56), .Y(n591) );
  INVX1 U643 ( .A(n591), .Y(n592) );
  AND2X1 U644 ( .A(n659), .B(n56), .Y(n593) );
  INVX1 U645 ( .A(n593), .Y(n594) );
  AND2X1 U646 ( .A(n661), .B(n56), .Y(n595) );
  INVX1 U647 ( .A(n595), .Y(n596) );
  AND2X1 U648 ( .A(n663), .B(n56), .Y(n597) );
  INVX1 U649 ( .A(n597), .Y(n598) );
  AND2X1 U650 ( .A(n665), .B(n56), .Y(n599) );
  INVX1 U651 ( .A(n599), .Y(n600) );
  AND2X1 U652 ( .A(n667), .B(n56), .Y(n601) );
  INVX1 U653 ( .A(n601), .Y(n602) );
  AND2X1 U654 ( .A(n669), .B(n56), .Y(n603) );
  INVX1 U655 ( .A(n603), .Y(n604) );
  AND2X1 U656 ( .A(n671), .B(n56), .Y(n605) );
  INVX1 U657 ( .A(n605), .Y(n606) );
  AND2X1 U658 ( .A(n609), .B(n56), .Y(n607) );
  INVX1 U659 ( .A(n607), .Y(n608) );
  AND2X1 U660 ( .A(n57), .B(n803), .Y(n609) );
  INVX1 U661 ( .A(n609), .Y(n610) );
  INVX1 U662 ( .A(n612), .Y(n611) );
  AND2X1 U663 ( .A(n801), .B(n113), .Y(n612) );
  INVX1 U664 ( .A(n614), .Y(n613) );
  AND2X1 U665 ( .A(n801), .B(n105), .Y(n614) );
  AND2X1 U666 ( .A(n801), .B(n97), .Y(n615) );
  INVX1 U667 ( .A(n615), .Y(n616) );
  AND2X1 U668 ( .A(n801), .B(n89), .Y(n617) );
  INVX1 U669 ( .A(n617), .Y(n618) );
  AND2X1 U670 ( .A(n801), .B(n81), .Y(n619) );
  INVX1 U671 ( .A(n619), .Y(n620) );
  AND2X1 U672 ( .A(n801), .B(n73), .Y(n621) );
  INVX1 U673 ( .A(n621), .Y(n622) );
  AND2X1 U674 ( .A(n801), .B(n65), .Y(n623) );
  INVX1 U675 ( .A(n623), .Y(n624) );
  AND2X1 U676 ( .A(n801), .B(n57), .Y(n625) );
  INVX1 U677 ( .A(n625), .Y(n626) );
  INVX1 U678 ( .A(n628), .Y(n627) );
  AND2X1 U679 ( .A(n804), .B(n113), .Y(n628) );
  INVX1 U680 ( .A(n630), .Y(n629) );
  AND2X1 U681 ( .A(n804), .B(n105), .Y(n630) );
  AND2X1 U682 ( .A(n804), .B(n97), .Y(n631) );
  INVX1 U683 ( .A(n631), .Y(n632) );
  AND2X1 U684 ( .A(n804), .B(n89), .Y(n633) );
  INVX1 U685 ( .A(n633), .Y(n634) );
  AND2X1 U686 ( .A(n804), .B(n81), .Y(n635) );
  INVX1 U687 ( .A(n635), .Y(n636) );
  AND2X1 U688 ( .A(n804), .B(n73), .Y(n637) );
  INVX1 U689 ( .A(n637), .Y(n638) );
  AND2X1 U690 ( .A(n804), .B(n65), .Y(n639) );
  INVX1 U691 ( .A(n639), .Y(n640) );
  AND2X1 U692 ( .A(n804), .B(n57), .Y(n641) );
  INVX1 U693 ( .A(n641), .Y(n642) );
  INVX1 U694 ( .A(n644), .Y(n643) );
  AND2X1 U695 ( .A(n802), .B(n113), .Y(n644) );
  INVX1 U696 ( .A(n646), .Y(n645) );
  AND2X1 U697 ( .A(n802), .B(n105), .Y(n646) );
  AND2X1 U698 ( .A(n802), .B(n97), .Y(n647) );
  INVX1 U699 ( .A(n647), .Y(n648) );
  AND2X1 U700 ( .A(n802), .B(n89), .Y(n649) );
  INVX1 U701 ( .A(n649), .Y(n650) );
  AND2X1 U702 ( .A(n802), .B(n81), .Y(n651) );
  INVX1 U703 ( .A(n651), .Y(n652) );
  AND2X1 U704 ( .A(n802), .B(n73), .Y(n653) );
  INVX1 U705 ( .A(n653), .Y(n654) );
  AND2X1 U706 ( .A(n802), .B(n65), .Y(n655) );
  INVX1 U707 ( .A(n655), .Y(n656) );
  AND2X1 U708 ( .A(n802), .B(n57), .Y(n657) );
  INVX1 U709 ( .A(n657), .Y(n658) );
  AND2X1 U710 ( .A(n113), .B(n803), .Y(n659) );
  INVX1 U711 ( .A(n659), .Y(n660) );
  AND2X1 U712 ( .A(n105), .B(n803), .Y(n661) );
  INVX1 U713 ( .A(n661), .Y(n662) );
  AND2X1 U714 ( .A(n97), .B(n803), .Y(n663) );
  INVX1 U715 ( .A(n663), .Y(n664) );
  AND2X1 U716 ( .A(n89), .B(n803), .Y(n665) );
  INVX1 U717 ( .A(n665), .Y(n666) );
  AND2X1 U718 ( .A(n81), .B(n803), .Y(n667) );
  INVX1 U719 ( .A(n667), .Y(n668) );
  AND2X1 U720 ( .A(n73), .B(n803), .Y(n669) );
  INVX1 U721 ( .A(n669), .Y(n670) );
  AND2X1 U722 ( .A(n65), .B(n803), .Y(n671) );
  INVX1 U723 ( .A(n671), .Y(n672) );
  INVX8 U724 ( .A(net60296), .Y(net60284) );
  INVX1 U725 ( .A(net60300), .Y(net72479) );
  INVX1 U726 ( .A(net72479), .Y(net72480) );
  MUX2X1 U727 ( .B(n758), .A(n759), .S(net59578), .Y(n767) );
  INVX1 U728 ( .A(net59842), .Y(net72395) );
  MUX2X1 U729 ( .B(\mem<5><0> ), .A(\mem<4><0> ), .S(net72480), .Y(n681) );
  INVX1 U730 ( .A(net60286), .Y(net66027) );
  MUX2X1 U731 ( .B(n706), .A(n707), .S(net59300), .Y(n708) );
  INVX4 U732 ( .A(N11), .Y(net59846) );
  MUX2X1 U733 ( .B(n796), .A(n797), .S(net59428), .Y(n798) );
  INVX8 U734 ( .A(net60296), .Y(net60282) );
  INVX8 U735 ( .A(net60300), .Y(net60292) );
  INVX8 U736 ( .A(net59846), .Y(net59840) );
  INVX8 U737 ( .A(N12), .Y(net59578) );
  INVX8 U738 ( .A(N14), .Y(net59300) );
  MUX2X1 U739 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(net60284), .Y(n679) );
  MUX2X1 U740 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(net101796), .Y(n678) );
  MUX2X1 U741 ( .B(n679), .A(n678), .S(net59842), .Y(n683) );
  MUX2X1 U742 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(net60284), .Y(n680) );
  MUX2X1 U743 ( .B(n681), .A(n680), .S(net59838), .Y(n682) );
  MUX2X1 U744 ( .B(n683), .A(n682), .S(N12), .Y(n691) );
  MUX2X1 U745 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(net60284), .Y(n685) );
  MUX2X1 U746 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(net60286), .Y(n684) );
  MUX2X1 U747 ( .B(n685), .A(n684), .S(net59842), .Y(n689) );
  MUX2X1 U748 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(net60282), .Y(n687) );
  MUX2X1 U749 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(net60282), .Y(n686) );
  MUX2X1 U750 ( .B(n687), .A(n686), .S(net59838), .Y(n688) );
  MUX2X1 U751 ( .B(n689), .A(n688), .S(N12), .Y(n690) );
  MUX2X1 U752 ( .B(n691), .A(n690), .S(net59426), .Y(n707) );
  MUX2X1 U753 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(net60288), .Y(n693) );
  MUX2X1 U754 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(net60292), .Y(n692) );
  MUX2X1 U755 ( .B(n693), .A(n692), .S(net59838), .Y(n697) );
  MUX2X1 U756 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(net60286), .Y(n695) );
  MUX2X1 U757 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(net60292), .Y(n694) );
  MUX2X1 U758 ( .B(n695), .A(n694), .S(net59836), .Y(n696) );
  MUX2X1 U759 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(net60292), .Y(n699) );
  MUX2X1 U760 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(net60292), .Y(n698) );
  MUX2X1 U761 ( .B(n699), .A(n698), .S(net59836), .Y(n703) );
  MUX2X1 U762 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(net60292), .Y(n701) );
  MUX2X1 U763 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(net60292), .Y(n700) );
  MUX2X1 U764 ( .B(n701), .A(n700), .S(net59838), .Y(n702) );
  MUX2X1 U765 ( .B(n703), .A(n702), .S(N12), .Y(n704) );
  MUX2X1 U766 ( .B(n705), .A(n704), .S(net59426), .Y(n706) );
  MUX2X1 U767 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(net60292), .Y(n709) );
  MUX2X1 U768 ( .B(n710), .A(n709), .S(net59836), .Y(n714) );
  MUX2X1 U769 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(net60288), .Y(n712) );
  MUX2X1 U770 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(net60288), .Y(n711) );
  MUX2X1 U771 ( .B(n712), .A(n711), .S(net59838), .Y(n713) );
  MUX2X1 U772 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(net101551), .Y(n716) );
  MUX2X1 U773 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(net60288), .Y(n715) );
  MUX2X1 U774 ( .B(n716), .A(n715), .S(net59838), .Y(n720) );
  MUX2X1 U775 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(net101667), .Y(n718) );
  MUX2X1 U776 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(net60292), .Y(n717) );
  MUX2X1 U777 ( .B(n718), .A(n717), .S(net59836), .Y(n719) );
  MUX2X1 U778 ( .B(n722), .A(n721), .S(net59426), .Y(n738) );
  MUX2X1 U779 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(net101551), .Y(n724) );
  MUX2X1 U780 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(net60282), .Y(n723) );
  MUX2X1 U781 ( .B(n724), .A(n723), .S(net59838), .Y(n728) );
  MUX2X1 U782 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(net101667), .Y(n726) );
  MUX2X1 U783 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(net101667), .Y(n725) );
  MUX2X1 U784 ( .B(n726), .A(n725), .S(net59838), .Y(n727) );
  MUX2X1 U785 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(net60286), .Y(n730) );
  MUX2X1 U786 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(net60286), .Y(n729) );
  MUX2X1 U787 ( .B(n730), .A(n729), .S(net59838), .Y(n734) );
  MUX2X1 U788 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(net60284), .Y(n732) );
  MUX2X1 U789 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(net60284), .Y(n731) );
  MUX2X1 U790 ( .B(n732), .A(n731), .S(net59838), .Y(n733) );
  MUX2X1 U791 ( .B(n734), .A(n733), .S(N12), .Y(n735) );
  MUX2X1 U792 ( .B(n736), .A(n735), .S(net59426), .Y(n737) );
  MUX2X1 U793 ( .B(n738), .A(n737), .S(net59298), .Y(n739) );
  MUX2X1 U794 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(net60282), .Y(n741) );
  MUX2X1 U795 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(net60284), .Y(n740) );
  MUX2X1 U796 ( .B(n741), .A(n740), .S(net59840), .Y(n745) );
  MUX2X1 U797 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(net60282), .Y(n743) );
  MUX2X1 U798 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(net60282), .Y(n742) );
  MUX2X1 U799 ( .B(n743), .A(n742), .S(net59840), .Y(n744) );
  MUX2X1 U800 ( .B(n745), .A(n744), .S(net59576), .Y(n753) );
  MUX2X1 U801 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(net60282), .Y(n747) );
  MUX2X1 U802 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(net60282), .Y(n746) );
  MUX2X1 U803 ( .B(n747), .A(n746), .S(net59840), .Y(n751) );
  MUX2X1 U804 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(net60284), .Y(n749) );
  MUX2X1 U805 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(net60284), .Y(n748) );
  MUX2X1 U806 ( .B(n749), .A(n748), .S(net59840), .Y(n750) );
  MUX2X1 U807 ( .B(n751), .A(n750), .S(net59576), .Y(n752) );
  MUX2X1 U808 ( .B(n753), .A(n752), .S(net59426), .Y(n769) );
  MUX2X1 U809 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(net101551), .Y(n755) );
  MUX2X1 U810 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(net60284), .Y(n754) );
  MUX2X1 U811 ( .B(n755), .A(n754), .S(net59840), .Y(n759) );
  MUX2X1 U812 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(net60286), .Y(n757) );
  MUX2X1 U813 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(net60286), .Y(n756) );
  MUX2X1 U814 ( .B(n757), .A(n756), .S(net59840), .Y(n758) );
  MUX2X1 U815 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(net60286), .Y(n761) );
  MUX2X1 U816 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(net60286), .Y(n760) );
  MUX2X1 U817 ( .B(n761), .A(n760), .S(net59840), .Y(n765) );
  MUX2X1 U818 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(net60282), .Y(n763) );
  MUX2X1 U819 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(net101667), .Y(n762) );
  MUX2X1 U820 ( .B(n763), .A(n762), .S(net59840), .Y(n764) );
  MUX2X1 U821 ( .B(n765), .A(n764), .S(net59576), .Y(n766) );
  MUX2X1 U822 ( .B(n767), .A(n766), .S(net59426), .Y(n768) );
  MUX2X1 U823 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(net60284), .Y(n772) );
  MUX2X1 U824 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(net101711), .Y(n771) );
  MUX2X1 U825 ( .B(n772), .A(n771), .S(net59840), .Y(n776) );
  MUX2X1 U826 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(net60284), .Y(n774) );
  MUX2X1 U827 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(net101711), .Y(n773) );
  MUX2X1 U828 ( .B(n774), .A(n773), .S(net59840), .Y(n775) );
  MUX2X1 U829 ( .B(n776), .A(n775), .S(net59576), .Y(n784) );
  MUX2X1 U830 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(net60282), .Y(n778) );
  MUX2X1 U831 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(net60284), .Y(n777) );
  MUX2X1 U832 ( .B(n778), .A(n777), .S(net59840), .Y(n782) );
  MUX2X1 U833 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(net60282), .Y(n780) );
  MUX2X1 U834 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(net60282), .Y(n779) );
  MUX2X1 U835 ( .B(n780), .A(n779), .S(net59840), .Y(n781) );
  MUX2X1 U836 ( .B(n782), .A(n781), .S(net59576), .Y(n783) );
  MUX2X1 U837 ( .B(n784), .A(n783), .S(net59426), .Y(n799) );
  MUX2X1 U838 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(net60282), .Y(n786) );
  MUX2X1 U839 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(net60282), .Y(n785) );
  MUX2X1 U840 ( .B(n786), .A(n785), .S(net59838), .Y(n790) );
  MUX2X1 U841 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(net60282), .Y(n788) );
  MUX2X1 U842 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(net60282), .Y(n787) );
  MUX2X1 U843 ( .B(n788), .A(n787), .S(net59838), .Y(n789) );
  MUX2X1 U844 ( .B(n790), .A(n789), .S(net59576), .Y(n797) );
  MUX2X1 U845 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(net60284), .Y(n792) );
  MUX2X1 U846 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(net60284), .Y(n791) );
  MUX2X1 U847 ( .B(n792), .A(n791), .S(net59838), .Y(n795) );
  MUX2X1 U848 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(net60284), .Y(n794) );
  MUX2X1 U849 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(net60282), .Y(n793) );
  MUX2X1 U850 ( .B(n795), .A(n37), .S(net59576), .Y(n796) );
endmodule


module memc_Size1_1 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n92), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n91), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n90), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n89), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n88), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n87), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n86), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n85), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n84), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n83), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n82), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n81), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n80), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n79), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n78), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n77), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n76), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n75), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n74), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n73), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n72), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n71), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n70), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n69), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n68), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n67), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n66), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n65), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n64), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n63), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n62), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n61), .CLK(clk), .Q(\mem<31><0> ) );
  INVX2 U2 ( .A(n193), .Y(n3) );
  INVX1 U3 ( .A(n158), .Y(N17) );
  INVX1 U4 ( .A(rst), .Y(n174) );
  INVX1 U5 ( .A(n167), .Y(n159) );
  INVX1 U6 ( .A(N12), .Y(n169) );
  INVX2 U7 ( .A(n122), .Y(n123) );
  INVX1 U8 ( .A(n108), .Y(n204) );
  INVX1 U9 ( .A(n109), .Y(n207) );
  INVX2 U10 ( .A(n165), .Y(n160) );
  AND2X1 U11 ( .A(n165), .B(n99), .Y(n119) );
  INVX1 U12 ( .A(n9), .Y(n1) );
  INVX1 U13 ( .A(n126), .Y(n2) );
  INVX2 U14 ( .A(n126), .Y(n127) );
  INVX4 U15 ( .A(n97), .Y(n163) );
  AND2X2 U16 ( .A(n5), .B(\data_in<0> ), .Y(n105) );
  INVX1 U17 ( .A(n7), .Y(n4) );
  INVX1 U18 ( .A(n11), .Y(n5) );
  INVX1 U19 ( .A(n193), .Y(n6) );
  INVX1 U20 ( .A(n9), .Y(n193) );
  AND2X2 U21 ( .A(n1), .B(\data_in<0> ), .Y(n104) );
  AND2X2 U22 ( .A(\data_in<0> ), .B(n4), .Y(n103) );
  AND2X2 U23 ( .A(\data_in<0> ), .B(n161), .Y(n97) );
  OR2X2 U24 ( .A(n173), .B(n8), .Y(n7) );
  OR2X2 U25 ( .A(n124), .B(n14), .Y(n8) );
  OR2X2 U26 ( .A(n171), .B(n10), .Y(n9) );
  OR2X2 U27 ( .A(n125), .B(n14), .Y(n10) );
  OR2X2 U28 ( .A(n124), .B(n10), .Y(n11) );
  OR2X2 U29 ( .A(write), .B(n101), .Y(n12) );
  INVX1 U30 ( .A(n12), .Y(\data_out<0> ) );
  OR2X2 U31 ( .A(n96), .B(\addr<5> ), .Y(n14) );
  INVX1 U32 ( .A(n14), .Y(n15) );
  AND2X2 U33 ( .A(n120), .B(n103), .Y(n16) );
  INVX1 U34 ( .A(n16), .Y(n17) );
  AND2X2 U35 ( .A(n117), .B(n103), .Y(n18) );
  INVX1 U36 ( .A(n18), .Y(n19) );
  AND2X2 U37 ( .A(n204), .B(n103), .Y(n20) );
  INVX1 U38 ( .A(n20), .Y(n21) );
  AND2X2 U39 ( .A(n207), .B(n103), .Y(n22) );
  INVX1 U40 ( .A(n22), .Y(n23) );
  AND2X2 U41 ( .A(n110), .B(n103), .Y(n24) );
  INVX1 U42 ( .A(n24), .Y(n25) );
  AND2X2 U43 ( .A(n112), .B(n103), .Y(n26) );
  INVX1 U44 ( .A(n26), .Y(n27) );
  AND2X2 U45 ( .A(n114), .B(n103), .Y(n28) );
  INVX1 U46 ( .A(n28), .Y(n29) );
  AND2X2 U47 ( .A(n119), .B(n103), .Y(n30) );
  INVX1 U48 ( .A(n30), .Y(n31) );
  AND2X2 U49 ( .A(n120), .B(n104), .Y(n32) );
  INVX1 U50 ( .A(n32), .Y(n33) );
  AND2X2 U51 ( .A(n117), .B(n104), .Y(n34) );
  INVX1 U52 ( .A(n34), .Y(n35) );
  AND2X2 U53 ( .A(n204), .B(n104), .Y(n36) );
  INVX1 U54 ( .A(n36), .Y(n37) );
  AND2X2 U55 ( .A(n207), .B(n104), .Y(n38) );
  INVX1 U56 ( .A(n38), .Y(n39) );
  AND2X2 U57 ( .A(n110), .B(n104), .Y(n40) );
  INVX1 U58 ( .A(n40), .Y(n41) );
  AND2X2 U59 ( .A(n112), .B(n104), .Y(n42) );
  INVX1 U60 ( .A(n42), .Y(n43) );
  AND2X2 U61 ( .A(n104), .B(n114), .Y(n44) );
  INVX1 U62 ( .A(n44), .Y(n45) );
  AND2X2 U63 ( .A(n119), .B(n104), .Y(n46) );
  INVX1 U64 ( .A(n46), .Y(n47) );
  AND2X2 U65 ( .A(n120), .B(n105), .Y(n48) );
  INVX1 U66 ( .A(n48), .Y(n49) );
  AND2X2 U67 ( .A(n117), .B(n105), .Y(n50) );
  INVX1 U68 ( .A(n50), .Y(n51) );
  AND2X2 U69 ( .A(n204), .B(n105), .Y(n52) );
  INVX1 U70 ( .A(n52), .Y(n53) );
  AND2X2 U71 ( .A(n207), .B(n105), .Y(n54) );
  INVX1 U72 ( .A(n54), .Y(n55) );
  AND2X2 U73 ( .A(n110), .B(n105), .Y(n56) );
  INVX1 U74 ( .A(n56), .Y(n57) );
  AND2X2 U75 ( .A(n112), .B(n105), .Y(n58) );
  INVX1 U76 ( .A(n58), .Y(n59) );
  AND2X2 U77 ( .A(n114), .B(n105), .Y(n60) );
  INVX1 U78 ( .A(n60), .Y(n93) );
  AND2X2 U79 ( .A(n119), .B(n105), .Y(n94) );
  INVX1 U80 ( .A(n94), .Y(n95) );
  BUFX2 U81 ( .A(n175), .Y(n96) );
  INVX1 U82 ( .A(n169), .Y(n168) );
  INVX1 U83 ( .A(n167), .Y(n166) );
  INVX1 U84 ( .A(n165), .Y(n164) );
  OR2X1 U85 ( .A(n166), .B(n168), .Y(n98) );
  INVX1 U86 ( .A(n98), .Y(n99) );
  AND2X1 U87 ( .A(N17), .B(n174), .Y(n100) );
  INVX1 U88 ( .A(n100), .Y(n101) );
  AND2X1 U89 ( .A(n168), .B(n166), .Y(n102) );
  OR2X1 U90 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n106) );
  INVX1 U91 ( .A(n106), .Y(n107) );
  BUFX2 U92 ( .A(n205), .Y(n108) );
  BUFX2 U93 ( .A(n208), .Y(n109) );
  INVX1 U94 ( .A(n111), .Y(n110) );
  BUFX2 U95 ( .A(n210), .Y(n111) );
  INVX1 U96 ( .A(n113), .Y(n112) );
  BUFX2 U97 ( .A(n212), .Y(n113) );
  INVX1 U98 ( .A(n115), .Y(n114) );
  BUFX2 U99 ( .A(n214), .Y(n115) );
  INVX1 U100 ( .A(n117), .Y(n116) );
  AND2X1 U101 ( .A(n165), .B(n102), .Y(n117) );
  INVX1 U102 ( .A(n119), .Y(n118) );
  AND2X1 U103 ( .A(n164), .B(n102), .Y(n120) );
  INVX1 U104 ( .A(n120), .Y(n121) );
  INVX1 U105 ( .A(n7), .Y(n122) );
  INVX1 U106 ( .A(n171), .Y(n124) );
  INVX1 U107 ( .A(n173), .Y(n172) );
  INVX1 U108 ( .A(n173), .Y(n125) );
  INVX1 U109 ( .A(n171), .Y(n170) );
  INVX1 U110 ( .A(n11), .Y(n126) );
  INVX1 U111 ( .A(N13), .Y(n171) );
  INVX1 U112 ( .A(N14), .Y(n173) );
  MUX2X1 U113 ( .B(n129), .A(n130), .S(n159), .Y(n128) );
  MUX2X1 U114 ( .B(n132), .A(n133), .S(n159), .Y(n131) );
  MUX2X1 U115 ( .B(n135), .A(n136), .S(n159), .Y(n134) );
  MUX2X1 U116 ( .B(n138), .A(n139), .S(n159), .Y(n137) );
  MUX2X1 U117 ( .B(n141), .A(n142), .S(n170), .Y(n140) );
  MUX2X1 U118 ( .B(n144), .A(n145), .S(n159), .Y(n143) );
  MUX2X1 U119 ( .B(n147), .A(n148), .S(n159), .Y(n146) );
  MUX2X1 U120 ( .B(n150), .A(n151), .S(n159), .Y(n149) );
  MUX2X1 U121 ( .B(n153), .A(n154), .S(n159), .Y(n152) );
  MUX2X1 U122 ( .B(n156), .A(n157), .S(n170), .Y(n155) );
  MUX2X1 U123 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n160), .Y(n130) );
  MUX2X1 U124 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n160), .Y(n129) );
  MUX2X1 U125 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n160), .Y(n133) );
  MUX2X1 U126 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n160), .Y(n132) );
  MUX2X1 U127 ( .B(n131), .A(n128), .S(n168), .Y(n142) );
  MUX2X1 U128 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n160), .Y(n136) );
  MUX2X1 U129 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n160), .Y(n135) );
  MUX2X1 U130 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n160), .Y(n139) );
  MUX2X1 U131 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n160), .Y(n138) );
  MUX2X1 U132 ( .B(n137), .A(n134), .S(n168), .Y(n141) );
  MUX2X1 U133 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n160), .Y(n145) );
  MUX2X1 U134 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n160), .Y(n144) );
  MUX2X1 U135 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n160), .Y(n148) );
  MUX2X1 U136 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n160), .Y(n147) );
  MUX2X1 U137 ( .B(n146), .A(n143), .S(n168), .Y(n157) );
  MUX2X1 U138 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n160), .Y(n151) );
  MUX2X1 U139 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n160), .Y(n150) );
  MUX2X1 U140 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n160), .Y(n154) );
  MUX2X1 U141 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n160), .Y(n153) );
  MUX2X1 U142 ( .B(n152), .A(n149), .S(n168), .Y(n156) );
  MUX2X1 U143 ( .B(n155), .A(n140), .S(n172), .Y(n158) );
  INVX1 U144 ( .A(N11), .Y(n167) );
  INVX1 U145 ( .A(n183), .Y(n161) );
  INVX1 U146 ( .A(n161), .Y(n162) );
  INVX1 U147 ( .A(N10), .Y(n165) );
  NAND3X1 U148 ( .A(n107), .B(n174), .C(write), .Y(n175) );
  NAND3X1 U149 ( .A(n172), .B(n170), .C(n15), .Y(n183) );
  OAI21X1 U150 ( .A(n162), .B(n121), .C(\mem<31><0> ), .Y(n176) );
  OAI21X1 U151 ( .A(n163), .B(n121), .C(n176), .Y(n61) );
  OAI21X1 U152 ( .A(n116), .B(n162), .C(\mem<30><0> ), .Y(n177) );
  OAI21X1 U153 ( .A(n116), .B(n163), .C(n177), .Y(n62) );
  NAND3X1 U154 ( .A(n164), .B(n168), .C(n167), .Y(n205) );
  OAI21X1 U155 ( .A(n108), .B(n162), .C(\mem<29><0> ), .Y(n178) );
  OAI21X1 U156 ( .A(n108), .B(n163), .C(n178), .Y(n63) );
  NAND3X1 U157 ( .A(n168), .B(n167), .C(n165), .Y(n208) );
  OAI21X1 U158 ( .A(n109), .B(n162), .C(\mem<28><0> ), .Y(n179) );
  OAI21X1 U159 ( .A(n109), .B(n163), .C(n179), .Y(n64) );
  NAND3X1 U160 ( .A(n164), .B(n166), .C(n169), .Y(n210) );
  OAI21X1 U161 ( .A(n111), .B(n162), .C(\mem<27><0> ), .Y(n180) );
  OAI21X1 U162 ( .A(n111), .B(n163), .C(n180), .Y(n65) );
  NAND3X1 U163 ( .A(n169), .B(n166), .C(n165), .Y(n212) );
  OAI21X1 U164 ( .A(n113), .B(n162), .C(\mem<26><0> ), .Y(n181) );
  OAI21X1 U165 ( .A(n113), .B(n163), .C(n181), .Y(n66) );
  NAND3X1 U166 ( .A(n164), .B(n169), .C(n167), .Y(n214) );
  OAI21X1 U167 ( .A(n115), .B(n162), .C(\mem<25><0> ), .Y(n182) );
  OAI21X1 U168 ( .A(n115), .B(n163), .C(n182), .Y(n67) );
  OAI21X1 U169 ( .A(n118), .B(n162), .C(\mem<24><0> ), .Y(n184) );
  OAI21X1 U170 ( .A(n118), .B(n163), .C(n184), .Y(n68) );
  OAI21X1 U171 ( .A(n123), .B(n121), .C(\mem<23><0> ), .Y(n185) );
  NAND2X1 U172 ( .A(n17), .B(n185), .Y(n69) );
  OAI21X1 U173 ( .A(n123), .B(n116), .C(\mem<22><0> ), .Y(n186) );
  NAND2X1 U174 ( .A(n19), .B(n186), .Y(n70) );
  OAI21X1 U175 ( .A(n123), .B(n108), .C(\mem<21><0> ), .Y(n187) );
  NAND2X1 U176 ( .A(n21), .B(n187), .Y(n71) );
  OAI21X1 U177 ( .A(n123), .B(n109), .C(\mem<20><0> ), .Y(n188) );
  NAND2X1 U178 ( .A(n23), .B(n188), .Y(n72) );
  OAI21X1 U179 ( .A(n123), .B(n111), .C(\mem<19><0> ), .Y(n189) );
  NAND2X1 U180 ( .A(n25), .B(n189), .Y(n73) );
  OAI21X1 U181 ( .A(n123), .B(n113), .C(\mem<18><0> ), .Y(n190) );
  NAND2X1 U182 ( .A(n27), .B(n190), .Y(n74) );
  OAI21X1 U183 ( .A(n123), .B(n115), .C(\mem<17><0> ), .Y(n191) );
  NAND2X1 U184 ( .A(n29), .B(n191), .Y(n75) );
  OAI21X1 U185 ( .A(n123), .B(n118), .C(\mem<16><0> ), .Y(n192) );
  NAND2X1 U186 ( .A(n31), .B(n192), .Y(n76) );
  OAI21X1 U187 ( .A(n6), .B(n121), .C(\mem<15><0> ), .Y(n194) );
  NAND2X1 U188 ( .A(n33), .B(n194), .Y(n77) );
  OAI21X1 U189 ( .A(n6), .B(n116), .C(\mem<14><0> ), .Y(n195) );
  NAND2X1 U190 ( .A(n35), .B(n195), .Y(n78) );
  OAI21X1 U191 ( .A(n3), .B(n108), .C(\mem<13><0> ), .Y(n196) );
  NAND2X1 U192 ( .A(n37), .B(n196), .Y(n79) );
  OAI21X1 U193 ( .A(n3), .B(n109), .C(\mem<12><0> ), .Y(n197) );
  NAND2X1 U194 ( .A(n39), .B(n197), .Y(n80) );
  OAI21X1 U195 ( .A(n3), .B(n111), .C(\mem<11><0> ), .Y(n198) );
  NAND2X1 U196 ( .A(n41), .B(n198), .Y(n81) );
  OAI21X1 U197 ( .A(n3), .B(n113), .C(\mem<10><0> ), .Y(n199) );
  NAND2X1 U198 ( .A(n43), .B(n199), .Y(n82) );
  OAI21X1 U199 ( .A(n6), .B(n115), .C(\mem<9><0> ), .Y(n200) );
  NAND2X1 U200 ( .A(n45), .B(n200), .Y(n83) );
  OAI21X1 U201 ( .A(n3), .B(n118), .C(\mem<8><0> ), .Y(n201) );
  NAND2X1 U202 ( .A(n47), .B(n201), .Y(n84) );
  OAI21X1 U203 ( .A(n127), .B(n121), .C(\mem<7><0> ), .Y(n202) );
  NAND2X1 U204 ( .A(n49), .B(n202), .Y(n85) );
  OAI21X1 U205 ( .A(n127), .B(n116), .C(\mem<6><0> ), .Y(n203) );
  NAND2X1 U206 ( .A(n51), .B(n203), .Y(n86) );
  OAI21X1 U207 ( .A(n127), .B(n108), .C(\mem<5><0> ), .Y(n206) );
  NAND2X1 U208 ( .A(n53), .B(n206), .Y(n87) );
  OAI21X1 U209 ( .A(n127), .B(n109), .C(\mem<4><0> ), .Y(n209) );
  NAND2X1 U210 ( .A(n55), .B(n209), .Y(n88) );
  OAI21X1 U211 ( .A(n2), .B(n111), .C(\mem<3><0> ), .Y(n211) );
  NAND2X1 U212 ( .A(n57), .B(n211), .Y(n89) );
  OAI21X1 U213 ( .A(n127), .B(n113), .C(\mem<2><0> ), .Y(n213) );
  NAND2X1 U214 ( .A(n59), .B(n213), .Y(n90) );
  OAI21X1 U215 ( .A(n127), .B(n115), .C(\mem<1><0> ), .Y(n215) );
  NAND2X1 U216 ( .A(n93), .B(n215), .Y(n91) );
  OAI21X1 U217 ( .A(n2), .B(n118), .C(\mem<0><0> ), .Y(n216) );
  NAND2X1 U218 ( .A(n95), .B(n216), .Y(n92) );
endmodule


module memv_1 ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , n42, n46, n49, n52, n55, n58, n61, n64, n67, n70, n73,
         n76, n79, n82, n85, n88, n90, n91, n92, n94, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n113, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n132, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n151,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n170, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n206, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n224, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n243, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n261, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n279, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n297, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n334, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n352, n355, n356, n357, n358, n359, n361, n363, n364, n365, n366,
         n367, n368, n370, n371, n372, n373, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43,
         n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62, n63,
         n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83, n84,
         n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149, n150,
         n152, n169, n171, n187, n189, n205, n207, n223, n225, n241, n242,
         n244, n260, n262, n278, n280, n296, n298, n314, n315, n317, n333,
         n335, n351, n353, n354, n360, n362, n369, n374, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n633), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n632), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n631), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n630), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n629), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n628), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n627), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n626), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n625), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n624), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n623), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n622), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n621), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n620), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n619), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n618), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n617), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n616), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n615), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n614), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n613), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n612), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n611), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n610), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n609), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n608), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n607), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n606), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n605), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n604), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n603), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n602), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n601), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n600), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n599), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n598), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n597), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n596), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n595), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n594), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n593), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n592), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n591), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n590), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n589), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n588), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n587), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n586), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n585), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n584), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n583), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n582), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n581), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n580), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n579), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n578), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n577), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n576), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n575), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n574), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n573), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n572), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n571), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n570), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n569), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n568), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n567), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n566), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n565), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n564), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n563), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n562), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n561), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n560), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n559), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n558), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n557), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n556), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n555), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n554), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n553), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n552), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n551), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n550), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n549), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n548), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n547), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n546), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n545), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n544), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n543), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n542), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n541), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n540), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n539), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n538), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n537), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n536), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n535), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n534), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n533), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n532), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n531), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n530), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n529), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n528), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n527), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n526), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n525), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n524), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n523), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n522), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n521), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n520), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n519), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n518), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n517), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n516), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n515), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n514), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n513), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n512), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n511), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n510), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n509), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n508), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n507), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n506), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n505), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n504), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n503), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n502), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n501), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n500), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n499), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n498), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n497), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n496), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n495), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n494), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n493), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n492), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n491), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n490), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n489), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n488), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n487), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n486), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n485), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n484), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n483), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n482), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n481), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n480), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n479), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n478), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n477), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n476), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n475), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n474), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n473), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n472), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n471), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n470), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n469), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n468), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n467), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n466), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n465), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n464), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n463), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n462), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n461), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n460), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n459), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n458), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n457), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n456), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n455), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n454), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n453), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n452), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n451), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n450), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n449), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n448), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n447), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n446), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n445), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n444), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n443), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n442), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n441), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n440), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n439), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n438), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n437), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n436), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n435), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n434), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n433), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n432), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n431), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n430), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n429), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n428), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n427), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n426), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n425), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n424), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n423), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n422), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n421), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n420), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n419), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n418), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n417), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n416), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n415), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n414), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n413), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n412), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n411), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n410), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n409), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n408), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n407), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n406), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n405), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n404), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n403), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n402), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n401), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n400), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n399), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n398), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n397), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n396), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n395), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n394), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n393), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n392), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n391), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n390), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n389), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n388), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n387), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n386), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n385), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n384), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n383), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n382), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n381), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n380), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n379), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n378), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U6 ( .A(N21), .B(n757), .Y(n355) );
  AND2X2 U7 ( .A(N21), .B(n758), .Y(n364) );
  AND2X2 U8 ( .A(n752), .B(n744), .Y(n356) );
  AND2X2 U9 ( .A(n752), .B(n746), .Y(n358) );
  OAI21X1 U49 ( .A(n133), .B(n729), .C(n42), .Y(n378) );
  OAI21X1 U50 ( .A(n45), .B(n727), .C(\mem<255> ), .Y(n42) );
  OAI21X1 U51 ( .A(n730), .B(n130), .C(n46), .Y(n379) );
  OAI21X1 U52 ( .A(n728), .B(n43), .C(\mem<254> ), .Y(n46) );
  OAI21X1 U53 ( .A(n730), .B(n679), .C(n49), .Y(n380) );
  OAI21X1 U54 ( .A(n728), .B(n40), .C(\mem<253> ), .Y(n49) );
  OAI21X1 U55 ( .A(n730), .B(n678), .C(n52), .Y(n381) );
  OAI21X1 U56 ( .A(n728), .B(n38), .C(\mem<252> ), .Y(n52) );
  OAI21X1 U57 ( .A(n730), .B(n112), .C(n55), .Y(n382) );
  OAI21X1 U58 ( .A(n728), .B(n36), .C(\mem<251> ), .Y(n55) );
  OAI21X1 U59 ( .A(n730), .B(n93), .C(n58), .Y(n383) );
  OAI21X1 U60 ( .A(n728), .B(n34), .C(\mem<250> ), .Y(n58) );
  OAI21X1 U61 ( .A(n730), .B(n87), .C(n61), .Y(n384) );
  OAI21X1 U62 ( .A(n728), .B(n32), .C(\mem<249> ), .Y(n61) );
  OAI21X1 U63 ( .A(n730), .B(n84), .C(n64), .Y(n385) );
  OAI21X1 U64 ( .A(n728), .B(n30), .C(\mem<248> ), .Y(n64) );
  OAI21X1 U65 ( .A(n730), .B(n677), .C(n67), .Y(n386) );
  OAI21X1 U66 ( .A(n728), .B(n28), .C(\mem<247> ), .Y(n67) );
  OAI21X1 U67 ( .A(n729), .B(n676), .C(n70), .Y(n387) );
  OAI21X1 U68 ( .A(n727), .B(n26), .C(\mem<246> ), .Y(n70) );
  OAI21X1 U69 ( .A(n729), .B(n675), .C(n73), .Y(n388) );
  OAI21X1 U70 ( .A(n727), .B(n24), .C(\mem<245> ), .Y(n73) );
  OAI21X1 U71 ( .A(n729), .B(n674), .C(n76), .Y(n389) );
  OAI21X1 U72 ( .A(n727), .B(n22), .C(\mem<244> ), .Y(n76) );
  OAI21X1 U73 ( .A(n729), .B(n673), .C(n79), .Y(n390) );
  OAI21X1 U74 ( .A(n727), .B(n20), .C(\mem<243> ), .Y(n79) );
  OAI21X1 U75 ( .A(n729), .B(n672), .C(n82), .Y(n391) );
  OAI21X1 U76 ( .A(n727), .B(n18), .C(\mem<242> ), .Y(n82) );
  OAI21X1 U77 ( .A(n729), .B(n671), .C(n85), .Y(n392) );
  OAI21X1 U78 ( .A(n727), .B(n16), .C(\mem<241> ), .Y(n85) );
  OAI21X1 U79 ( .A(n729), .B(n665), .C(n88), .Y(n393) );
  OAI21X1 U80 ( .A(n727), .B(n14), .C(\mem<240> ), .Y(n88) );
  OAI21X1 U83 ( .A(n133), .B(n726), .C(n94), .Y(n394) );
  OAI21X1 U84 ( .A(n45), .B(n724), .C(\mem<239> ), .Y(n94) );
  OAI21X1 U85 ( .A(n130), .B(n726), .C(n96), .Y(n395) );
  OAI21X1 U86 ( .A(n43), .B(n724), .C(\mem<238> ), .Y(n96) );
  OAI21X1 U87 ( .A(n679), .B(n726), .C(n97), .Y(n396) );
  OAI21X1 U88 ( .A(n40), .B(n724), .C(\mem<237> ), .Y(n97) );
  OAI21X1 U89 ( .A(n678), .B(n726), .C(n98), .Y(n397) );
  OAI21X1 U90 ( .A(n38), .B(n724), .C(\mem<236> ), .Y(n98) );
  OAI21X1 U91 ( .A(n112), .B(n726), .C(n99), .Y(n398) );
  OAI21X1 U92 ( .A(n36), .B(n724), .C(\mem<235> ), .Y(n99) );
  OAI21X1 U93 ( .A(n93), .B(n726), .C(n100), .Y(n399) );
  OAI21X1 U94 ( .A(n34), .B(n724), .C(\mem<234> ), .Y(n100) );
  OAI21X1 U95 ( .A(n87), .B(n726), .C(n101), .Y(n400) );
  OAI21X1 U96 ( .A(n32), .B(n724), .C(\mem<233> ), .Y(n101) );
  OAI21X1 U97 ( .A(n84), .B(n726), .C(n102), .Y(n401) );
  OAI21X1 U98 ( .A(n30), .B(n724), .C(\mem<232> ), .Y(n102) );
  OAI21X1 U99 ( .A(n677), .B(n725), .C(n103), .Y(n402) );
  OAI21X1 U100 ( .A(n28), .B(n723), .C(\mem<231> ), .Y(n103) );
  OAI21X1 U101 ( .A(n676), .B(n725), .C(n104), .Y(n403) );
  OAI21X1 U102 ( .A(n26), .B(n723), .C(\mem<230> ), .Y(n104) );
  OAI21X1 U103 ( .A(n675), .B(n725), .C(n105), .Y(n404) );
  OAI21X1 U104 ( .A(n24), .B(n723), .C(\mem<229> ), .Y(n105) );
  OAI21X1 U105 ( .A(n674), .B(n725), .C(n106), .Y(n405) );
  OAI21X1 U106 ( .A(n22), .B(n723), .C(\mem<228> ), .Y(n106) );
  OAI21X1 U107 ( .A(n673), .B(n725), .C(n107), .Y(n406) );
  OAI21X1 U108 ( .A(n20), .B(n723), .C(\mem<227> ), .Y(n107) );
  OAI21X1 U109 ( .A(n672), .B(n725), .C(n108), .Y(n407) );
  OAI21X1 U110 ( .A(n18), .B(n723), .C(\mem<226> ), .Y(n108) );
  OAI21X1 U111 ( .A(n671), .B(n725), .C(n109), .Y(n408) );
  OAI21X1 U112 ( .A(n16), .B(n723), .C(\mem<225> ), .Y(n109) );
  OAI21X1 U113 ( .A(n665), .B(n725), .C(n110), .Y(n409) );
  OAI21X1 U114 ( .A(n14), .B(n723), .C(\mem<224> ), .Y(n110) );
  OAI21X1 U117 ( .A(n133), .B(n722), .C(n113), .Y(n410) );
  OAI21X1 U118 ( .A(n45), .B(n720), .C(\mem<223> ), .Y(n113) );
  OAI21X1 U119 ( .A(n130), .B(n722), .C(n115), .Y(n411) );
  OAI21X1 U120 ( .A(n43), .B(n720), .C(\mem<222> ), .Y(n115) );
  OAI21X1 U121 ( .A(n679), .B(n722), .C(n116), .Y(n412) );
  OAI21X1 U122 ( .A(n40), .B(n720), .C(\mem<221> ), .Y(n116) );
  OAI21X1 U123 ( .A(n678), .B(n722), .C(n117), .Y(n413) );
  OAI21X1 U124 ( .A(n38), .B(n720), .C(\mem<220> ), .Y(n117) );
  OAI21X1 U125 ( .A(n112), .B(n722), .C(n118), .Y(n414) );
  OAI21X1 U126 ( .A(n36), .B(n720), .C(\mem<219> ), .Y(n118) );
  OAI21X1 U127 ( .A(n93), .B(n722), .C(n119), .Y(n415) );
  OAI21X1 U128 ( .A(n34), .B(n720), .C(\mem<218> ), .Y(n119) );
  OAI21X1 U129 ( .A(n87), .B(n722), .C(n120), .Y(n416) );
  OAI21X1 U130 ( .A(n32), .B(n720), .C(\mem<217> ), .Y(n120) );
  OAI21X1 U131 ( .A(n84), .B(n722), .C(n121), .Y(n417) );
  OAI21X1 U132 ( .A(n30), .B(n720), .C(\mem<216> ), .Y(n121) );
  OAI21X1 U133 ( .A(n677), .B(n721), .C(n122), .Y(n418) );
  OAI21X1 U134 ( .A(n28), .B(n720), .C(\mem<215> ), .Y(n122) );
  OAI21X1 U135 ( .A(n676), .B(n721), .C(n123), .Y(n419) );
  OAI21X1 U136 ( .A(n26), .B(n720), .C(\mem<214> ), .Y(n123) );
  OAI21X1 U137 ( .A(n675), .B(n721), .C(n124), .Y(n420) );
  OAI21X1 U138 ( .A(n24), .B(n720), .C(\mem<213> ), .Y(n124) );
  OAI21X1 U139 ( .A(n674), .B(n721), .C(n125), .Y(n421) );
  OAI21X1 U140 ( .A(n22), .B(n720), .C(\mem<212> ), .Y(n125) );
  OAI21X1 U141 ( .A(n673), .B(n721), .C(n126), .Y(n422) );
  OAI21X1 U142 ( .A(n20), .B(n720), .C(\mem<211> ), .Y(n126) );
  OAI21X1 U143 ( .A(n672), .B(n721), .C(n127), .Y(n423) );
  OAI21X1 U144 ( .A(n18), .B(n720), .C(\mem<210> ), .Y(n127) );
  OAI21X1 U145 ( .A(n671), .B(n721), .C(n128), .Y(n424) );
  OAI21X1 U146 ( .A(n16), .B(n720), .C(\mem<209> ), .Y(n128) );
  OAI21X1 U147 ( .A(n665), .B(n721), .C(n129), .Y(n425) );
  OAI21X1 U148 ( .A(n14), .B(n720), .C(\mem<208> ), .Y(n129) );
  OAI21X1 U151 ( .A(n133), .B(n719), .C(n132), .Y(n426) );
  OAI21X1 U152 ( .A(n45), .B(n717), .C(\mem<207> ), .Y(n132) );
  OAI21X1 U153 ( .A(n130), .B(n719), .C(n134), .Y(n427) );
  OAI21X1 U154 ( .A(n43), .B(n717), .C(\mem<206> ), .Y(n134) );
  OAI21X1 U155 ( .A(n679), .B(n719), .C(n135), .Y(n428) );
  OAI21X1 U156 ( .A(n40), .B(n717), .C(\mem<205> ), .Y(n135) );
  OAI21X1 U157 ( .A(n678), .B(n719), .C(n136), .Y(n429) );
  OAI21X1 U158 ( .A(n38), .B(n717), .C(\mem<204> ), .Y(n136) );
  OAI21X1 U159 ( .A(n112), .B(n719), .C(n137), .Y(n430) );
  OAI21X1 U160 ( .A(n36), .B(n717), .C(\mem<203> ), .Y(n137) );
  OAI21X1 U161 ( .A(n93), .B(n719), .C(n138), .Y(n431) );
  OAI21X1 U162 ( .A(n34), .B(n717), .C(\mem<202> ), .Y(n138) );
  OAI21X1 U163 ( .A(n87), .B(n719), .C(n139), .Y(n432) );
  OAI21X1 U164 ( .A(n32), .B(n717), .C(\mem<201> ), .Y(n139) );
  OAI21X1 U165 ( .A(n84), .B(n719), .C(n140), .Y(n433) );
  OAI21X1 U166 ( .A(n30), .B(n717), .C(\mem<200> ), .Y(n140) );
  OAI21X1 U167 ( .A(n677), .B(n718), .C(n141), .Y(n434) );
  OAI21X1 U168 ( .A(n28), .B(n717), .C(\mem<199> ), .Y(n141) );
  OAI21X1 U169 ( .A(n676), .B(n718), .C(n142), .Y(n435) );
  OAI21X1 U170 ( .A(n26), .B(n717), .C(\mem<198> ), .Y(n142) );
  OAI21X1 U171 ( .A(n675), .B(n718), .C(n143), .Y(n436) );
  OAI21X1 U172 ( .A(n24), .B(n717), .C(\mem<197> ), .Y(n143) );
  OAI21X1 U173 ( .A(n674), .B(n718), .C(n144), .Y(n437) );
  OAI21X1 U174 ( .A(n22), .B(n717), .C(\mem<196> ), .Y(n144) );
  OAI21X1 U175 ( .A(n673), .B(n718), .C(n145), .Y(n438) );
  OAI21X1 U176 ( .A(n20), .B(n717), .C(\mem<195> ), .Y(n145) );
  OAI21X1 U177 ( .A(n672), .B(n718), .C(n146), .Y(n439) );
  OAI21X1 U178 ( .A(n18), .B(n717), .C(\mem<194> ), .Y(n146) );
  OAI21X1 U179 ( .A(n671), .B(n718), .C(n147), .Y(n440) );
  OAI21X1 U180 ( .A(n16), .B(n717), .C(\mem<193> ), .Y(n147) );
  OAI21X1 U181 ( .A(n665), .B(n718), .C(n148), .Y(n441) );
  OAI21X1 U182 ( .A(n14), .B(n717), .C(\mem<192> ), .Y(n148) );
  OAI21X1 U185 ( .A(n133), .B(n716), .C(n151), .Y(n442) );
  OAI21X1 U186 ( .A(n45), .B(n714), .C(\mem<191> ), .Y(n151) );
  OAI21X1 U187 ( .A(n130), .B(n716), .C(n153), .Y(n443) );
  OAI21X1 U188 ( .A(n43), .B(n714), .C(\mem<190> ), .Y(n153) );
  OAI21X1 U189 ( .A(n679), .B(n716), .C(n154), .Y(n444) );
  OAI21X1 U190 ( .A(n40), .B(n714), .C(\mem<189> ), .Y(n154) );
  OAI21X1 U191 ( .A(n678), .B(n716), .C(n155), .Y(n445) );
  OAI21X1 U192 ( .A(n38), .B(n714), .C(\mem<188> ), .Y(n155) );
  OAI21X1 U193 ( .A(n112), .B(n716), .C(n156), .Y(n446) );
  OAI21X1 U194 ( .A(n36), .B(n714), .C(\mem<187> ), .Y(n156) );
  OAI21X1 U195 ( .A(n93), .B(n716), .C(n157), .Y(n447) );
  OAI21X1 U196 ( .A(n34), .B(n714), .C(\mem<186> ), .Y(n157) );
  OAI21X1 U197 ( .A(n87), .B(n716), .C(n158), .Y(n448) );
  OAI21X1 U198 ( .A(n32), .B(n714), .C(\mem<185> ), .Y(n158) );
  OAI21X1 U199 ( .A(n84), .B(n716), .C(n159), .Y(n449) );
  OAI21X1 U200 ( .A(n30), .B(n714), .C(\mem<184> ), .Y(n159) );
  OAI21X1 U201 ( .A(n677), .B(n715), .C(n160), .Y(n450) );
  OAI21X1 U202 ( .A(n28), .B(n713), .C(\mem<183> ), .Y(n160) );
  OAI21X1 U203 ( .A(n676), .B(n715), .C(n161), .Y(n451) );
  OAI21X1 U204 ( .A(n26), .B(n713), .C(\mem<182> ), .Y(n161) );
  OAI21X1 U205 ( .A(n675), .B(n715), .C(n162), .Y(n452) );
  OAI21X1 U206 ( .A(n24), .B(n713), .C(\mem<181> ), .Y(n162) );
  OAI21X1 U207 ( .A(n674), .B(n715), .C(n163), .Y(n453) );
  OAI21X1 U208 ( .A(n22), .B(n713), .C(\mem<180> ), .Y(n163) );
  OAI21X1 U209 ( .A(n673), .B(n715), .C(n164), .Y(n454) );
  OAI21X1 U210 ( .A(n20), .B(n713), .C(\mem<179> ), .Y(n164) );
  OAI21X1 U211 ( .A(n672), .B(n715), .C(n165), .Y(n455) );
  OAI21X1 U212 ( .A(n18), .B(n713), .C(\mem<178> ), .Y(n165) );
  OAI21X1 U213 ( .A(n671), .B(n715), .C(n166), .Y(n456) );
  OAI21X1 U214 ( .A(n16), .B(n713), .C(\mem<177> ), .Y(n166) );
  OAI21X1 U215 ( .A(n665), .B(n715), .C(n167), .Y(n457) );
  OAI21X1 U216 ( .A(n14), .B(n713), .C(\mem<176> ), .Y(n167) );
  OAI21X1 U219 ( .A(n133), .B(n712), .C(n170), .Y(n458) );
  OAI21X1 U220 ( .A(n45), .B(n710), .C(\mem<175> ), .Y(n170) );
  OAI21X1 U221 ( .A(n130), .B(n712), .C(n172), .Y(n459) );
  OAI21X1 U222 ( .A(n43), .B(n710), .C(\mem<174> ), .Y(n172) );
  OAI21X1 U223 ( .A(n679), .B(n712), .C(n173), .Y(n460) );
  OAI21X1 U224 ( .A(n40), .B(n710), .C(\mem<173> ), .Y(n173) );
  OAI21X1 U225 ( .A(n678), .B(n712), .C(n174), .Y(n461) );
  OAI21X1 U226 ( .A(n38), .B(n710), .C(\mem<172> ), .Y(n174) );
  OAI21X1 U227 ( .A(n112), .B(n712), .C(n175), .Y(n462) );
  OAI21X1 U228 ( .A(n36), .B(n710), .C(\mem<171> ), .Y(n175) );
  OAI21X1 U229 ( .A(n93), .B(n712), .C(n176), .Y(n463) );
  OAI21X1 U230 ( .A(n34), .B(n710), .C(\mem<170> ), .Y(n176) );
  OAI21X1 U231 ( .A(n87), .B(n712), .C(n177), .Y(n464) );
  OAI21X1 U232 ( .A(n32), .B(n710), .C(\mem<169> ), .Y(n177) );
  OAI21X1 U233 ( .A(n84), .B(n712), .C(n178), .Y(n465) );
  OAI21X1 U234 ( .A(n30), .B(n710), .C(\mem<168> ), .Y(n178) );
  OAI21X1 U235 ( .A(n677), .B(n711), .C(n179), .Y(n466) );
  OAI21X1 U236 ( .A(n28), .B(n709), .C(\mem<167> ), .Y(n179) );
  OAI21X1 U237 ( .A(n676), .B(n711), .C(n180), .Y(n467) );
  OAI21X1 U238 ( .A(n26), .B(n709), .C(\mem<166> ), .Y(n180) );
  OAI21X1 U239 ( .A(n675), .B(n711), .C(n181), .Y(n468) );
  OAI21X1 U240 ( .A(n24), .B(n709), .C(\mem<165> ), .Y(n181) );
  OAI21X1 U241 ( .A(n674), .B(n711), .C(n182), .Y(n469) );
  OAI21X1 U242 ( .A(n22), .B(n709), .C(\mem<164> ), .Y(n182) );
  OAI21X1 U243 ( .A(n673), .B(n711), .C(n183), .Y(n470) );
  OAI21X1 U244 ( .A(n20), .B(n709), .C(\mem<163> ), .Y(n183) );
  OAI21X1 U245 ( .A(n672), .B(n711), .C(n184), .Y(n471) );
  OAI21X1 U246 ( .A(n18), .B(n709), .C(\mem<162> ), .Y(n184) );
  OAI21X1 U247 ( .A(n671), .B(n711), .C(n185), .Y(n472) );
  OAI21X1 U248 ( .A(n16), .B(n709), .C(\mem<161> ), .Y(n185) );
  OAI21X1 U249 ( .A(n665), .B(n711), .C(n186), .Y(n473) );
  OAI21X1 U250 ( .A(n14), .B(n709), .C(\mem<160> ), .Y(n186) );
  OAI21X1 U253 ( .A(n133), .B(n708), .C(n188), .Y(n474) );
  OAI21X1 U254 ( .A(n45), .B(n706), .C(\mem<159> ), .Y(n188) );
  OAI21X1 U255 ( .A(n130), .B(n708), .C(n190), .Y(n475) );
  OAI21X1 U256 ( .A(n43), .B(n706), .C(\mem<158> ), .Y(n190) );
  OAI21X1 U257 ( .A(n679), .B(n708), .C(n191), .Y(n476) );
  OAI21X1 U258 ( .A(n40), .B(n706), .C(\mem<157> ), .Y(n191) );
  OAI21X1 U259 ( .A(n678), .B(n708), .C(n192), .Y(n477) );
  OAI21X1 U260 ( .A(n38), .B(n706), .C(\mem<156> ), .Y(n192) );
  OAI21X1 U261 ( .A(n112), .B(n708), .C(n193), .Y(n478) );
  OAI21X1 U262 ( .A(n36), .B(n706), .C(\mem<155> ), .Y(n193) );
  OAI21X1 U263 ( .A(n93), .B(n708), .C(n194), .Y(n479) );
  OAI21X1 U264 ( .A(n34), .B(n706), .C(\mem<154> ), .Y(n194) );
  OAI21X1 U265 ( .A(n87), .B(n708), .C(n195), .Y(n480) );
  OAI21X1 U266 ( .A(n32), .B(n706), .C(\mem<153> ), .Y(n195) );
  OAI21X1 U267 ( .A(n84), .B(n708), .C(n196), .Y(n481) );
  OAI21X1 U268 ( .A(n30), .B(n706), .C(\mem<152> ), .Y(n196) );
  OAI21X1 U269 ( .A(n677), .B(n707), .C(n197), .Y(n482) );
  OAI21X1 U270 ( .A(n28), .B(n705), .C(\mem<151> ), .Y(n197) );
  OAI21X1 U271 ( .A(n676), .B(n707), .C(n198), .Y(n483) );
  OAI21X1 U272 ( .A(n26), .B(n705), .C(\mem<150> ), .Y(n198) );
  OAI21X1 U273 ( .A(n675), .B(n707), .C(n199), .Y(n484) );
  OAI21X1 U274 ( .A(n24), .B(n705), .C(\mem<149> ), .Y(n199) );
  OAI21X1 U275 ( .A(n674), .B(n707), .C(n200), .Y(n485) );
  OAI21X1 U276 ( .A(n22), .B(n705), .C(\mem<148> ), .Y(n200) );
  OAI21X1 U277 ( .A(n673), .B(n707), .C(n201), .Y(n486) );
  OAI21X1 U278 ( .A(n20), .B(n705), .C(\mem<147> ), .Y(n201) );
  OAI21X1 U279 ( .A(n672), .B(n707), .C(n202), .Y(n487) );
  OAI21X1 U280 ( .A(n18), .B(n705), .C(\mem<146> ), .Y(n202) );
  OAI21X1 U281 ( .A(n671), .B(n707), .C(n203), .Y(n488) );
  OAI21X1 U282 ( .A(n16), .B(n705), .C(\mem<145> ), .Y(n203) );
  OAI21X1 U283 ( .A(n665), .B(n707), .C(n204), .Y(n489) );
  OAI21X1 U284 ( .A(n14), .B(n705), .C(\mem<144> ), .Y(n204) );
  OAI21X1 U287 ( .A(n133), .B(n704), .C(n206), .Y(n490) );
  OAI21X1 U288 ( .A(n45), .B(n702), .C(\mem<143> ), .Y(n206) );
  OAI21X1 U289 ( .A(n130), .B(n704), .C(n208), .Y(n491) );
  OAI21X1 U290 ( .A(n43), .B(n702), .C(\mem<142> ), .Y(n208) );
  OAI21X1 U291 ( .A(n679), .B(n704), .C(n209), .Y(n492) );
  OAI21X1 U292 ( .A(n40), .B(n702), .C(\mem<141> ), .Y(n209) );
  OAI21X1 U293 ( .A(n678), .B(n704), .C(n210), .Y(n493) );
  OAI21X1 U294 ( .A(n38), .B(n702), .C(\mem<140> ), .Y(n210) );
  OAI21X1 U295 ( .A(n112), .B(n704), .C(n211), .Y(n494) );
  OAI21X1 U296 ( .A(n36), .B(n702), .C(\mem<139> ), .Y(n211) );
  OAI21X1 U297 ( .A(n93), .B(n704), .C(n212), .Y(n495) );
  OAI21X1 U298 ( .A(n34), .B(n702), .C(\mem<138> ), .Y(n212) );
  OAI21X1 U299 ( .A(n87), .B(n704), .C(n213), .Y(n496) );
  OAI21X1 U300 ( .A(n32), .B(n702), .C(\mem<137> ), .Y(n213) );
  OAI21X1 U301 ( .A(n84), .B(n704), .C(n214), .Y(n497) );
  OAI21X1 U302 ( .A(n30), .B(n702), .C(\mem<136> ), .Y(n214) );
  OAI21X1 U303 ( .A(n677), .B(n703), .C(n215), .Y(n498) );
  OAI21X1 U304 ( .A(n28), .B(n701), .C(\mem<135> ), .Y(n215) );
  OAI21X1 U305 ( .A(n676), .B(n703), .C(n216), .Y(n499) );
  OAI21X1 U306 ( .A(n26), .B(n701), .C(\mem<134> ), .Y(n216) );
  OAI21X1 U307 ( .A(n675), .B(n703), .C(n217), .Y(n500) );
  OAI21X1 U308 ( .A(n24), .B(n701), .C(\mem<133> ), .Y(n217) );
  OAI21X1 U309 ( .A(n674), .B(n703), .C(n218), .Y(n501) );
  OAI21X1 U310 ( .A(n22), .B(n701), .C(\mem<132> ), .Y(n218) );
  OAI21X1 U311 ( .A(n673), .B(n703), .C(n219), .Y(n502) );
  OAI21X1 U312 ( .A(n20), .B(n701), .C(\mem<131> ), .Y(n219) );
  OAI21X1 U313 ( .A(n672), .B(n703), .C(n220), .Y(n503) );
  OAI21X1 U314 ( .A(n18), .B(n701), .C(\mem<130> ), .Y(n220) );
  OAI21X1 U315 ( .A(n671), .B(n703), .C(n221), .Y(n504) );
  OAI21X1 U316 ( .A(n16), .B(n701), .C(\mem<129> ), .Y(n221) );
  OAI21X1 U317 ( .A(n665), .B(n703), .C(n222), .Y(n505) );
  OAI21X1 U318 ( .A(n14), .B(n701), .C(\mem<128> ), .Y(n222) );
  OAI21X1 U321 ( .A(n133), .B(n700), .C(n224), .Y(n506) );
  OAI21X1 U322 ( .A(n45), .B(n698), .C(\mem<127> ), .Y(n224) );
  OAI21X1 U323 ( .A(n130), .B(n700), .C(n226), .Y(n507) );
  OAI21X1 U324 ( .A(n43), .B(n698), .C(\mem<126> ), .Y(n226) );
  OAI21X1 U325 ( .A(n679), .B(n700), .C(n227), .Y(n508) );
  OAI21X1 U326 ( .A(n40), .B(n698), .C(\mem<125> ), .Y(n227) );
  OAI21X1 U327 ( .A(n678), .B(n700), .C(n228), .Y(n509) );
  OAI21X1 U328 ( .A(n38), .B(n698), .C(\mem<124> ), .Y(n228) );
  OAI21X1 U329 ( .A(n112), .B(n700), .C(n229), .Y(n510) );
  OAI21X1 U330 ( .A(n36), .B(n698), .C(\mem<123> ), .Y(n229) );
  OAI21X1 U331 ( .A(n93), .B(n700), .C(n230), .Y(n511) );
  OAI21X1 U332 ( .A(n34), .B(n698), .C(\mem<122> ), .Y(n230) );
  OAI21X1 U333 ( .A(n87), .B(n700), .C(n231), .Y(n512) );
  OAI21X1 U334 ( .A(n32), .B(n698), .C(\mem<121> ), .Y(n231) );
  OAI21X1 U335 ( .A(n84), .B(n700), .C(n232), .Y(n513) );
  OAI21X1 U336 ( .A(n30), .B(n698), .C(\mem<120> ), .Y(n232) );
  OAI21X1 U337 ( .A(n677), .B(n699), .C(n233), .Y(n514) );
  OAI21X1 U338 ( .A(n28), .B(n698), .C(\mem<119> ), .Y(n233) );
  OAI21X1 U339 ( .A(n676), .B(n699), .C(n234), .Y(n515) );
  OAI21X1 U340 ( .A(n26), .B(n698), .C(\mem<118> ), .Y(n234) );
  OAI21X1 U341 ( .A(n675), .B(n699), .C(n235), .Y(n516) );
  OAI21X1 U342 ( .A(n24), .B(n698), .C(\mem<117> ), .Y(n235) );
  OAI21X1 U343 ( .A(n674), .B(n699), .C(n236), .Y(n517) );
  OAI21X1 U344 ( .A(n22), .B(n698), .C(\mem<116> ), .Y(n236) );
  OAI21X1 U345 ( .A(n673), .B(n699), .C(n237), .Y(n518) );
  OAI21X1 U346 ( .A(n20), .B(n698), .C(\mem<115> ), .Y(n237) );
  OAI21X1 U347 ( .A(n672), .B(n699), .C(n238), .Y(n519) );
  OAI21X1 U348 ( .A(n18), .B(n698), .C(\mem<114> ), .Y(n238) );
  OAI21X1 U349 ( .A(n671), .B(n699), .C(n239), .Y(n520) );
  OAI21X1 U350 ( .A(n16), .B(n698), .C(\mem<113> ), .Y(n239) );
  OAI21X1 U351 ( .A(n665), .B(n699), .C(n240), .Y(n521) );
  OAI21X1 U352 ( .A(n14), .B(n698), .C(\mem<112> ), .Y(n240) );
  OAI21X1 U355 ( .A(n133), .B(n697), .C(n243), .Y(n522) );
  OAI21X1 U356 ( .A(n45), .B(n695), .C(\mem<111> ), .Y(n243) );
  OAI21X1 U357 ( .A(n130), .B(n697), .C(n245), .Y(n523) );
  OAI21X1 U358 ( .A(n43), .B(n695), .C(\mem<110> ), .Y(n245) );
  OAI21X1 U359 ( .A(n679), .B(n697), .C(n246), .Y(n524) );
  OAI21X1 U360 ( .A(n40), .B(n695), .C(\mem<109> ), .Y(n246) );
  OAI21X1 U361 ( .A(n678), .B(n697), .C(n247), .Y(n525) );
  OAI21X1 U362 ( .A(n38), .B(n695), .C(\mem<108> ), .Y(n247) );
  OAI21X1 U363 ( .A(n112), .B(n697), .C(n248), .Y(n526) );
  OAI21X1 U364 ( .A(n36), .B(n695), .C(\mem<107> ), .Y(n248) );
  OAI21X1 U365 ( .A(n93), .B(n697), .C(n249), .Y(n527) );
  OAI21X1 U366 ( .A(n34), .B(n695), .C(\mem<106> ), .Y(n249) );
  OAI21X1 U367 ( .A(n87), .B(n697), .C(n250), .Y(n528) );
  OAI21X1 U368 ( .A(n32), .B(n695), .C(\mem<105> ), .Y(n250) );
  OAI21X1 U369 ( .A(n84), .B(n697), .C(n251), .Y(n529) );
  OAI21X1 U370 ( .A(n30), .B(n695), .C(\mem<104> ), .Y(n251) );
  OAI21X1 U371 ( .A(n677), .B(n696), .C(n252), .Y(n530) );
  OAI21X1 U372 ( .A(n28), .B(n695), .C(\mem<103> ), .Y(n252) );
  OAI21X1 U373 ( .A(n676), .B(n696), .C(n253), .Y(n531) );
  OAI21X1 U374 ( .A(n26), .B(n695), .C(\mem<102> ), .Y(n253) );
  OAI21X1 U375 ( .A(n675), .B(n696), .C(n254), .Y(n532) );
  OAI21X1 U376 ( .A(n24), .B(n695), .C(\mem<101> ), .Y(n254) );
  OAI21X1 U377 ( .A(n674), .B(n696), .C(n255), .Y(n533) );
  OAI21X1 U378 ( .A(n22), .B(n695), .C(\mem<100> ), .Y(n255) );
  OAI21X1 U379 ( .A(n673), .B(n696), .C(n256), .Y(n534) );
  OAI21X1 U380 ( .A(n20), .B(n695), .C(\mem<99> ), .Y(n256) );
  OAI21X1 U381 ( .A(n672), .B(n696), .C(n257), .Y(n535) );
  OAI21X1 U382 ( .A(n18), .B(n695), .C(\mem<98> ), .Y(n257) );
  OAI21X1 U383 ( .A(n671), .B(n696), .C(n258), .Y(n536) );
  OAI21X1 U384 ( .A(n16), .B(n695), .C(\mem<97> ), .Y(n258) );
  OAI21X1 U385 ( .A(n665), .B(n696), .C(n259), .Y(n537) );
  OAI21X1 U386 ( .A(n14), .B(n695), .C(\mem<96> ), .Y(n259) );
  OAI21X1 U389 ( .A(n133), .B(n694), .C(n261), .Y(n538) );
  OAI21X1 U390 ( .A(n45), .B(n692), .C(\mem<95> ), .Y(n261) );
  OAI21X1 U391 ( .A(n130), .B(n694), .C(n263), .Y(n539) );
  OAI21X1 U392 ( .A(n43), .B(n692), .C(\mem<94> ), .Y(n263) );
  OAI21X1 U393 ( .A(n679), .B(n694), .C(n264), .Y(n540) );
  OAI21X1 U394 ( .A(n40), .B(n692), .C(\mem<93> ), .Y(n264) );
  OAI21X1 U395 ( .A(n678), .B(n694), .C(n265), .Y(n541) );
  OAI21X1 U396 ( .A(n38), .B(n692), .C(\mem<92> ), .Y(n265) );
  OAI21X1 U397 ( .A(n112), .B(n694), .C(n266), .Y(n542) );
  OAI21X1 U398 ( .A(n36), .B(n692), .C(\mem<91> ), .Y(n266) );
  OAI21X1 U399 ( .A(n93), .B(n694), .C(n267), .Y(n543) );
  OAI21X1 U400 ( .A(n34), .B(n692), .C(\mem<90> ), .Y(n267) );
  OAI21X1 U401 ( .A(n87), .B(n694), .C(n268), .Y(n544) );
  OAI21X1 U402 ( .A(n32), .B(n692), .C(\mem<89> ), .Y(n268) );
  OAI21X1 U403 ( .A(n84), .B(n694), .C(n269), .Y(n545) );
  OAI21X1 U404 ( .A(n30), .B(n692), .C(\mem<88> ), .Y(n269) );
  OAI21X1 U405 ( .A(n677), .B(n693), .C(n270), .Y(n546) );
  OAI21X1 U406 ( .A(n28), .B(n692), .C(\mem<87> ), .Y(n270) );
  OAI21X1 U407 ( .A(n676), .B(n693), .C(n271), .Y(n547) );
  OAI21X1 U408 ( .A(n26), .B(n692), .C(\mem<86> ), .Y(n271) );
  OAI21X1 U409 ( .A(n675), .B(n693), .C(n272), .Y(n548) );
  OAI21X1 U410 ( .A(n24), .B(n692), .C(\mem<85> ), .Y(n272) );
  OAI21X1 U411 ( .A(n674), .B(n693), .C(n273), .Y(n549) );
  OAI21X1 U412 ( .A(n22), .B(n692), .C(\mem<84> ), .Y(n273) );
  OAI21X1 U413 ( .A(n673), .B(n693), .C(n274), .Y(n550) );
  OAI21X1 U414 ( .A(n20), .B(n692), .C(\mem<83> ), .Y(n274) );
  OAI21X1 U415 ( .A(n672), .B(n693), .C(n275), .Y(n551) );
  OAI21X1 U416 ( .A(n18), .B(n692), .C(\mem<82> ), .Y(n275) );
  OAI21X1 U417 ( .A(n671), .B(n693), .C(n276), .Y(n552) );
  OAI21X1 U418 ( .A(n16), .B(n692), .C(\mem<81> ), .Y(n276) );
  OAI21X1 U419 ( .A(n665), .B(n693), .C(n277), .Y(n553) );
  OAI21X1 U420 ( .A(n14), .B(n692), .C(\mem<80> ), .Y(n277) );
  OAI21X1 U423 ( .A(n133), .B(n691), .C(n279), .Y(n554) );
  OAI21X1 U424 ( .A(n45), .B(n689), .C(\mem<79> ), .Y(n279) );
  OAI21X1 U425 ( .A(n130), .B(n691), .C(n281), .Y(n555) );
  OAI21X1 U426 ( .A(n43), .B(n689), .C(\mem<78> ), .Y(n281) );
  OAI21X1 U427 ( .A(n679), .B(n691), .C(n282), .Y(n556) );
  OAI21X1 U428 ( .A(n40), .B(n689), .C(\mem<77> ), .Y(n282) );
  OAI21X1 U429 ( .A(n678), .B(n691), .C(n283), .Y(n557) );
  OAI21X1 U430 ( .A(n38), .B(n689), .C(\mem<76> ), .Y(n283) );
  OAI21X1 U431 ( .A(n112), .B(n691), .C(n284), .Y(n558) );
  OAI21X1 U432 ( .A(n36), .B(n689), .C(\mem<75> ), .Y(n284) );
  OAI21X1 U433 ( .A(n93), .B(n691), .C(n285), .Y(n559) );
  OAI21X1 U434 ( .A(n34), .B(n689), .C(\mem<74> ), .Y(n285) );
  OAI21X1 U435 ( .A(n87), .B(n691), .C(n286), .Y(n560) );
  OAI21X1 U436 ( .A(n32), .B(n689), .C(\mem<73> ), .Y(n286) );
  OAI21X1 U437 ( .A(n84), .B(n691), .C(n287), .Y(n561) );
  OAI21X1 U438 ( .A(n30), .B(n689), .C(\mem<72> ), .Y(n287) );
  OAI21X1 U439 ( .A(n677), .B(n690), .C(n288), .Y(n562) );
  OAI21X1 U440 ( .A(n28), .B(n689), .C(\mem<71> ), .Y(n288) );
  OAI21X1 U441 ( .A(n676), .B(n690), .C(n289), .Y(n563) );
  OAI21X1 U442 ( .A(n26), .B(n689), .C(\mem<70> ), .Y(n289) );
  OAI21X1 U443 ( .A(n675), .B(n690), .C(n290), .Y(n564) );
  OAI21X1 U444 ( .A(n24), .B(n689), .C(\mem<69> ), .Y(n290) );
  OAI21X1 U445 ( .A(n674), .B(n690), .C(n291), .Y(n565) );
  OAI21X1 U446 ( .A(n22), .B(n689), .C(\mem<68> ), .Y(n291) );
  OAI21X1 U447 ( .A(n673), .B(n690), .C(n292), .Y(n566) );
  OAI21X1 U448 ( .A(n20), .B(n689), .C(\mem<67> ), .Y(n292) );
  OAI21X1 U449 ( .A(n672), .B(n690), .C(n293), .Y(n567) );
  OAI21X1 U450 ( .A(n18), .B(n689), .C(\mem<66> ), .Y(n293) );
  OAI21X1 U451 ( .A(n671), .B(n690), .C(n294), .Y(n568) );
  OAI21X1 U452 ( .A(n16), .B(n689), .C(\mem<65> ), .Y(n294) );
  OAI21X1 U453 ( .A(n665), .B(n690), .C(n295), .Y(n569) );
  OAI21X1 U454 ( .A(n14), .B(n689), .C(\mem<64> ), .Y(n295) );
  OAI21X1 U458 ( .A(n133), .B(n688), .C(n297), .Y(n570) );
  OAI21X1 U459 ( .A(n45), .B(n686), .C(\mem<63> ), .Y(n297) );
  OAI21X1 U460 ( .A(n130), .B(n688), .C(n299), .Y(n571) );
  OAI21X1 U461 ( .A(n43), .B(n686), .C(\mem<62> ), .Y(n299) );
  OAI21X1 U462 ( .A(n679), .B(n688), .C(n300), .Y(n572) );
  OAI21X1 U463 ( .A(n40), .B(n686), .C(\mem<61> ), .Y(n300) );
  OAI21X1 U464 ( .A(n678), .B(n688), .C(n301), .Y(n573) );
  OAI21X1 U465 ( .A(n38), .B(n686), .C(\mem<60> ), .Y(n301) );
  OAI21X1 U466 ( .A(n112), .B(n688), .C(n302), .Y(n574) );
  OAI21X1 U467 ( .A(n36), .B(n686), .C(\mem<59> ), .Y(n302) );
  OAI21X1 U468 ( .A(n93), .B(n688), .C(n303), .Y(n575) );
  OAI21X1 U469 ( .A(n34), .B(n686), .C(\mem<58> ), .Y(n303) );
  OAI21X1 U470 ( .A(n87), .B(n688), .C(n304), .Y(n576) );
  OAI21X1 U471 ( .A(n32), .B(n686), .C(\mem<57> ), .Y(n304) );
  OAI21X1 U472 ( .A(n84), .B(n688), .C(n305), .Y(n577) );
  OAI21X1 U473 ( .A(n30), .B(n686), .C(\mem<56> ), .Y(n305) );
  OAI21X1 U474 ( .A(n677), .B(n687), .C(n306), .Y(n578) );
  OAI21X1 U475 ( .A(n28), .B(n686), .C(\mem<55> ), .Y(n306) );
  OAI21X1 U476 ( .A(n676), .B(n687), .C(n307), .Y(n579) );
  OAI21X1 U477 ( .A(n26), .B(n686), .C(\mem<54> ), .Y(n307) );
  OAI21X1 U478 ( .A(n675), .B(n687), .C(n308), .Y(n580) );
  OAI21X1 U479 ( .A(n24), .B(n686), .C(\mem<53> ), .Y(n308) );
  OAI21X1 U480 ( .A(n674), .B(n687), .C(n309), .Y(n581) );
  OAI21X1 U481 ( .A(n22), .B(n686), .C(\mem<52> ), .Y(n309) );
  OAI21X1 U482 ( .A(n673), .B(n687), .C(n310), .Y(n582) );
  OAI21X1 U483 ( .A(n20), .B(n686), .C(\mem<51> ), .Y(n310) );
  OAI21X1 U484 ( .A(n672), .B(n687), .C(n311), .Y(n583) );
  OAI21X1 U485 ( .A(n18), .B(n686), .C(\mem<50> ), .Y(n311) );
  OAI21X1 U486 ( .A(n671), .B(n687), .C(n312), .Y(n584) );
  OAI21X1 U487 ( .A(n16), .B(n686), .C(\mem<49> ), .Y(n312) );
  OAI21X1 U488 ( .A(n665), .B(n687), .C(n313), .Y(n585) );
  OAI21X1 U489 ( .A(n14), .B(n686), .C(\mem<48> ), .Y(n313) );
  OAI21X1 U492 ( .A(n133), .B(n685), .C(n316), .Y(n586) );
  OAI21X1 U493 ( .A(n45), .B(n683), .C(\mem<47> ), .Y(n316) );
  OAI21X1 U494 ( .A(n130), .B(n685), .C(n318), .Y(n587) );
  OAI21X1 U495 ( .A(n43), .B(n683), .C(\mem<46> ), .Y(n318) );
  OAI21X1 U496 ( .A(n679), .B(n685), .C(n319), .Y(n588) );
  OAI21X1 U497 ( .A(n40), .B(n683), .C(\mem<45> ), .Y(n319) );
  OAI21X1 U498 ( .A(n678), .B(n685), .C(n320), .Y(n589) );
  OAI21X1 U499 ( .A(n38), .B(n683), .C(\mem<44> ), .Y(n320) );
  OAI21X1 U500 ( .A(n112), .B(n685), .C(n321), .Y(n590) );
  OAI21X1 U501 ( .A(n36), .B(n683), .C(\mem<43> ), .Y(n321) );
  OAI21X1 U502 ( .A(n93), .B(n685), .C(n322), .Y(n591) );
  OAI21X1 U503 ( .A(n34), .B(n683), .C(\mem<42> ), .Y(n322) );
  OAI21X1 U504 ( .A(n87), .B(n685), .C(n323), .Y(n592) );
  OAI21X1 U505 ( .A(n32), .B(n683), .C(\mem<41> ), .Y(n323) );
  OAI21X1 U506 ( .A(n84), .B(n685), .C(n324), .Y(n593) );
  OAI21X1 U507 ( .A(n30), .B(n683), .C(\mem<40> ), .Y(n324) );
  OAI21X1 U508 ( .A(n677), .B(n684), .C(n325), .Y(n594) );
  OAI21X1 U509 ( .A(n28), .B(n683), .C(\mem<39> ), .Y(n325) );
  OAI21X1 U510 ( .A(n676), .B(n684), .C(n326), .Y(n595) );
  OAI21X1 U511 ( .A(n26), .B(n683), .C(\mem<38> ), .Y(n326) );
  OAI21X1 U512 ( .A(n675), .B(n684), .C(n327), .Y(n596) );
  OAI21X1 U513 ( .A(n24), .B(n683), .C(\mem<37> ), .Y(n327) );
  OAI21X1 U514 ( .A(n674), .B(n684), .C(n328), .Y(n597) );
  OAI21X1 U515 ( .A(n22), .B(n683), .C(\mem<36> ), .Y(n328) );
  OAI21X1 U516 ( .A(n673), .B(n684), .C(n329), .Y(n598) );
  OAI21X1 U517 ( .A(n20), .B(n683), .C(\mem<35> ), .Y(n329) );
  OAI21X1 U518 ( .A(n672), .B(n684), .C(n330), .Y(n599) );
  OAI21X1 U519 ( .A(n18), .B(n683), .C(\mem<34> ), .Y(n330) );
  OAI21X1 U520 ( .A(n671), .B(n684), .C(n331), .Y(n600) );
  OAI21X1 U521 ( .A(n16), .B(n683), .C(\mem<33> ), .Y(n331) );
  OAI21X1 U522 ( .A(n665), .B(n684), .C(n332), .Y(n601) );
  OAI21X1 U523 ( .A(n14), .B(n683), .C(\mem<32> ), .Y(n332) );
  OAI21X1 U526 ( .A(n133), .B(n682), .C(n334), .Y(n602) );
  OAI21X1 U527 ( .A(n45), .B(n680), .C(\mem<31> ), .Y(n334) );
  OAI21X1 U528 ( .A(n130), .B(n682), .C(n336), .Y(n603) );
  OAI21X1 U529 ( .A(n43), .B(n680), .C(\mem<30> ), .Y(n336) );
  OAI21X1 U530 ( .A(n679), .B(n682), .C(n337), .Y(n604) );
  OAI21X1 U531 ( .A(n40), .B(n680), .C(\mem<29> ), .Y(n337) );
  OAI21X1 U532 ( .A(n678), .B(n682), .C(n338), .Y(n605) );
  OAI21X1 U533 ( .A(n38), .B(n680), .C(\mem<28> ), .Y(n338) );
  OAI21X1 U534 ( .A(n112), .B(n682), .C(n339), .Y(n606) );
  OAI21X1 U535 ( .A(n36), .B(n680), .C(\mem<27> ), .Y(n339) );
  OAI21X1 U536 ( .A(n93), .B(n682), .C(n340), .Y(n607) );
  OAI21X1 U537 ( .A(n34), .B(n680), .C(\mem<26> ), .Y(n340) );
  OAI21X1 U538 ( .A(n87), .B(n682), .C(n341), .Y(n608) );
  OAI21X1 U539 ( .A(n32), .B(n680), .C(\mem<25> ), .Y(n341) );
  OAI21X1 U540 ( .A(n84), .B(n682), .C(n342), .Y(n609) );
  OAI21X1 U541 ( .A(n30), .B(n680), .C(\mem<24> ), .Y(n342) );
  OAI21X1 U542 ( .A(n677), .B(n681), .C(n343), .Y(n610) );
  OAI21X1 U543 ( .A(n28), .B(n680), .C(\mem<23> ), .Y(n343) );
  OAI21X1 U544 ( .A(n676), .B(n681), .C(n344), .Y(n611) );
  OAI21X1 U545 ( .A(n26), .B(n680), .C(\mem<22> ), .Y(n344) );
  OAI21X1 U546 ( .A(n675), .B(n681), .C(n345), .Y(n612) );
  OAI21X1 U547 ( .A(n24), .B(n680), .C(\mem<21> ), .Y(n345) );
  OAI21X1 U548 ( .A(n674), .B(n681), .C(n346), .Y(n613) );
  OAI21X1 U549 ( .A(n22), .B(n680), .C(\mem<20> ), .Y(n346) );
  OAI21X1 U550 ( .A(n673), .B(n681), .C(n347), .Y(n614) );
  OAI21X1 U551 ( .A(n20), .B(n680), .C(\mem<19> ), .Y(n347) );
  OAI21X1 U552 ( .A(n672), .B(n681), .C(n348), .Y(n615) );
  OAI21X1 U553 ( .A(n18), .B(n680), .C(\mem<18> ), .Y(n348) );
  OAI21X1 U554 ( .A(n671), .B(n681), .C(n349), .Y(n616) );
  OAI21X1 U555 ( .A(n16), .B(n680), .C(\mem<17> ), .Y(n349) );
  OAI21X1 U556 ( .A(n665), .B(n681), .C(n350), .Y(n617) );
  OAI21X1 U557 ( .A(n14), .B(n680), .C(\mem<16> ), .Y(n350) );
  OAI21X1 U561 ( .A(n133), .B(n670), .C(n352), .Y(n618) );
  OAI21X1 U562 ( .A(n45), .B(n666), .C(\mem<15> ), .Y(n352) );
  OAI21X1 U565 ( .A(n130), .B(n670), .C(n357), .Y(n619) );
  OAI21X1 U566 ( .A(n43), .B(n666), .C(\mem<14> ), .Y(n357) );
  OAI21X1 U569 ( .A(n679), .B(n670), .C(n359), .Y(n620) );
  OAI21X1 U570 ( .A(n40), .B(n666), .C(\mem<13> ), .Y(n359) );
  OAI21X1 U573 ( .A(n678), .B(n670), .C(n361), .Y(n621) );
  OAI21X1 U574 ( .A(n38), .B(n666), .C(\mem<12> ), .Y(n361) );
  OAI21X1 U577 ( .A(n112), .B(n670), .C(n363), .Y(n622) );
  OAI21X1 U578 ( .A(n36), .B(n666), .C(\mem<11> ), .Y(n363) );
  OAI21X1 U581 ( .A(n93), .B(n670), .C(n365), .Y(n623) );
  OAI21X1 U582 ( .A(n34), .B(n666), .C(\mem<10> ), .Y(n365) );
  OAI21X1 U585 ( .A(n87), .B(n670), .C(n366), .Y(n624) );
  OAI21X1 U586 ( .A(n32), .B(n666), .C(\mem<9> ), .Y(n366) );
  OAI21X1 U589 ( .A(n84), .B(n670), .C(n367), .Y(n625) );
  OAI21X1 U590 ( .A(n30), .B(n666), .C(\mem<8> ), .Y(n367) );
  OAI21X1 U593 ( .A(n677), .B(n669), .C(n368), .Y(n626) );
  OAI21X1 U594 ( .A(n28), .B(n666), .C(\mem<7> ), .Y(n368) );
  OAI21X1 U597 ( .A(n676), .B(n669), .C(n370), .Y(n627) );
  OAI21X1 U598 ( .A(n26), .B(n666), .C(\mem<6> ), .Y(n370) );
  OAI21X1 U601 ( .A(n675), .B(n669), .C(n371), .Y(n628) );
  OAI21X1 U602 ( .A(n24), .B(n666), .C(\mem<5> ), .Y(n371) );
  OAI21X1 U605 ( .A(n674), .B(n669), .C(n372), .Y(n629) );
  OAI21X1 U606 ( .A(n22), .B(n666), .C(\mem<4> ), .Y(n372) );
  OAI21X1 U610 ( .A(n673), .B(n669), .C(n373), .Y(n630) );
  OAI21X1 U611 ( .A(n20), .B(n666), .C(\mem<3> ), .Y(n373) );
  OAI21X1 U614 ( .A(n672), .B(n669), .C(n375), .Y(n631) );
  OAI21X1 U615 ( .A(n18), .B(n666), .C(\mem<2> ), .Y(n375) );
  OAI21X1 U618 ( .A(n671), .B(n669), .C(n376), .Y(n632) );
  OAI21X1 U619 ( .A(n16), .B(n666), .C(\mem<1> ), .Y(n376) );
  OAI21X1 U623 ( .A(n665), .B(n669), .C(n377), .Y(n633) );
  OAI21X1 U624 ( .A(n14), .B(n666), .C(\mem<0> ), .Y(n377) );
  AND2X1 U2 ( .A(n830), .B(n750), .Y(n3) );
  INVX1 U3 ( .A(N21), .Y(n762) );
  INVX2 U4 ( .A(N20), .Y(n760) );
  AND2X1 U5 ( .A(n831), .B(n660), .Y(n1) );
  INVX1 U10 ( .A(n750), .Y(n663) );
  AND2X1 U11 ( .A(n854), .B(n664), .Y(n11) );
  INVX2 U12 ( .A(N20), .Y(n759) );
  INVX1 U13 ( .A(N23), .Y(n662) );
  AND2X1 U14 ( .A(N25), .B(n765), .Y(n168) );
  AND2X1 U15 ( .A(data_in), .B(n668), .Y(n90) );
  AND2X1 U16 ( .A(N25), .B(N24), .Y(n91) );
  BUFX2 U17 ( .A(n90), .Y(n732) );
  AND2X1 U18 ( .A(N23), .B(n763), .Y(n92) );
  AND2X1 U19 ( .A(N23), .B(n764), .Y(n111) );
  INVX1 U20 ( .A(write), .Y(n1019) );
  BUFX2 U21 ( .A(n90), .Y(n731) );
  BUFX2 U22 ( .A(n78), .Y(n668) );
  BUFX2 U23 ( .A(n78), .Y(n667) );
  BUFX2 U24 ( .A(n643), .Y(n730) );
  BUFX2 U25 ( .A(n641), .Y(n727) );
  BUFX2 U26 ( .A(n643), .Y(n729) );
  BUFX2 U27 ( .A(n639), .Y(n726) );
  BUFX2 U28 ( .A(n637), .Y(n723) );
  BUFX2 U29 ( .A(n639), .Y(n725) );
  BUFX2 U30 ( .A(n635), .Y(n722) );
  BUFX2 U31 ( .A(n635), .Y(n721) );
  BUFX2 U32 ( .A(n374), .Y(n719) );
  BUFX2 U33 ( .A(n374), .Y(n718) );
  BUFX2 U34 ( .A(n362), .Y(n716) );
  BUFX2 U35 ( .A(n354), .Y(n713) );
  BUFX2 U36 ( .A(n362), .Y(n715) );
  BUFX2 U37 ( .A(n351), .Y(n712) );
  BUFX2 U38 ( .A(n333), .Y(n709) );
  BUFX2 U39 ( .A(n351), .Y(n711) );
  BUFX2 U40 ( .A(n315), .Y(n708) );
  BUFX2 U41 ( .A(n298), .Y(n705) );
  BUFX2 U42 ( .A(n315), .Y(n707) );
  BUFX2 U43 ( .A(n280), .Y(n704) );
  BUFX2 U44 ( .A(n262), .Y(n701) );
  BUFX2 U45 ( .A(n280), .Y(n703) );
  BUFX2 U46 ( .A(n244), .Y(n700) );
  BUFX2 U47 ( .A(n244), .Y(n699) );
  BUFX2 U48 ( .A(n241), .Y(n697) );
  BUFX2 U81 ( .A(n241), .Y(n696) );
  BUFX2 U82 ( .A(n223), .Y(n694) );
  BUFX2 U115 ( .A(n223), .Y(n693) );
  BUFX2 U116 ( .A(n205), .Y(n691) );
  BUFX2 U149 ( .A(n205), .Y(n690) );
  BUFX2 U150 ( .A(n187), .Y(n688) );
  BUFX2 U183 ( .A(n187), .Y(n687) );
  BUFX2 U184 ( .A(n169), .Y(n685) );
  BUFX2 U217 ( .A(n169), .Y(n684) );
  BUFX2 U218 ( .A(n150), .Y(n682) );
  BUFX2 U251 ( .A(n150), .Y(n681) );
  BUFX2 U252 ( .A(n81), .Y(n670) );
  BUFX2 U285 ( .A(n81), .Y(n669) );
  INVX1 U286 ( .A(n753), .Y(n752) );
  INVX1 U319 ( .A(n48), .Y(n666) );
  INVX1 U320 ( .A(n63), .Y(n680) );
  INVX1 U353 ( .A(n68), .Y(n689) );
  INVX1 U354 ( .A(n69), .Y(n692) );
  INVX1 U387 ( .A(n74), .Y(n717) );
  INVX1 U388 ( .A(n75), .Y(n720) );
  INVX1 U421 ( .A(n65), .Y(n683) );
  INVX1 U422 ( .A(n71), .Y(n695) );
  INVX1 U455 ( .A(n51), .Y(n672) );
  INVX1 U456 ( .A(n57), .Y(n676) );
  INVX1 U457 ( .A(n66), .Y(n686) );
  INVX1 U490 ( .A(n72), .Y(n698) );
  INVX1 U491 ( .A(n53), .Y(n673) );
  INVX1 U524 ( .A(n59), .Y(n677) );
  INVX1 U525 ( .A(N24), .Y(n765) );
  BUFX2 U558 ( .A(n262), .Y(n702) );
  BUFX2 U559 ( .A(n298), .Y(n706) );
  BUFX2 U560 ( .A(n333), .Y(n710) );
  BUFX2 U563 ( .A(n354), .Y(n714) );
  BUFX2 U564 ( .A(n637), .Y(n724) );
  BUFX2 U567 ( .A(n641), .Y(n728) );
  INVX1 U568 ( .A(n47), .Y(n665) );
  INVX1 U571 ( .A(n50), .Y(n671) );
  INVX1 U572 ( .A(n54), .Y(n674) );
  INVX1 U575 ( .A(n56), .Y(n675) );
  INVX1 U576 ( .A(n60), .Y(n678) );
  INVX1 U579 ( .A(n62), .Y(n679) );
  INVX1 U580 ( .A(n1), .Y(n2) );
  INVX1 U583 ( .A(n3), .Y(n4) );
  AND2X2 U584 ( .A(n2), .B(n4), .Y(n5) );
  AND2X2 U587 ( .A(n12), .B(n8), .Y(n6) );
  AND2X1 U588 ( .A(n853), .B(N21), .Y(n7) );
  INVX1 U591 ( .A(n7), .Y(n8) );
  OR2X1 U592 ( .A(rst), .B(write), .Y(n9) );
  INVX1 U595 ( .A(n9), .Y(n10) );
  INVX1 U596 ( .A(n11), .Y(n12) );
  AND2X1 U599 ( .A(n47), .B(n667), .Y(n13) );
  INVX1 U600 ( .A(n13), .Y(n14) );
  AND2X1 U603 ( .A(n50), .B(n667), .Y(n15) );
  INVX1 U604 ( .A(n15), .Y(n16) );
  AND2X1 U607 ( .A(n51), .B(n667), .Y(n17) );
  INVX1 U608 ( .A(n17), .Y(n18) );
  AND2X1 U609 ( .A(n53), .B(n667), .Y(n19) );
  INVX1 U612 ( .A(n19), .Y(n20) );
  AND2X1 U613 ( .A(n54), .B(n667), .Y(n21) );
  INVX1 U616 ( .A(n21), .Y(n22) );
  AND2X1 U617 ( .A(n56), .B(n667), .Y(n23) );
  INVX1 U620 ( .A(n23), .Y(n24) );
  AND2X1 U621 ( .A(n57), .B(n667), .Y(n25) );
  INVX1 U622 ( .A(n25), .Y(n26) );
  AND2X1 U625 ( .A(n59), .B(n667), .Y(n27) );
  INVX1 U626 ( .A(n27), .Y(n28) );
  AND2X1 U627 ( .A(n83), .B(n668), .Y(n29) );
  INVX1 U628 ( .A(n29), .Y(n30) );
  AND2X1 U629 ( .A(n86), .B(n668), .Y(n31) );
  INVX1 U630 ( .A(n31), .Y(n32) );
  AND2X1 U631 ( .A(n89), .B(n668), .Y(n33) );
  INVX1 U632 ( .A(n33), .Y(n34) );
  AND2X1 U633 ( .A(n95), .B(n668), .Y(n35) );
  INVX1 U634 ( .A(n35), .Y(n36) );
  AND2X1 U635 ( .A(n60), .B(n668), .Y(n37) );
  INVX1 U636 ( .A(n37), .Y(n38) );
  AND2X1 U637 ( .A(n62), .B(n668), .Y(n39) );
  INVX1 U638 ( .A(n39), .Y(n40) );
  AND2X1 U639 ( .A(n114), .B(n668), .Y(n41) );
  INVX1 U640 ( .A(n41), .Y(n43) );
  AND2X1 U641 ( .A(n131), .B(n668), .Y(n44) );
  INVX1 U642 ( .A(n44), .Y(n45) );
  AND2X1 U643 ( .A(n653), .B(n645), .Y(n47) );
  AND2X1 U644 ( .A(n655), .B(n647), .Y(n48) );
  AND2X1 U645 ( .A(n653), .B(n649), .Y(n50) );
  AND2X1 U646 ( .A(n653), .B(n358), .Y(n51) );
  AND2X1 U647 ( .A(n653), .B(n356), .Y(n53) );
  AND2X1 U648 ( .A(n657), .B(n645), .Y(n54) );
  AND2X1 U649 ( .A(n657), .B(n649), .Y(n56) );
  AND2X1 U650 ( .A(n657), .B(n358), .Y(n57) );
  AND2X1 U651 ( .A(n657), .B(n356), .Y(n59) );
  AND2X1 U652 ( .A(n645), .B(n355), .Y(n60) );
  AND2X1 U653 ( .A(n649), .B(n355), .Y(n62) );
  AND2X1 U654 ( .A(n655), .B(n651), .Y(n63) );
  AND2X1 U655 ( .A(n655), .B(n111), .Y(n65) );
  AND2X1 U656 ( .A(n655), .B(n92), .Y(n66) );
  AND2X1 U657 ( .A(n659), .B(n647), .Y(n68) );
  AND2X1 U658 ( .A(n659), .B(n651), .Y(n69) );
  AND2X1 U659 ( .A(n659), .B(n111), .Y(n71) );
  AND2X1 U660 ( .A(n659), .B(n92), .Y(n72) );
  AND2X1 U661 ( .A(n647), .B(n91), .Y(n74) );
  AND2X1 U662 ( .A(n651), .B(n91), .Y(n75) );
  OR2X1 U663 ( .A(n1019), .B(rst), .Y(n77) );
  INVX1 U664 ( .A(n77), .Y(n78) );
  AND2X1 U665 ( .A(n48), .B(n731), .Y(n80) );
  INVX1 U666 ( .A(n80), .Y(n81) );
  AND2X1 U667 ( .A(n364), .B(n645), .Y(n83) );
  INVX1 U668 ( .A(n83), .Y(n84) );
  AND2X1 U669 ( .A(n364), .B(n649), .Y(n86) );
  INVX1 U670 ( .A(n86), .Y(n87) );
  AND2X1 U671 ( .A(n364), .B(n358), .Y(n89) );
  INVX1 U672 ( .A(n89), .Y(n93) );
  AND2X1 U673 ( .A(n364), .B(n356), .Y(n95) );
  INVX1 U674 ( .A(n95), .Y(n112) );
  AND2X1 U675 ( .A(n358), .B(n355), .Y(n114) );
  INVX1 U676 ( .A(n114), .Y(n130) );
  AND2X1 U677 ( .A(n355), .B(n356), .Y(n131) );
  INVX1 U678 ( .A(n131), .Y(n133) );
  AND2X1 U679 ( .A(n63), .B(n731), .Y(n149) );
  INVX1 U680 ( .A(n149), .Y(n150) );
  AND2X1 U681 ( .A(n65), .B(n731), .Y(n152) );
  INVX1 U682 ( .A(n152), .Y(n169) );
  AND2X1 U683 ( .A(n66), .B(n731), .Y(n171) );
  INVX1 U684 ( .A(n171), .Y(n187) );
  AND2X1 U685 ( .A(n68), .B(n731), .Y(n189) );
  INVX1 U686 ( .A(n189), .Y(n205) );
  AND2X1 U687 ( .A(n69), .B(n731), .Y(n207) );
  INVX1 U688 ( .A(n207), .Y(n223) );
  AND2X1 U689 ( .A(n71), .B(n731), .Y(n225) );
  INVX1 U690 ( .A(n225), .Y(n241) );
  AND2X1 U691 ( .A(n72), .B(n732), .Y(n242) );
  INVX1 U692 ( .A(n242), .Y(n244) );
  AND2X1 U693 ( .A(n168), .B(n647), .Y(n260) );
  INVX1 U694 ( .A(n260), .Y(n262) );
  AND2X1 U695 ( .A(n260), .B(n732), .Y(n278) );
  INVX1 U696 ( .A(n278), .Y(n280) );
  AND2X1 U697 ( .A(n168), .B(n651), .Y(n296) );
  INVX1 U698 ( .A(n296), .Y(n298) );
  AND2X1 U699 ( .A(n296), .B(n732), .Y(n314) );
  INVX1 U700 ( .A(n314), .Y(n315) );
  AND2X1 U701 ( .A(n168), .B(n111), .Y(n317) );
  INVX1 U702 ( .A(n317), .Y(n333) );
  AND2X1 U703 ( .A(n317), .B(n732), .Y(n335) );
  INVX1 U704 ( .A(n335), .Y(n351) );
  AND2X1 U705 ( .A(n168), .B(n92), .Y(n353) );
  INVX1 U706 ( .A(n353), .Y(n354) );
  AND2X1 U707 ( .A(n353), .B(n732), .Y(n360) );
  INVX1 U708 ( .A(n360), .Y(n362) );
  AND2X1 U709 ( .A(n74), .B(n732), .Y(n369) );
  INVX1 U710 ( .A(n369), .Y(n374) );
  AND2X1 U711 ( .A(n75), .B(n732), .Y(n634) );
  INVX1 U712 ( .A(n634), .Y(n635) );
  AND2X1 U713 ( .A(n111), .B(n91), .Y(n636) );
  INVX1 U714 ( .A(n636), .Y(n637) );
  AND2X1 U715 ( .A(n636), .B(n732), .Y(n638) );
  INVX1 U716 ( .A(n638), .Y(n639) );
  AND2X1 U717 ( .A(n91), .B(n92), .Y(n640) );
  INVX1 U718 ( .A(n640), .Y(n641) );
  AND2X1 U719 ( .A(n731), .B(n640), .Y(n642) );
  INVX1 U720 ( .A(n642), .Y(n643) );
  OR2X1 U721 ( .A(n744), .B(n752), .Y(n644) );
  INVX1 U722 ( .A(n644), .Y(n645) );
  OR2X1 U723 ( .A(n763), .B(N23), .Y(n646) );
  INVX1 U724 ( .A(n646), .Y(n647) );
  OR2X1 U725 ( .A(n745), .B(n752), .Y(n648) );
  INVX1 U726 ( .A(n648), .Y(n649) );
  OR2X1 U727 ( .A(n764), .B(N23), .Y(n650) );
  INVX1 U728 ( .A(n650), .Y(n651) );
  OR2X1 U729 ( .A(n757), .B(N21), .Y(n652) );
  INVX1 U730 ( .A(n652), .Y(n653) );
  OR2X1 U731 ( .A(N24), .B(N25), .Y(n654) );
  INVX1 U732 ( .A(n654), .Y(n655) );
  OR2X1 U733 ( .A(n758), .B(N21), .Y(n656) );
  INVX1 U734 ( .A(n656), .Y(n657) );
  OR2X1 U735 ( .A(n765), .B(N25), .Y(n658) );
  INVX1 U736 ( .A(n658), .Y(n659) );
  INVX8 U737 ( .A(n747), .Y(n742) );
  INVX1 U738 ( .A(n749), .Y(n660) );
  MUX2X1 U739 ( .B(n851), .A(n852), .S(n760), .Y(n853) );
  INVX2 U740 ( .A(n760), .Y(n756) );
  MUX2X1 U741 ( .B(\mem<85> ), .A(\mem<84> ), .S(n747), .Y(n844) );
  INVX1 U742 ( .A(N18), .Y(n661) );
  INVX4 U743 ( .A(n734), .Y(n748) );
  INVX2 U744 ( .A(N19), .Y(n753) );
  INVX4 U745 ( .A(N19), .Y(n754) );
  INVX1 U746 ( .A(N18), .Y(n735) );
  INVX4 U747 ( .A(n661), .Y(n733) );
  INVX1 U748 ( .A(n735), .Y(n734) );
  MUX2X1 U749 ( .B(n884), .A(n885), .S(n764), .Y(n886) );
  MUX2X1 U750 ( .B(n826), .A(n827), .S(n662), .Y(n889) );
  MUX2X1 U751 ( .B(n5), .A(n832), .S(n759), .Y(n840) );
  INVX2 U752 ( .A(n759), .Y(n757) );
  MUX2X1 U753 ( .B(\mem<87> ), .A(\mem<86> ), .S(n747), .Y(n843) );
  MUX2X1 U754 ( .B(\mem<81> ), .A(\mem<80> ), .S(n747), .Y(n842) );
  MUX2X1 U755 ( .B(n770), .A(n771), .S(n758), .Y(n779) );
  INVX2 U756 ( .A(n758), .Y(n755) );
  MUX2X1 U757 ( .B(n766), .A(n767), .S(n663), .Y(n771) );
  MUX2X1 U758 ( .B(\mem<83> ), .A(\mem<82> ), .S(n747), .Y(n841) );
  INVX1 U759 ( .A(N21), .Y(n664) );
  INVX2 U760 ( .A(n762), .Y(n761) );
  MUX2X1 U761 ( .B(n855), .A(n6), .S(N22), .Y(n887) );
  INVX1 U762 ( .A(N22), .Y(n764) );
  MUX2X1 U763 ( .B(n888), .A(n889), .S(n765), .Y(n1017) );
  INVX1 U764 ( .A(n764), .Y(n763) );
  INVX8 U765 ( .A(n745), .Y(n736) );
  INVX8 U766 ( .A(n745), .Y(n737) );
  INVX8 U767 ( .A(n746), .Y(n738) );
  INVX8 U768 ( .A(n746), .Y(n739) );
  INVX8 U769 ( .A(n747), .Y(n740) );
  INVX8 U770 ( .A(n747), .Y(n741) );
  INVX8 U771 ( .A(n748), .Y(n743) );
  INVX8 U772 ( .A(n748), .Y(n744) );
  INVX8 U773 ( .A(n733), .Y(n745) );
  INVX8 U774 ( .A(n733), .Y(n746) );
  INVX8 U775 ( .A(n733), .Y(n747) );
  INVX8 U776 ( .A(n754), .Y(n749) );
  INVX8 U777 ( .A(n754), .Y(n750) );
  INVX8 U778 ( .A(n753), .Y(n751) );
  INVX4 U779 ( .A(N20), .Y(n758) );
  MUX2X1 U780 ( .B(\mem<0> ), .A(\mem<1> ), .S(n736), .Y(n767) );
  MUX2X1 U781 ( .B(\mem<2> ), .A(\mem<3> ), .S(n744), .Y(n766) );
  MUX2X1 U782 ( .B(\mem<4> ), .A(\mem<5> ), .S(n744), .Y(n769) );
  MUX2X1 U783 ( .B(\mem<6> ), .A(\mem<7> ), .S(n738), .Y(n768) );
  MUX2X1 U784 ( .B(n769), .A(n768), .S(n749), .Y(n770) );
  MUX2X1 U785 ( .B(\mem<8> ), .A(\mem<9> ), .S(n738), .Y(n773) );
  MUX2X1 U786 ( .B(\mem<10> ), .A(\mem<11> ), .S(n738), .Y(n772) );
  MUX2X1 U787 ( .B(n773), .A(n772), .S(n749), .Y(n777) );
  MUX2X1 U788 ( .B(\mem<12> ), .A(\mem<13> ), .S(n738), .Y(n775) );
  MUX2X1 U789 ( .B(\mem<14> ), .A(\mem<15> ), .S(n738), .Y(n774) );
  MUX2X1 U790 ( .B(n775), .A(n774), .S(n749), .Y(n776) );
  MUX2X1 U791 ( .B(n777), .A(n776), .S(n757), .Y(n778) );
  MUX2X1 U792 ( .B(n779), .A(n778), .S(n761), .Y(n795) );
  MUX2X1 U793 ( .B(\mem<16> ), .A(\mem<17> ), .S(n744), .Y(n781) );
  MUX2X1 U794 ( .B(\mem<18> ), .A(\mem<19> ), .S(n738), .Y(n780) );
  MUX2X1 U795 ( .B(n781), .A(n780), .S(n749), .Y(n785) );
  MUX2X1 U796 ( .B(\mem<20> ), .A(\mem<21> ), .S(n744), .Y(n783) );
  MUX2X1 U797 ( .B(\mem<22> ), .A(\mem<23> ), .S(n744), .Y(n782) );
  MUX2X1 U798 ( .B(n783), .A(n782), .S(n749), .Y(n784) );
  MUX2X1 U799 ( .B(n785), .A(n784), .S(n757), .Y(n793) );
  MUX2X1 U800 ( .B(\mem<24> ), .A(\mem<25> ), .S(n744), .Y(n787) );
  MUX2X1 U801 ( .B(\mem<26> ), .A(\mem<27> ), .S(n744), .Y(n786) );
  MUX2X1 U802 ( .B(n787), .A(n786), .S(n749), .Y(n791) );
  MUX2X1 U803 ( .B(\mem<28> ), .A(\mem<29> ), .S(n744), .Y(n789) );
  MUX2X1 U804 ( .B(\mem<30> ), .A(\mem<31> ), .S(n744), .Y(n788) );
  MUX2X1 U805 ( .B(n789), .A(n788), .S(n749), .Y(n790) );
  MUX2X1 U806 ( .B(n791), .A(n790), .S(n757), .Y(n792) );
  MUX2X1 U807 ( .B(n793), .A(n792), .S(n761), .Y(n794) );
  MUX2X1 U808 ( .B(n795), .A(n794), .S(n763), .Y(n827) );
  MUX2X1 U809 ( .B(\mem<32> ), .A(\mem<33> ), .S(n744), .Y(n797) );
  MUX2X1 U810 ( .B(\mem<34> ), .A(\mem<35> ), .S(n744), .Y(n796) );
  MUX2X1 U811 ( .B(n797), .A(n796), .S(n749), .Y(n801) );
  MUX2X1 U812 ( .B(\mem<36> ), .A(\mem<37> ), .S(n744), .Y(n799) );
  MUX2X1 U813 ( .B(\mem<38> ), .A(\mem<39> ), .S(n744), .Y(n798) );
  MUX2X1 U814 ( .B(n799), .A(n798), .S(n749), .Y(n800) );
  MUX2X1 U815 ( .B(n801), .A(n800), .S(n757), .Y(n809) );
  MUX2X1 U816 ( .B(\mem<40> ), .A(\mem<41> ), .S(n743), .Y(n803) );
  MUX2X1 U817 ( .B(\mem<42> ), .A(\mem<43> ), .S(n744), .Y(n802) );
  MUX2X1 U818 ( .B(n803), .A(n802), .S(n749), .Y(n807) );
  MUX2X1 U819 ( .B(\mem<44> ), .A(\mem<45> ), .S(n743), .Y(n805) );
  MUX2X1 U820 ( .B(\mem<46> ), .A(\mem<47> ), .S(n743), .Y(n804) );
  MUX2X1 U821 ( .B(n805), .A(n804), .S(n749), .Y(n806) );
  MUX2X1 U822 ( .B(n807), .A(n806), .S(n757), .Y(n808) );
  MUX2X1 U823 ( .B(n809), .A(n808), .S(n761), .Y(n825) );
  MUX2X1 U824 ( .B(\mem<48> ), .A(\mem<49> ), .S(n743), .Y(n811) );
  MUX2X1 U825 ( .B(\mem<50> ), .A(\mem<51> ), .S(n743), .Y(n810) );
  MUX2X1 U826 ( .B(n811), .A(n810), .S(n749), .Y(n815) );
  MUX2X1 U827 ( .B(\mem<52> ), .A(\mem<53> ), .S(n743), .Y(n813) );
  MUX2X1 U828 ( .B(\mem<54> ), .A(\mem<55> ), .S(n743), .Y(n812) );
  MUX2X1 U829 ( .B(n813), .A(n812), .S(n750), .Y(n814) );
  MUX2X1 U830 ( .B(n815), .A(n814), .S(n757), .Y(n823) );
  MUX2X1 U831 ( .B(\mem<56> ), .A(\mem<57> ), .S(n743), .Y(n817) );
  MUX2X1 U832 ( .B(\mem<58> ), .A(\mem<59> ), .S(n743), .Y(n816) );
  MUX2X1 U833 ( .B(n817), .A(n816), .S(n749), .Y(n821) );
  MUX2X1 U834 ( .B(\mem<60> ), .A(\mem<61> ), .S(n743), .Y(n819) );
  MUX2X1 U835 ( .B(\mem<62> ), .A(\mem<63> ), .S(n743), .Y(n818) );
  MUX2X1 U836 ( .B(n819), .A(n818), .S(n750), .Y(n820) );
  MUX2X1 U837 ( .B(n821), .A(n820), .S(n757), .Y(n822) );
  MUX2X1 U838 ( .B(n823), .A(n822), .S(n761), .Y(n824) );
  MUX2X1 U839 ( .B(n825), .A(n824), .S(n763), .Y(n826) );
  MUX2X1 U840 ( .B(\mem<64> ), .A(\mem<65> ), .S(n743), .Y(n829) );
  MUX2X1 U841 ( .B(\mem<66> ), .A(\mem<67> ), .S(n742), .Y(n828) );
  MUX2X1 U842 ( .B(n829), .A(n828), .S(n749), .Y(n832) );
  MUX2X1 U843 ( .B(\mem<68> ), .A(\mem<69> ), .S(n742), .Y(n831) );
  MUX2X1 U844 ( .B(\mem<70> ), .A(\mem<71> ), .S(n742), .Y(n830) );
  MUX2X1 U845 ( .B(\mem<72> ), .A(\mem<73> ), .S(n742), .Y(n834) );
  MUX2X1 U846 ( .B(\mem<74> ), .A(\mem<75> ), .S(n742), .Y(n833) );
  MUX2X1 U847 ( .B(n834), .A(n833), .S(n752), .Y(n838) );
  MUX2X1 U848 ( .B(\mem<76> ), .A(\mem<77> ), .S(n742), .Y(n836) );
  MUX2X1 U849 ( .B(\mem<78> ), .A(\mem<79> ), .S(n742), .Y(n835) );
  MUX2X1 U850 ( .B(n836), .A(n835), .S(n752), .Y(n837) );
  MUX2X1 U851 ( .B(n838), .A(n837), .S(n756), .Y(n839) );
  MUX2X1 U852 ( .B(n840), .A(n839), .S(n761), .Y(n855) );
  MUX2X1 U853 ( .B(n842), .A(n841), .S(n750), .Y(n846) );
  MUX2X1 U854 ( .B(n844), .A(n843), .S(n749), .Y(n845) );
  MUX2X1 U855 ( .B(n846), .A(n845), .S(n756), .Y(n854) );
  MUX2X1 U856 ( .B(\mem<88> ), .A(\mem<89> ), .S(n742), .Y(n848) );
  MUX2X1 U857 ( .B(\mem<90> ), .A(\mem<91> ), .S(n741), .Y(n847) );
  MUX2X1 U858 ( .B(n848), .A(n847), .S(n750), .Y(n852) );
  MUX2X1 U859 ( .B(\mem<92> ), .A(\mem<93> ), .S(n741), .Y(n850) );
  MUX2X1 U860 ( .B(\mem<94> ), .A(\mem<95> ), .S(n741), .Y(n849) );
  MUX2X1 U861 ( .B(n850), .A(n849), .S(n749), .Y(n851) );
  MUX2X1 U862 ( .B(\mem<96> ), .A(\mem<97> ), .S(n741), .Y(n857) );
  MUX2X1 U863 ( .B(\mem<98> ), .A(\mem<99> ), .S(n741), .Y(n856) );
  MUX2X1 U864 ( .B(n857), .A(n856), .S(n752), .Y(n861) );
  MUX2X1 U865 ( .B(\mem<100> ), .A(\mem<101> ), .S(n741), .Y(n859) );
  MUX2X1 U866 ( .B(\mem<102> ), .A(\mem<103> ), .S(n741), .Y(n858) );
  MUX2X1 U867 ( .B(n859), .A(n858), .S(n750), .Y(n860) );
  MUX2X1 U868 ( .B(n861), .A(n860), .S(n756), .Y(n869) );
  MUX2X1 U869 ( .B(\mem<104> ), .A(\mem<105> ), .S(n741), .Y(n863) );
  MUX2X1 U870 ( .B(\mem<106> ), .A(\mem<107> ), .S(n741), .Y(n862) );
  MUX2X1 U871 ( .B(n863), .A(n862), .S(n750), .Y(n867) );
  MUX2X1 U872 ( .B(\mem<108> ), .A(\mem<109> ), .S(n741), .Y(n865) );
  MUX2X1 U873 ( .B(\mem<110> ), .A(\mem<111> ), .S(n741), .Y(n864) );
  MUX2X1 U874 ( .B(n865), .A(n864), .S(n750), .Y(n866) );
  MUX2X1 U875 ( .B(n867), .A(n866), .S(n756), .Y(n868) );
  MUX2X1 U876 ( .B(n869), .A(n868), .S(n761), .Y(n885) );
  MUX2X1 U877 ( .B(\mem<112> ), .A(\mem<113> ), .S(n741), .Y(n871) );
  MUX2X1 U878 ( .B(\mem<114> ), .A(\mem<115> ), .S(n740), .Y(n870) );
  MUX2X1 U879 ( .B(n871), .A(n870), .S(n750), .Y(n875) );
  MUX2X1 U880 ( .B(\mem<116> ), .A(\mem<117> ), .S(n740), .Y(n873) );
  MUX2X1 U881 ( .B(\mem<118> ), .A(\mem<119> ), .S(n740), .Y(n872) );
  MUX2X1 U882 ( .B(n873), .A(n872), .S(n750), .Y(n874) );
  MUX2X1 U883 ( .B(n875), .A(n874), .S(n756), .Y(n883) );
  MUX2X1 U884 ( .B(\mem<120> ), .A(\mem<121> ), .S(n740), .Y(n877) );
  MUX2X1 U885 ( .B(\mem<122> ), .A(\mem<123> ), .S(n740), .Y(n876) );
  MUX2X1 U886 ( .B(n877), .A(n876), .S(n750), .Y(n881) );
  MUX2X1 U887 ( .B(\mem<124> ), .A(\mem<125> ), .S(n740), .Y(n879) );
  MUX2X1 U888 ( .B(\mem<126> ), .A(\mem<127> ), .S(n740), .Y(n878) );
  MUX2X1 U889 ( .B(n879), .A(n878), .S(n750), .Y(n880) );
  MUX2X1 U890 ( .B(n881), .A(n880), .S(n756), .Y(n882) );
  MUX2X1 U891 ( .B(n883), .A(n882), .S(n761), .Y(n884) );
  MUX2X1 U892 ( .B(n887), .A(n886), .S(N23), .Y(n888) );
  MUX2X1 U893 ( .B(\mem<128> ), .A(\mem<129> ), .S(n740), .Y(n891) );
  MUX2X1 U894 ( .B(\mem<130> ), .A(\mem<131> ), .S(n740), .Y(n890) );
  MUX2X1 U895 ( .B(n891), .A(n890), .S(n750), .Y(n895) );
  MUX2X1 U896 ( .B(\mem<132> ), .A(\mem<133> ), .S(n740), .Y(n893) );
  MUX2X1 U897 ( .B(\mem<134> ), .A(\mem<135> ), .S(n740), .Y(n892) );
  MUX2X1 U898 ( .B(n893), .A(n892), .S(n750), .Y(n894) );
  MUX2X1 U899 ( .B(n895), .A(n894), .S(n756), .Y(n903) );
  MUX2X1 U900 ( .B(\mem<136> ), .A(\mem<137> ), .S(n739), .Y(n897) );
  MUX2X1 U901 ( .B(\mem<138> ), .A(\mem<139> ), .S(n739), .Y(n896) );
  MUX2X1 U902 ( .B(n897), .A(n896), .S(n750), .Y(n901) );
  MUX2X1 U903 ( .B(\mem<140> ), .A(\mem<141> ), .S(n739), .Y(n899) );
  MUX2X1 U904 ( .B(\mem<142> ), .A(\mem<143> ), .S(n739), .Y(n898) );
  MUX2X1 U905 ( .B(n899), .A(n898), .S(n750), .Y(n900) );
  MUX2X1 U906 ( .B(n901), .A(n900), .S(n756), .Y(n902) );
  MUX2X1 U907 ( .B(n903), .A(n902), .S(n761), .Y(n919) );
  MUX2X1 U908 ( .B(\mem<144> ), .A(\mem<145> ), .S(n739), .Y(n905) );
  MUX2X1 U909 ( .B(\mem<146> ), .A(\mem<147> ), .S(n739), .Y(n904) );
  MUX2X1 U910 ( .B(n905), .A(n904), .S(n751), .Y(n909) );
  MUX2X1 U911 ( .B(\mem<148> ), .A(\mem<149> ), .S(n739), .Y(n907) );
  MUX2X1 U912 ( .B(\mem<150> ), .A(\mem<151> ), .S(n739), .Y(n906) );
  MUX2X1 U913 ( .B(n907), .A(n906), .S(n751), .Y(n908) );
  MUX2X1 U914 ( .B(n909), .A(n908), .S(n756), .Y(n917) );
  MUX2X1 U915 ( .B(\mem<152> ), .A(\mem<153> ), .S(n739), .Y(n911) );
  MUX2X1 U916 ( .B(\mem<154> ), .A(\mem<155> ), .S(n739), .Y(n910) );
  MUX2X1 U917 ( .B(n911), .A(n910), .S(n751), .Y(n915) );
  MUX2X1 U918 ( .B(\mem<156> ), .A(\mem<157> ), .S(n739), .Y(n913) );
  MUX2X1 U919 ( .B(\mem<158> ), .A(\mem<159> ), .S(n739), .Y(n912) );
  MUX2X1 U920 ( .B(n913), .A(n912), .S(n751), .Y(n914) );
  MUX2X1 U921 ( .B(n915), .A(n914), .S(n756), .Y(n916) );
  MUX2X1 U922 ( .B(n917), .A(n916), .S(n761), .Y(n918) );
  MUX2X1 U923 ( .B(n919), .A(n918), .S(n763), .Y(n951) );
  MUX2X1 U924 ( .B(\mem<160> ), .A(\mem<161> ), .S(n738), .Y(n921) );
  MUX2X1 U925 ( .B(\mem<162> ), .A(\mem<163> ), .S(n738), .Y(n920) );
  MUX2X1 U926 ( .B(n921), .A(n920), .S(n751), .Y(n925) );
  MUX2X1 U927 ( .B(\mem<164> ), .A(\mem<165> ), .S(n738), .Y(n923) );
  MUX2X1 U928 ( .B(\mem<166> ), .A(\mem<167> ), .S(n738), .Y(n922) );
  MUX2X1 U929 ( .B(n923), .A(n922), .S(n751), .Y(n924) );
  MUX2X1 U930 ( .B(n925), .A(n924), .S(n755), .Y(n933) );
  MUX2X1 U931 ( .B(\mem<168> ), .A(\mem<169> ), .S(n738), .Y(n927) );
  MUX2X1 U932 ( .B(\mem<170> ), .A(\mem<171> ), .S(n738), .Y(n926) );
  MUX2X1 U933 ( .B(n927), .A(n926), .S(n751), .Y(n931) );
  MUX2X1 U934 ( .B(\mem<172> ), .A(\mem<173> ), .S(n738), .Y(n929) );
  MUX2X1 U935 ( .B(\mem<174> ), .A(\mem<175> ), .S(n738), .Y(n928) );
  MUX2X1 U936 ( .B(n929), .A(n928), .S(n751), .Y(n930) );
  MUX2X1 U937 ( .B(n931), .A(n930), .S(n755), .Y(n932) );
  MUX2X1 U938 ( .B(n933), .A(n932), .S(n761), .Y(n949) );
  MUX2X1 U939 ( .B(\mem<176> ), .A(\mem<177> ), .S(n738), .Y(n935) );
  MUX2X1 U940 ( .B(\mem<178> ), .A(\mem<179> ), .S(n738), .Y(n934) );
  MUX2X1 U941 ( .B(n935), .A(n934), .S(n751), .Y(n939) );
  MUX2X1 U942 ( .B(\mem<180> ), .A(\mem<181> ), .S(n738), .Y(n937) );
  MUX2X1 U943 ( .B(\mem<182> ), .A(\mem<183> ), .S(n738), .Y(n936) );
  MUX2X1 U944 ( .B(n937), .A(n936), .S(n751), .Y(n938) );
  MUX2X1 U945 ( .B(n939), .A(n938), .S(n755), .Y(n947) );
  MUX2X1 U946 ( .B(\mem<184> ), .A(\mem<185> ), .S(n738), .Y(n941) );
  MUX2X1 U947 ( .B(\mem<186> ), .A(\mem<187> ), .S(n744), .Y(n940) );
  MUX2X1 U948 ( .B(n941), .A(n940), .S(n751), .Y(n945) );
  MUX2X1 U949 ( .B(\mem<188> ), .A(\mem<189> ), .S(n738), .Y(n943) );
  MUX2X1 U950 ( .B(\mem<190> ), .A(\mem<191> ), .S(n743), .Y(n942) );
  MUX2X1 U951 ( .B(n943), .A(n942), .S(n751), .Y(n944) );
  MUX2X1 U952 ( .B(n945), .A(n944), .S(n755), .Y(n946) );
  MUX2X1 U953 ( .B(n947), .A(n946), .S(n761), .Y(n948) );
  MUX2X1 U954 ( .B(n949), .A(n948), .S(n763), .Y(n950) );
  MUX2X1 U955 ( .B(n951), .A(n950), .S(N23), .Y(n1015) );
  MUX2X1 U956 ( .B(\mem<192> ), .A(\mem<193> ), .S(n743), .Y(n953) );
  MUX2X1 U957 ( .B(\mem<194> ), .A(\mem<195> ), .S(n740), .Y(n952) );
  MUX2X1 U958 ( .B(n953), .A(n952), .S(n751), .Y(n957) );
  MUX2X1 U959 ( .B(\mem<196> ), .A(\mem<197> ), .S(n744), .Y(n955) );
  MUX2X1 U960 ( .B(\mem<198> ), .A(\mem<199> ), .S(n736), .Y(n954) );
  MUX2X1 U961 ( .B(n955), .A(n954), .S(n751), .Y(n956) );
  MUX2X1 U962 ( .B(n957), .A(n956), .S(n755), .Y(n965) );
  MUX2X1 U963 ( .B(\mem<200> ), .A(\mem<201> ), .S(n736), .Y(n959) );
  MUX2X1 U964 ( .B(\mem<202> ), .A(\mem<203> ), .S(n736), .Y(n958) );
  MUX2X1 U965 ( .B(n959), .A(n958), .S(n751), .Y(n963) );
  MUX2X1 U966 ( .B(\mem<204> ), .A(\mem<205> ), .S(n736), .Y(n961) );
  MUX2X1 U967 ( .B(\mem<206> ), .A(\mem<207> ), .S(n736), .Y(n960) );
  MUX2X1 U968 ( .B(n961), .A(n960), .S(n751), .Y(n962) );
  MUX2X1 U969 ( .B(n963), .A(n962), .S(n756), .Y(n964) );
  MUX2X1 U970 ( .B(n965), .A(n964), .S(N21), .Y(n981) );
  MUX2X1 U971 ( .B(\mem<208> ), .A(\mem<209> ), .S(n743), .Y(n967) );
  MUX2X1 U972 ( .B(\mem<210> ), .A(\mem<211> ), .S(n737), .Y(n966) );
  MUX2X1 U973 ( .B(n967), .A(n966), .S(n751), .Y(n971) );
  MUX2X1 U974 ( .B(\mem<212> ), .A(\mem<213> ), .S(n737), .Y(n969) );
  MUX2X1 U975 ( .B(\mem<214> ), .A(\mem<215> ), .S(n737), .Y(n968) );
  MUX2X1 U976 ( .B(n969), .A(n968), .S(n751), .Y(n970) );
  MUX2X1 U977 ( .B(n971), .A(n970), .S(n755), .Y(n979) );
  MUX2X1 U978 ( .B(\mem<216> ), .A(\mem<217> ), .S(n737), .Y(n973) );
  MUX2X1 U979 ( .B(\mem<218> ), .A(\mem<219> ), .S(n737), .Y(n972) );
  MUX2X1 U980 ( .B(n973), .A(n972), .S(n751), .Y(n977) );
  MUX2X1 U981 ( .B(\mem<220> ), .A(\mem<221> ), .S(n737), .Y(n975) );
  MUX2X1 U982 ( .B(\mem<222> ), .A(\mem<223> ), .S(n737), .Y(n974) );
  MUX2X1 U983 ( .B(n975), .A(n974), .S(n751), .Y(n976) );
  MUX2X1 U984 ( .B(n977), .A(n976), .S(n755), .Y(n978) );
  MUX2X1 U985 ( .B(n979), .A(n978), .S(N21), .Y(n980) );
  MUX2X1 U986 ( .B(n981), .A(n980), .S(n763), .Y(n1013) );
  MUX2X1 U987 ( .B(\mem<224> ), .A(\mem<225> ), .S(n737), .Y(n983) );
  MUX2X1 U988 ( .B(\mem<226> ), .A(\mem<227> ), .S(n737), .Y(n982) );
  MUX2X1 U989 ( .B(n983), .A(n982), .S(n751), .Y(n987) );
  MUX2X1 U990 ( .B(\mem<228> ), .A(\mem<229> ), .S(n737), .Y(n985) );
  MUX2X1 U991 ( .B(\mem<230> ), .A(\mem<231> ), .S(n737), .Y(n984) );
  MUX2X1 U992 ( .B(n985), .A(n984), .S(n751), .Y(n986) );
  MUX2X1 U993 ( .B(n987), .A(n986), .S(n755), .Y(n995) );
  MUX2X1 U994 ( .B(\mem<232> ), .A(\mem<233> ), .S(n737), .Y(n989) );
  MUX2X1 U995 ( .B(\mem<234> ), .A(\mem<235> ), .S(n736), .Y(n988) );
  MUX2X1 U996 ( .B(n989), .A(n988), .S(n751), .Y(n993) );
  MUX2X1 U997 ( .B(\mem<236> ), .A(\mem<237> ), .S(n736), .Y(n991) );
  MUX2X1 U998 ( .B(\mem<238> ), .A(\mem<239> ), .S(n736), .Y(n990) );
  MUX2X1 U999 ( .B(n991), .A(n990), .S(n751), .Y(n992) );
  MUX2X1 U1000 ( .B(n993), .A(n992), .S(n755), .Y(n994) );
  MUX2X1 U1001 ( .B(n995), .A(n994), .S(N21), .Y(n1011) );
  MUX2X1 U1002 ( .B(\mem<240> ), .A(\mem<241> ), .S(n736), .Y(n997) );
  MUX2X1 U1003 ( .B(\mem<242> ), .A(\mem<243> ), .S(n736), .Y(n996) );
  MUX2X1 U1004 ( .B(n997), .A(n996), .S(n752), .Y(n1001) );
  MUX2X1 U1005 ( .B(\mem<244> ), .A(\mem<245> ), .S(n736), .Y(n999) );
  MUX2X1 U1006 ( .B(\mem<246> ), .A(\mem<247> ), .S(n736), .Y(n998) );
  MUX2X1 U1007 ( .B(n999), .A(n998), .S(n752), .Y(n1000) );
  MUX2X1 U1008 ( .B(n1001), .A(n1000), .S(n755), .Y(n1009) );
  MUX2X1 U1009 ( .B(\mem<248> ), .A(\mem<249> ), .S(n736), .Y(n1003) );
  MUX2X1 U1010 ( .B(\mem<250> ), .A(\mem<251> ), .S(n736), .Y(n1002) );
  MUX2X1 U1011 ( .B(n1003), .A(n1002), .S(n752), .Y(n1007) );
  MUX2X1 U1012 ( .B(\mem<252> ), .A(\mem<253> ), .S(n736), .Y(n1005) );
  MUX2X1 U1013 ( .B(\mem<254> ), .A(\mem<255> ), .S(n736), .Y(n1004) );
  MUX2X1 U1014 ( .B(n1005), .A(n1004), .S(n752), .Y(n1006) );
  MUX2X1 U1015 ( .B(n1007), .A(n1006), .S(n755), .Y(n1008) );
  MUX2X1 U1016 ( .B(n1009), .A(n1008), .S(N21), .Y(n1010) );
  MUX2X1 U1017 ( .B(n1011), .A(n1010), .S(n763), .Y(n1012) );
  MUX2X1 U1018 ( .B(n1013), .A(n1012), .S(N23), .Y(n1014) );
  MUX2X1 U1019 ( .B(n1015), .A(n1014), .S(N24), .Y(n1016) );
  MUX2X1 U1020 ( .B(n1017), .A(n1016), .S(N25), .Y(n1018) );
  AND2X2 U1021 ( .A(n1018), .B(n10), .Y(data_out) );
endmodule


module memc_Size16_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2070), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2071), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2072), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2073), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2074), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2075), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2076), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2077), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2078), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2079), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2080), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2081), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2082), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2083), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2084), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2085), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2086), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2087), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2088), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2089), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2090), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2091), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2092), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2093), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2094), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2095), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2096), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2097), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2098), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2099), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2100), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2101), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2102), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2103), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2104), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2105), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2106), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2107), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2108), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2109), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2110), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2111), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2112), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2113), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2114), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2115), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2116), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2117), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2118), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2119), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2120), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2121), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2122), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2123), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2124), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2125), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2126), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2127), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2128), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2129), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2130), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2131), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2132), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2133), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2134), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2135), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2136), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2137), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2138), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2139), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2140), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2141), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2142), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2143), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2144), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2145), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2146), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2147), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2148), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2149), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2150), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2151), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2152), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2153), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2154), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2155), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2156), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2157), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2158), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2159), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2160), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2161), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2162), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2163), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2164), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2165), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2166), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2167), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2168), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2169), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2170), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2171), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2172), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2173), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2174), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2175), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2176), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2177), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2178), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2179), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2180), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2181), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2182), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2183), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2184), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2185), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2186), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2187), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2188), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2189), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2190), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2191), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2192), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2193), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2194), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2195), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2196), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2197), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2198), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2199), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2200), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2201), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2202), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2203), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2204), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2205), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2206), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2207), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2208), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2209), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2210), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2211), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2212), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2213), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2214), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2215), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2216), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2217), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2218), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2219), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2220), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2221), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2222), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2223), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2224), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2225), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2226), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2227), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2228), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2229), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2230), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2231), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2232), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2233), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2234), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2235), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2236), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2237), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2238), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2239), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2240), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2241), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2242), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2243), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2244), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2245), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2246), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2247), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2248), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2249), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2250), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2251), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2252), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2253), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2254), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2255), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2256), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2257), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2258), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2259), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2260), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2261), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2262), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2263), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2264), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2265), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2266), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2267), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2268), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2269), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2270), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2271), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2272), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2273), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2274), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2275), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2276), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2277), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2278), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2279), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2280), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2281), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2282), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2283), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2284), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2285), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2286), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2287), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2288), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2289), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2290), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2291), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2292), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2293), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2294), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2295), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2296), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2297), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2298), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2299), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2300), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2301), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2302), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2303), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2304), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2305), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2306), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2307), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2308), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2309), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2310), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2311), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2312), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2313), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2314), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2315), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2316), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2317), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2318), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2319), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2320), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2321), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2322), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2323), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2324), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2325), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2326), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2327), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2328), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2329), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2330), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2331), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2332), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2333), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2334), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2335), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2336), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2337), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2338), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2339), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2340), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2341), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2342), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2343), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2344), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2345), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2346), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2347), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2348), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2349), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2350), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2351), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2352), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2353), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2354), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2355), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2356), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2357), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2358), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2359), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2360), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2361), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2362), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2363), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2364), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2365), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2366), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2367), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2368), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2369), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2370), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2371), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2372), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2373), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2374), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2375), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2376), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2377), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2378), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2379), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2380), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2381), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2382), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2383), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2384), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2385), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2386), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2387), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2388), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2389), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2390), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2391), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2392), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2393), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2394), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2395), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2396), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2397), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2398), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2399), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2400), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2401), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2402), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2403), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2404), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2405), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2406), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2407), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2408), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2409), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2410), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2411), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2412), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2413), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2414), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2415), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2416), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2417), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2418), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2419), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2420), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2421), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2422), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2423), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2424), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2425), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2426), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2427), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2428), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2429), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2430), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2431), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2432), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2433), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2434), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2435), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2436), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2437), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2438), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2439), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2440), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2441), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2442), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2443), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2444), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2445), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2446), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2447), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2448), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2449), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2450), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2451), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2452), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2453), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2454), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2455), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2456), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2457), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2458), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2459), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2460), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2461), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2462), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2463), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2464), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2465), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2466), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2467), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2468), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2469), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2470), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2471), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2472), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2473), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2474), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2475), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2476), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2477), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2478), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2479), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2480), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2481), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2482), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2483), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2484), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2485), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2486), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2487), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2488), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2489), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2490), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2491), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2492), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2493), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2494), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2495), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2496), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2497), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2498), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2499), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2500), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2501), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2502), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2503), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2504), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2505), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2506), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2507), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2508), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2509), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2510), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2511), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2512), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2513), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2514), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2515), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2516), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2517), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2518), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2519), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2520), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2521), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2522), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2523), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2524), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2525), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2526), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2527), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2528), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2529), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2530), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2531), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2532), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2533), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2534), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2535), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2536), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2537), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2538), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2539), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2540), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2541), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2542), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2543), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2544), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2545), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2546), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2547), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2548), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2549), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2550), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2551), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2552), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2553), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2554), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2555), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2556), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2557), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2558), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2559), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2560), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2561), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2562), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2563), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2564), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2565), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2566), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2567), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2568), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2569), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2570), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2571), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2572), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2573), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2574), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2575), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2576), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2577), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2578), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2579), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2580), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2581), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2582) );
  AND2X1 U2 ( .A(\data_in<10> ), .B(n1740), .Y(n476) );
  AND2X2 U3 ( .A(\data_in<9> ), .B(n1740), .Y(n475) );
  AND2X2 U4 ( .A(\data_in<8> ), .B(n1740), .Y(n474) );
  AND2X1 U5 ( .A(\data_in<7> ), .B(n1740), .Y(n473) );
  AND2X1 U6 ( .A(\data_in<6> ), .B(n1740), .Y(n472) );
  AND2X2 U7 ( .A(\data_in<5> ), .B(n1740), .Y(n471) );
  AND2X2 U8 ( .A(\data_in<4> ), .B(n1740), .Y(n470) );
  AND2X1 U9 ( .A(\data_in<3> ), .B(n1740), .Y(n469) );
  AND2X1 U10 ( .A(\data_in<2> ), .B(n1740), .Y(n468) );
  AND2X2 U11 ( .A(\data_in<1> ), .B(n1740), .Y(n467) );
  AND2X2 U12 ( .A(\data_in<0> ), .B(n1740), .Y(n466) );
  AND2X1 U13 ( .A(\data_in<14> ), .B(n1739), .Y(n494) );
  AND2X1 U14 ( .A(\data_in<12> ), .B(n1739), .Y(n492) );
  INVX1 U15 ( .A(n1654), .Y(n1655) );
  INVX1 U16 ( .A(n1654), .Y(n1656) );
  INVX2 U17 ( .A(n1653), .Y(n1661) );
  INVX2 U18 ( .A(n1671), .Y(n1652) );
  INVX1 U19 ( .A(n1671), .Y(n1653) );
  INVX2 U20 ( .A(n1652), .Y(n1665) );
  INVX2 U21 ( .A(n1653), .Y(n1663) );
  INVX2 U22 ( .A(n1653), .Y(n1662) );
  INVX1 U23 ( .A(n1654), .Y(n1658) );
  INVX1 U24 ( .A(n1654), .Y(n1670) );
  INVX1 U25 ( .A(n1654), .Y(n1669) );
  INVX1 U26 ( .A(n1764), .Y(n1667) );
  INVX1 U27 ( .A(n1764), .Y(n1666) );
  INVX1 U28 ( .A(n1769), .Y(n1633) );
  INVX1 U29 ( .A(n1769), .Y(n1631) );
  INVX1 U30 ( .A(n1769), .Y(n1632) );
  INVX1 U31 ( .A(n1615), .Y(N31) );
  INVX1 U32 ( .A(N10), .Y(n1654) );
  INVX1 U33 ( .A(n1639), .Y(n1640) );
  INVX1 U34 ( .A(n1639), .Y(n1642) );
  INVX1 U35 ( .A(n1638), .Y(n1645) );
  INVX1 U36 ( .A(n1651), .Y(n1647) );
  INVX1 U37 ( .A(n1651), .Y(n1648) );
  INVX1 U38 ( .A(n1639), .Y(n1649) );
  INVX2 U39 ( .A(n1654), .Y(n1657) );
  INVX1 U40 ( .A(n1638), .Y(n1650) );
  INVX1 U41 ( .A(n1639), .Y(n1641) );
  INVX1 U42 ( .A(n1638), .Y(n1643) );
  INVX1 U43 ( .A(n1638), .Y(n1644) );
  INVX1 U44 ( .A(n1651), .Y(n1646) );
  INVX1 U45 ( .A(n1626), .Y(N20) );
  INVX1 U46 ( .A(n1628), .Y(N18) );
  INVX1 U47 ( .A(n1614), .Y(N32) );
  INVX1 U48 ( .A(n1616), .Y(N30) );
  INVX1 U49 ( .A(n1617), .Y(N29) );
  INVX1 U50 ( .A(n1618), .Y(N28) );
  INVX1 U51 ( .A(n1619), .Y(N27) );
  INVX1 U52 ( .A(n1620), .Y(N26) );
  INVX1 U53 ( .A(n1621), .Y(N25) );
  INVX1 U54 ( .A(n1622), .Y(N24) );
  INVX1 U55 ( .A(n1623), .Y(N23) );
  INVX1 U56 ( .A(n1624), .Y(N22) );
  INVX1 U57 ( .A(n1625), .Y(N21) );
  INVX1 U58 ( .A(n1627), .Y(N19) );
  INVX1 U59 ( .A(n1629), .Y(N17) );
  INVX2 U60 ( .A(n1767), .Y(n1634) );
  INVX1 U61 ( .A(n1764), .Y(n1671) );
  INVX1 U62 ( .A(N12), .Y(n1767) );
  INVX1 U63 ( .A(n1767), .Y(n1636) );
  INVX1 U64 ( .A(n1767), .Y(n1637) );
  INVX1 U65 ( .A(n1767), .Y(n1635) );
  INVX1 U66 ( .A(n1765), .Y(n1651) );
  INVX1 U67 ( .A(n1765), .Y(n1638) );
  INVX1 U68 ( .A(n1765), .Y(n1639) );
  INVX1 U69 ( .A(N13), .Y(n1769) );
  INVX1 U70 ( .A(N14), .Y(n1771) );
  INVX1 U71 ( .A(n1771), .Y(n1630) );
  INVX1 U72 ( .A(n496), .Y(n1686) );
  INVX1 U73 ( .A(n497), .Y(n1703) );
  INVX1 U74 ( .A(rst), .Y(n1772) );
  BUFX2 U75 ( .A(n505), .Y(n1672) );
  AND2X2 U76 ( .A(\mem<31><8> ), .B(n1673), .Y(n1) );
  INVX1 U77 ( .A(n1), .Y(n2) );
  AND2X2 U78 ( .A(\mem<31><9> ), .B(n1673), .Y(n3) );
  INVX1 U79 ( .A(n3), .Y(n4) );
  AND2X2 U80 ( .A(\mem<31><10> ), .B(n1673), .Y(n5) );
  INVX1 U81 ( .A(n5), .Y(n6) );
  AND2X2 U82 ( .A(\mem<31><11> ), .B(n1673), .Y(n7) );
  INVX1 U83 ( .A(n7), .Y(n8) );
  AND2X2 U84 ( .A(\mem<31><12> ), .B(n1673), .Y(n9) );
  INVX1 U85 ( .A(n9), .Y(n10) );
  AND2X2 U86 ( .A(\mem<31><13> ), .B(n1673), .Y(n11) );
  INVX1 U87 ( .A(n11), .Y(n12) );
  AND2X2 U88 ( .A(\mem<31><14> ), .B(n1673), .Y(n13) );
  INVX1 U89 ( .A(n13), .Y(n14) );
  AND2X2 U90 ( .A(\mem<31><15> ), .B(n1673), .Y(n15) );
  INVX1 U91 ( .A(n15), .Y(n16) );
  BUFX2 U92 ( .A(n505), .Y(n1673) );
  BUFX2 U93 ( .A(n509), .Y(n1674) );
  AND2X2 U94 ( .A(\mem<30><8> ), .B(n1675), .Y(n17) );
  INVX1 U95 ( .A(n17), .Y(n18) );
  AND2X2 U96 ( .A(\mem<30><9> ), .B(n1675), .Y(n19) );
  INVX1 U97 ( .A(n19), .Y(n20) );
  AND2X2 U98 ( .A(\mem<30><10> ), .B(n1675), .Y(n21) );
  INVX1 U99 ( .A(n21), .Y(n22) );
  AND2X2 U100 ( .A(\mem<30><11> ), .B(n1675), .Y(n23) );
  INVX1 U101 ( .A(n23), .Y(n24) );
  AND2X2 U102 ( .A(\mem<30><12> ), .B(n1675), .Y(n25) );
  INVX1 U103 ( .A(n25), .Y(n26) );
  AND2X2 U104 ( .A(\mem<30><13> ), .B(n1675), .Y(n27) );
  INVX1 U105 ( .A(n27), .Y(n28) );
  AND2X2 U106 ( .A(\mem<30><14> ), .B(n1675), .Y(n29) );
  INVX1 U107 ( .A(n29), .Y(n30) );
  AND2X2 U108 ( .A(\mem<30><15> ), .B(n1675), .Y(n31) );
  INVX1 U109 ( .A(n31), .Y(n32) );
  BUFX2 U110 ( .A(n509), .Y(n1675) );
  BUFX2 U111 ( .A(n513), .Y(n1676) );
  AND2X2 U112 ( .A(\mem<29><8> ), .B(n1677), .Y(n33) );
  INVX1 U113 ( .A(n33), .Y(n34) );
  AND2X2 U114 ( .A(\mem<29><9> ), .B(n1677), .Y(n35) );
  INVX1 U115 ( .A(n35), .Y(n36) );
  AND2X2 U116 ( .A(\mem<29><10> ), .B(n1677), .Y(n37) );
  INVX1 U117 ( .A(n37), .Y(n38) );
  AND2X2 U118 ( .A(\mem<29><11> ), .B(n1677), .Y(n39) );
  INVX1 U119 ( .A(n39), .Y(n40) );
  AND2X2 U120 ( .A(\mem<29><12> ), .B(n1677), .Y(n41) );
  INVX1 U121 ( .A(n41), .Y(n42) );
  AND2X2 U122 ( .A(\mem<29><13> ), .B(n1677), .Y(n43) );
  INVX1 U123 ( .A(n43), .Y(n44) );
  AND2X2 U124 ( .A(\mem<29><14> ), .B(n1677), .Y(n45) );
  INVX1 U125 ( .A(n45), .Y(n46) );
  AND2X2 U126 ( .A(\mem<29><15> ), .B(n1677), .Y(n47) );
  INVX1 U127 ( .A(n47), .Y(n48) );
  BUFX2 U128 ( .A(n513), .Y(n1677) );
  BUFX2 U129 ( .A(n517), .Y(n1678) );
  AND2X2 U130 ( .A(\mem<28><8> ), .B(n1679), .Y(n49) );
  INVX1 U131 ( .A(n49), .Y(n50) );
  AND2X2 U132 ( .A(\mem<28><9> ), .B(n1679), .Y(n51) );
  INVX1 U133 ( .A(n51), .Y(n52) );
  AND2X2 U134 ( .A(\mem<28><10> ), .B(n1679), .Y(n53) );
  INVX1 U135 ( .A(n53), .Y(n54) );
  AND2X2 U136 ( .A(\mem<28><11> ), .B(n1679), .Y(n55) );
  INVX1 U137 ( .A(n55), .Y(n56) );
  AND2X2 U138 ( .A(\mem<28><12> ), .B(n1679), .Y(n57) );
  INVX1 U139 ( .A(n57), .Y(n58) );
  AND2X2 U140 ( .A(\mem<28><13> ), .B(n1679), .Y(n59) );
  INVX1 U141 ( .A(n59), .Y(n60) );
  AND2X2 U142 ( .A(\mem<28><14> ), .B(n1679), .Y(n61) );
  INVX1 U143 ( .A(n61), .Y(n62) );
  AND2X2 U144 ( .A(\mem<28><15> ), .B(n1679), .Y(n63) );
  INVX1 U145 ( .A(n63), .Y(n64) );
  BUFX2 U146 ( .A(n517), .Y(n1679) );
  BUFX2 U147 ( .A(n521), .Y(n1680) );
  AND2X2 U148 ( .A(\mem<27><8> ), .B(n1681), .Y(n65) );
  INVX1 U149 ( .A(n65), .Y(n66) );
  AND2X2 U150 ( .A(\mem<27><9> ), .B(n1681), .Y(n67) );
  INVX1 U151 ( .A(n67), .Y(n68) );
  AND2X2 U152 ( .A(\mem<27><10> ), .B(n1681), .Y(n69) );
  INVX1 U153 ( .A(n69), .Y(n70) );
  AND2X2 U154 ( .A(\mem<27><11> ), .B(n1681), .Y(n71) );
  INVX1 U155 ( .A(n71), .Y(n72) );
  AND2X2 U156 ( .A(\mem<27><12> ), .B(n1681), .Y(n73) );
  INVX1 U157 ( .A(n73), .Y(n74) );
  AND2X2 U158 ( .A(\mem<27><13> ), .B(n1681), .Y(n75) );
  INVX1 U159 ( .A(n75), .Y(n76) );
  AND2X2 U160 ( .A(\mem<27><14> ), .B(n1681), .Y(n77) );
  INVX1 U161 ( .A(n77), .Y(n78) );
  AND2X2 U162 ( .A(\mem<27><15> ), .B(n1681), .Y(n79) );
  INVX1 U163 ( .A(n79), .Y(n80) );
  BUFX2 U164 ( .A(n521), .Y(n1681) );
  BUFX2 U165 ( .A(n525), .Y(n1682) );
  AND2X2 U166 ( .A(\mem<26><8> ), .B(n1683), .Y(n81) );
  INVX1 U167 ( .A(n81), .Y(n82) );
  AND2X2 U168 ( .A(\mem<26><9> ), .B(n1683), .Y(n83) );
  INVX1 U169 ( .A(n83), .Y(n84) );
  AND2X2 U170 ( .A(\mem<26><10> ), .B(n1683), .Y(n85) );
  INVX1 U171 ( .A(n85), .Y(n86) );
  AND2X2 U172 ( .A(\mem<26><11> ), .B(n1683), .Y(n87) );
  INVX1 U173 ( .A(n87), .Y(n88) );
  AND2X2 U174 ( .A(\mem<26><12> ), .B(n1683), .Y(n89) );
  INVX1 U175 ( .A(n89), .Y(n90) );
  AND2X2 U176 ( .A(\mem<26><13> ), .B(n1683), .Y(n91) );
  INVX1 U177 ( .A(n91), .Y(n92) );
  AND2X2 U178 ( .A(\mem<26><14> ), .B(n1683), .Y(n93) );
  INVX1 U179 ( .A(n93), .Y(n94) );
  AND2X2 U180 ( .A(\mem<26><15> ), .B(n1683), .Y(n95) );
  INVX1 U181 ( .A(n95), .Y(n96) );
  BUFX2 U182 ( .A(n525), .Y(n1683) );
  BUFX2 U183 ( .A(n529), .Y(n1684) );
  AND2X2 U184 ( .A(\mem<25><8> ), .B(n1685), .Y(n97) );
  INVX1 U185 ( .A(n97), .Y(n98) );
  AND2X2 U186 ( .A(\mem<25><9> ), .B(n1685), .Y(n99) );
  INVX1 U187 ( .A(n99), .Y(n100) );
  AND2X2 U188 ( .A(\mem<25><10> ), .B(n1685), .Y(n101) );
  INVX1 U189 ( .A(n101), .Y(n102) );
  AND2X2 U190 ( .A(\mem<25><11> ), .B(n1685), .Y(n103) );
  INVX1 U191 ( .A(n103), .Y(n104) );
  AND2X2 U192 ( .A(\mem<25><12> ), .B(n1685), .Y(n105) );
  INVX1 U193 ( .A(n105), .Y(n106) );
  AND2X2 U194 ( .A(\mem<25><13> ), .B(n1685), .Y(n107) );
  INVX1 U195 ( .A(n107), .Y(n108) );
  AND2X2 U196 ( .A(\mem<25><14> ), .B(n1685), .Y(n109) );
  INVX1 U197 ( .A(n109), .Y(n110) );
  AND2X2 U198 ( .A(\mem<25><15> ), .B(n1685), .Y(n111) );
  INVX1 U199 ( .A(n111), .Y(n112) );
  BUFX2 U200 ( .A(n529), .Y(n1685) );
  BUFX2 U201 ( .A(n531), .Y(n1687) );
  AND2X2 U202 ( .A(\mem<24><8> ), .B(n1688), .Y(n113) );
  INVX1 U203 ( .A(n113), .Y(n114) );
  AND2X2 U204 ( .A(\mem<24><9> ), .B(n1688), .Y(n115) );
  INVX1 U205 ( .A(n115), .Y(n116) );
  AND2X2 U206 ( .A(\mem<24><10> ), .B(n1688), .Y(n117) );
  INVX1 U207 ( .A(n117), .Y(n118) );
  AND2X2 U208 ( .A(\mem<24><11> ), .B(n1688), .Y(n119) );
  INVX1 U209 ( .A(n119), .Y(n120) );
  AND2X2 U210 ( .A(\mem<24><12> ), .B(n1688), .Y(n121) );
  INVX1 U211 ( .A(n121), .Y(n122) );
  AND2X2 U212 ( .A(\mem<24><13> ), .B(n1688), .Y(n123) );
  INVX1 U213 ( .A(n123), .Y(n124) );
  AND2X2 U214 ( .A(\mem<24><14> ), .B(n1688), .Y(n125) );
  INVX1 U215 ( .A(n125), .Y(n126) );
  AND2X2 U216 ( .A(\mem<24><15> ), .B(n1688), .Y(n127) );
  INVX1 U217 ( .A(n127), .Y(n128) );
  BUFX2 U218 ( .A(n531), .Y(n1688) );
  BUFX2 U219 ( .A(n535), .Y(n1689) );
  AND2X2 U220 ( .A(\mem<23><8> ), .B(n1690), .Y(n129) );
  INVX1 U221 ( .A(n129), .Y(n130) );
  AND2X2 U222 ( .A(\mem<23><9> ), .B(n1690), .Y(n131) );
  INVX1 U223 ( .A(n131), .Y(n132) );
  AND2X2 U224 ( .A(\mem<23><10> ), .B(n1690), .Y(n133) );
  INVX1 U225 ( .A(n133), .Y(n134) );
  AND2X2 U226 ( .A(\mem<23><11> ), .B(n1690), .Y(n135) );
  INVX1 U227 ( .A(n135), .Y(n136) );
  AND2X2 U228 ( .A(\mem<23><12> ), .B(n1690), .Y(n137) );
  INVX1 U229 ( .A(n137), .Y(n138) );
  AND2X2 U230 ( .A(\mem<23><13> ), .B(n1690), .Y(n139) );
  INVX1 U231 ( .A(n139), .Y(n140) );
  AND2X2 U232 ( .A(\mem<23><14> ), .B(n1690), .Y(n141) );
  INVX1 U233 ( .A(n141), .Y(n142) );
  AND2X2 U234 ( .A(\mem<23><15> ), .B(n1690), .Y(n143) );
  INVX1 U235 ( .A(n143), .Y(n144) );
  BUFX2 U236 ( .A(n535), .Y(n1690) );
  BUFX2 U237 ( .A(n539), .Y(n1691) );
  AND2X2 U238 ( .A(\mem<22><8> ), .B(n1692), .Y(n145) );
  INVX1 U239 ( .A(n145), .Y(n146) );
  AND2X2 U240 ( .A(\mem<22><9> ), .B(n1692), .Y(n147) );
  INVX1 U241 ( .A(n147), .Y(n148) );
  AND2X2 U242 ( .A(\mem<22><10> ), .B(n1692), .Y(n149) );
  INVX1 U243 ( .A(n149), .Y(n150) );
  AND2X2 U244 ( .A(\mem<22><11> ), .B(n1692), .Y(n151) );
  INVX1 U245 ( .A(n151), .Y(n152) );
  AND2X2 U246 ( .A(\mem<22><12> ), .B(n1692), .Y(n153) );
  INVX1 U247 ( .A(n153), .Y(n154) );
  AND2X2 U248 ( .A(\mem<22><13> ), .B(n1692), .Y(n155) );
  INVX1 U249 ( .A(n155), .Y(n156) );
  AND2X2 U250 ( .A(\mem<22><14> ), .B(n1692), .Y(n157) );
  INVX1 U251 ( .A(n157), .Y(n158) );
  AND2X2 U252 ( .A(\mem<22><15> ), .B(n1692), .Y(n159) );
  INVX1 U253 ( .A(n159), .Y(n160) );
  BUFX2 U254 ( .A(n539), .Y(n1692) );
  BUFX2 U255 ( .A(n543), .Y(n1693) );
  AND2X2 U256 ( .A(\mem<21><8> ), .B(n1694), .Y(n161) );
  INVX1 U257 ( .A(n161), .Y(n162) );
  AND2X2 U258 ( .A(\mem<21><9> ), .B(n1694), .Y(n163) );
  INVX1 U259 ( .A(n163), .Y(n164) );
  AND2X2 U260 ( .A(\mem<21><10> ), .B(n1694), .Y(n165) );
  INVX1 U261 ( .A(n165), .Y(n166) );
  AND2X2 U262 ( .A(\mem<21><11> ), .B(n1694), .Y(n167) );
  INVX1 U263 ( .A(n167), .Y(n168) );
  AND2X2 U264 ( .A(\mem<21><12> ), .B(n1694), .Y(n169) );
  INVX1 U265 ( .A(n169), .Y(n170) );
  AND2X2 U266 ( .A(\mem<21><13> ), .B(n1694), .Y(n171) );
  INVX1 U267 ( .A(n171), .Y(n172) );
  AND2X2 U268 ( .A(\mem<21><14> ), .B(n1694), .Y(n173) );
  INVX1 U269 ( .A(n173), .Y(n174) );
  AND2X2 U270 ( .A(\mem<21><15> ), .B(n1694), .Y(n175) );
  INVX1 U271 ( .A(n175), .Y(n176) );
  BUFX2 U272 ( .A(n543), .Y(n1694) );
  BUFX2 U273 ( .A(n547), .Y(n1695) );
  AND2X2 U274 ( .A(\mem<20><8> ), .B(n1696), .Y(n177) );
  INVX1 U275 ( .A(n177), .Y(n178) );
  AND2X2 U276 ( .A(\mem<20><9> ), .B(n1696), .Y(n179) );
  INVX1 U277 ( .A(n179), .Y(n180) );
  AND2X2 U278 ( .A(\mem<20><10> ), .B(n1696), .Y(n181) );
  INVX1 U279 ( .A(n181), .Y(n182) );
  AND2X2 U280 ( .A(\mem<20><11> ), .B(n1696), .Y(n183) );
  INVX1 U281 ( .A(n183), .Y(n184) );
  AND2X2 U282 ( .A(\mem<20><12> ), .B(n1696), .Y(n185) );
  INVX1 U283 ( .A(n185), .Y(n186) );
  AND2X2 U284 ( .A(\mem<20><13> ), .B(n1696), .Y(n187) );
  INVX1 U285 ( .A(n187), .Y(n188) );
  AND2X2 U286 ( .A(\mem<20><14> ), .B(n1696), .Y(n189) );
  INVX1 U287 ( .A(n189), .Y(n190) );
  AND2X2 U288 ( .A(\mem<20><15> ), .B(n1696), .Y(n191) );
  INVX1 U289 ( .A(n191), .Y(n192) );
  BUFX2 U290 ( .A(n547), .Y(n1696) );
  BUFX2 U291 ( .A(n551), .Y(n1697) );
  AND2X2 U292 ( .A(\mem<19><8> ), .B(n1698), .Y(n193) );
  INVX1 U293 ( .A(n193), .Y(n194) );
  AND2X2 U294 ( .A(\mem<19><9> ), .B(n1698), .Y(n195) );
  INVX1 U295 ( .A(n195), .Y(n196) );
  AND2X2 U296 ( .A(\mem<19><10> ), .B(n1698), .Y(n197) );
  INVX1 U297 ( .A(n197), .Y(n198) );
  AND2X2 U298 ( .A(\mem<19><11> ), .B(n1698), .Y(n199) );
  INVX1 U299 ( .A(n199), .Y(n200) );
  AND2X2 U300 ( .A(\mem<19><12> ), .B(n1698), .Y(n201) );
  INVX1 U301 ( .A(n201), .Y(n202) );
  AND2X2 U302 ( .A(\mem<19><13> ), .B(n1698), .Y(n203) );
  INVX1 U303 ( .A(n203), .Y(n204) );
  AND2X2 U304 ( .A(\mem<19><14> ), .B(n1698), .Y(n205) );
  INVX1 U305 ( .A(n205), .Y(n206) );
  AND2X2 U306 ( .A(\mem<19><15> ), .B(n1698), .Y(n207) );
  INVX1 U307 ( .A(n207), .Y(n208) );
  BUFX2 U308 ( .A(n551), .Y(n1698) );
  BUFX2 U309 ( .A(n555), .Y(n1699) );
  AND2X2 U310 ( .A(\mem<18><8> ), .B(n1700), .Y(n209) );
  INVX1 U311 ( .A(n209), .Y(n210) );
  AND2X2 U312 ( .A(\mem<18><9> ), .B(n1700), .Y(n211) );
  INVX1 U313 ( .A(n211), .Y(n212) );
  AND2X2 U314 ( .A(\mem<18><10> ), .B(n1700), .Y(n213) );
  INVX1 U315 ( .A(n213), .Y(n215) );
  AND2X2 U316 ( .A(\mem<18><11> ), .B(n1700), .Y(n216) );
  INVX1 U317 ( .A(n216), .Y(n217) );
  AND2X2 U318 ( .A(\mem<18><12> ), .B(n1700), .Y(n218) );
  INVX1 U319 ( .A(n218), .Y(n219) );
  AND2X2 U320 ( .A(\mem<18><13> ), .B(n1700), .Y(n220) );
  INVX1 U321 ( .A(n220), .Y(n221) );
  AND2X2 U322 ( .A(\mem<18><14> ), .B(n1700), .Y(n222) );
  INVX1 U323 ( .A(n222), .Y(n223) );
  AND2X2 U324 ( .A(\mem<18><15> ), .B(n1700), .Y(n224) );
  INVX1 U325 ( .A(n224), .Y(n225) );
  BUFX2 U326 ( .A(n555), .Y(n1700) );
  BUFX2 U327 ( .A(n559), .Y(n1701) );
  AND2X2 U328 ( .A(\mem<17><8> ), .B(n1702), .Y(n226) );
  INVX1 U329 ( .A(n226), .Y(n227) );
  AND2X2 U330 ( .A(\mem<17><9> ), .B(n1702), .Y(n228) );
  INVX1 U331 ( .A(n228), .Y(n229) );
  AND2X2 U332 ( .A(\mem<17><10> ), .B(n1702), .Y(n230) );
  INVX1 U333 ( .A(n230), .Y(n231) );
  AND2X2 U334 ( .A(\mem<17><11> ), .B(n1702), .Y(n232) );
  INVX1 U335 ( .A(n232), .Y(n233) );
  AND2X2 U336 ( .A(\mem<17><12> ), .B(n1702), .Y(n234) );
  INVX1 U337 ( .A(n234), .Y(n235) );
  AND2X2 U338 ( .A(\mem<17><13> ), .B(n1702), .Y(n236) );
  INVX1 U339 ( .A(n236), .Y(n237) );
  AND2X2 U340 ( .A(\mem<17><14> ), .B(n1702), .Y(n238) );
  INVX1 U341 ( .A(n238), .Y(n239) );
  AND2X2 U342 ( .A(\mem<17><15> ), .B(n1702), .Y(n240) );
  INVX1 U343 ( .A(n240), .Y(n241) );
  BUFX2 U344 ( .A(n559), .Y(n1702) );
  BUFX2 U345 ( .A(n561), .Y(n1704) );
  AND2X2 U346 ( .A(\mem<16><8> ), .B(n1705), .Y(n242) );
  INVX1 U347 ( .A(n242), .Y(n243) );
  AND2X2 U348 ( .A(\mem<16><9> ), .B(n1705), .Y(n244) );
  INVX1 U349 ( .A(n244), .Y(n245) );
  AND2X2 U350 ( .A(\mem<16><10> ), .B(n1705), .Y(n246) );
  INVX1 U351 ( .A(n246), .Y(n247) );
  AND2X2 U352 ( .A(\mem<16><11> ), .B(n1705), .Y(n248) );
  INVX1 U353 ( .A(n248), .Y(n249) );
  AND2X2 U354 ( .A(\mem<16><12> ), .B(n1705), .Y(n250) );
  INVX1 U355 ( .A(n250), .Y(n251) );
  AND2X2 U356 ( .A(\mem<16><13> ), .B(n1705), .Y(n252) );
  INVX1 U357 ( .A(n252), .Y(n253) );
  AND2X2 U358 ( .A(\mem<16><14> ), .B(n1705), .Y(n254) );
  INVX1 U359 ( .A(n254), .Y(n255) );
  AND2X2 U360 ( .A(\mem<16><15> ), .B(n1705), .Y(n256) );
  INVX1 U361 ( .A(n256), .Y(n257) );
  BUFX2 U362 ( .A(n561), .Y(n1705) );
  BUFX2 U363 ( .A(n565), .Y(n1706) );
  AND2X2 U364 ( .A(\mem<15><8> ), .B(n1707), .Y(n258) );
  INVX1 U365 ( .A(n258), .Y(n259) );
  AND2X2 U366 ( .A(\mem<15><9> ), .B(n1707), .Y(n260) );
  INVX1 U367 ( .A(n260), .Y(n261) );
  AND2X2 U368 ( .A(\mem<15><10> ), .B(n1707), .Y(n262) );
  INVX1 U369 ( .A(n262), .Y(n263) );
  AND2X2 U370 ( .A(\mem<15><11> ), .B(n1707), .Y(n264) );
  INVX1 U371 ( .A(n264), .Y(n265) );
  AND2X2 U372 ( .A(\mem<15><12> ), .B(n1707), .Y(n266) );
  INVX1 U373 ( .A(n266), .Y(n267) );
  AND2X2 U374 ( .A(\mem<15><13> ), .B(n1707), .Y(n268) );
  INVX1 U375 ( .A(n268), .Y(n269) );
  AND2X2 U376 ( .A(\mem<15><14> ), .B(n1707), .Y(n270) );
  INVX1 U377 ( .A(n270), .Y(n271) );
  AND2X2 U378 ( .A(\mem<15><15> ), .B(n1707), .Y(n272) );
  INVX1 U379 ( .A(n272), .Y(n273) );
  BUFX2 U380 ( .A(n565), .Y(n1707) );
  BUFX2 U381 ( .A(n569), .Y(n1708) );
  AND2X2 U382 ( .A(\mem<14><8> ), .B(n1709), .Y(n274) );
  INVX1 U383 ( .A(n274), .Y(n275) );
  AND2X2 U384 ( .A(\mem<14><9> ), .B(n1709), .Y(n276) );
  INVX1 U385 ( .A(n276), .Y(n277) );
  AND2X2 U386 ( .A(\mem<14><10> ), .B(n1709), .Y(n278) );
  INVX1 U387 ( .A(n278), .Y(n279) );
  AND2X2 U388 ( .A(\mem<14><11> ), .B(n1709), .Y(n280) );
  INVX1 U389 ( .A(n280), .Y(n281) );
  AND2X2 U390 ( .A(\mem<14><12> ), .B(n1709), .Y(n282) );
  INVX1 U391 ( .A(n282), .Y(n283) );
  AND2X2 U392 ( .A(\mem<14><13> ), .B(n1709), .Y(n284) );
  INVX1 U393 ( .A(n284), .Y(n285) );
  AND2X2 U394 ( .A(\mem<14><14> ), .B(n1709), .Y(n286) );
  INVX1 U395 ( .A(n286), .Y(n287) );
  AND2X2 U396 ( .A(\mem<14><15> ), .B(n1709), .Y(n288) );
  INVX1 U397 ( .A(n288), .Y(n289) );
  BUFX2 U398 ( .A(n569), .Y(n1709) );
  BUFX2 U399 ( .A(n573), .Y(n1710) );
  AND2X2 U400 ( .A(\mem<13><8> ), .B(n1711), .Y(n290) );
  INVX1 U401 ( .A(n290), .Y(n291) );
  AND2X2 U402 ( .A(\mem<13><9> ), .B(n1711), .Y(n292) );
  INVX1 U403 ( .A(n292), .Y(n293) );
  AND2X2 U404 ( .A(\mem<13><10> ), .B(n1711), .Y(n294) );
  INVX1 U405 ( .A(n294), .Y(n295) );
  AND2X2 U406 ( .A(\mem<13><11> ), .B(n1711), .Y(n296) );
  INVX1 U407 ( .A(n296), .Y(n297) );
  AND2X2 U408 ( .A(\mem<13><12> ), .B(n1711), .Y(n298) );
  INVX1 U409 ( .A(n298), .Y(n299) );
  AND2X2 U410 ( .A(\mem<13><13> ), .B(n1711), .Y(n300) );
  INVX1 U411 ( .A(n300), .Y(n301) );
  AND2X2 U412 ( .A(\mem<13><14> ), .B(n1711), .Y(n302) );
  INVX1 U413 ( .A(n302), .Y(n303) );
  AND2X2 U414 ( .A(\mem<13><15> ), .B(n1711), .Y(n304) );
  INVX1 U415 ( .A(n304), .Y(n305) );
  BUFX2 U416 ( .A(n573), .Y(n1711) );
  BUFX2 U417 ( .A(n577), .Y(n1712) );
  AND2X2 U418 ( .A(\mem<12><8> ), .B(n1713), .Y(n306) );
  INVX1 U419 ( .A(n306), .Y(n307) );
  AND2X2 U420 ( .A(\mem<12><9> ), .B(n1713), .Y(n308) );
  INVX1 U421 ( .A(n308), .Y(n309) );
  AND2X2 U422 ( .A(\mem<12><10> ), .B(n1713), .Y(n310) );
  INVX1 U423 ( .A(n310), .Y(n311) );
  AND2X2 U424 ( .A(\mem<12><11> ), .B(n1713), .Y(n312) );
  INVX1 U425 ( .A(n312), .Y(n313) );
  AND2X2 U426 ( .A(\mem<12><12> ), .B(n1713), .Y(n314) );
  INVX1 U427 ( .A(n314), .Y(n315) );
  AND2X2 U428 ( .A(\mem<12><13> ), .B(n1713), .Y(n316) );
  INVX1 U429 ( .A(n316), .Y(n317) );
  AND2X2 U430 ( .A(\mem<12><14> ), .B(n1713), .Y(n318) );
  INVX1 U431 ( .A(n318), .Y(n319) );
  AND2X2 U432 ( .A(\mem<12><15> ), .B(n1713), .Y(n320) );
  INVX1 U433 ( .A(n320), .Y(n321) );
  BUFX2 U434 ( .A(n577), .Y(n1713) );
  BUFX2 U435 ( .A(n581), .Y(n1714) );
  AND2X2 U436 ( .A(\mem<11><8> ), .B(n1715), .Y(n322) );
  INVX1 U437 ( .A(n322), .Y(n323) );
  AND2X2 U438 ( .A(\mem<11><9> ), .B(n1715), .Y(n324) );
  INVX1 U439 ( .A(n324), .Y(n325) );
  AND2X2 U440 ( .A(\mem<11><10> ), .B(n1715), .Y(n326) );
  INVX1 U441 ( .A(n326), .Y(n327) );
  AND2X2 U442 ( .A(\mem<11><11> ), .B(n1715), .Y(n328) );
  INVX1 U443 ( .A(n328), .Y(n329) );
  AND2X2 U444 ( .A(\mem<11><12> ), .B(n1715), .Y(n330) );
  INVX1 U445 ( .A(n330), .Y(n331) );
  AND2X2 U446 ( .A(\mem<11><13> ), .B(n1715), .Y(n332) );
  INVX1 U447 ( .A(n332), .Y(n333) );
  AND2X2 U448 ( .A(\mem<11><14> ), .B(n1715), .Y(n334) );
  INVX1 U449 ( .A(n334), .Y(n335) );
  AND2X2 U450 ( .A(\mem<11><15> ), .B(n1715), .Y(n336) );
  INVX1 U451 ( .A(n336), .Y(n337) );
  BUFX2 U452 ( .A(n581), .Y(n1715) );
  BUFX2 U453 ( .A(n585), .Y(n1716) );
  AND2X2 U454 ( .A(\mem<10><8> ), .B(n1717), .Y(n338) );
  INVX1 U455 ( .A(n338), .Y(n339) );
  AND2X2 U456 ( .A(\mem<10><9> ), .B(n1717), .Y(n340) );
  INVX1 U457 ( .A(n340), .Y(n341) );
  AND2X2 U458 ( .A(\mem<10><10> ), .B(n1717), .Y(n342) );
  INVX1 U459 ( .A(n342), .Y(n343) );
  AND2X2 U460 ( .A(\mem<10><11> ), .B(n1717), .Y(n344) );
  INVX1 U461 ( .A(n344), .Y(n345) );
  AND2X2 U462 ( .A(\mem<10><12> ), .B(n1717), .Y(n346) );
  INVX1 U463 ( .A(n346), .Y(n347) );
  AND2X2 U464 ( .A(\mem<10><13> ), .B(n1717), .Y(n348) );
  INVX1 U465 ( .A(n348), .Y(n349) );
  AND2X2 U466 ( .A(\mem<10><14> ), .B(n1717), .Y(n350) );
  INVX1 U467 ( .A(n350), .Y(n351) );
  AND2X2 U468 ( .A(\mem<10><15> ), .B(n1717), .Y(n352) );
  INVX1 U469 ( .A(n352), .Y(n353) );
  BUFX2 U470 ( .A(n585), .Y(n1717) );
  BUFX2 U471 ( .A(n589), .Y(n1718) );
  AND2X2 U472 ( .A(\mem<9><8> ), .B(n1719), .Y(n354) );
  INVX1 U473 ( .A(n354), .Y(n355) );
  AND2X2 U474 ( .A(\mem<9><9> ), .B(n1719), .Y(n356) );
  INVX1 U475 ( .A(n356), .Y(n357) );
  AND2X2 U476 ( .A(\mem<9><10> ), .B(n1719), .Y(n358) );
  INVX1 U477 ( .A(n358), .Y(n359) );
  AND2X2 U478 ( .A(\mem<9><11> ), .B(n1719), .Y(n360) );
  INVX1 U479 ( .A(n360), .Y(n361) );
  AND2X2 U480 ( .A(\mem<9><12> ), .B(n1719), .Y(n362) );
  INVX1 U481 ( .A(n362), .Y(n363) );
  AND2X2 U482 ( .A(\mem<9><13> ), .B(n1719), .Y(n364) );
  INVX1 U483 ( .A(n364), .Y(n365) );
  AND2X2 U484 ( .A(\mem<9><14> ), .B(n1719), .Y(n366) );
  INVX1 U485 ( .A(n366), .Y(n367) );
  AND2X2 U486 ( .A(\mem<9><15> ), .B(n1719), .Y(n368) );
  INVX1 U487 ( .A(n368), .Y(n369) );
  BUFX2 U488 ( .A(n589), .Y(n1719) );
  BUFX2 U489 ( .A(n591), .Y(n1720) );
  AND2X2 U490 ( .A(\mem<8><11> ), .B(n1721), .Y(n370) );
  INVX1 U491 ( .A(n370), .Y(n371) );
  AND2X2 U492 ( .A(\mem<8><12> ), .B(n1721), .Y(n372) );
  INVX1 U493 ( .A(n372), .Y(n373) );
  AND2X2 U494 ( .A(\mem<8><13> ), .B(n1721), .Y(n374) );
  INVX1 U495 ( .A(n374), .Y(n375) );
  AND2X2 U496 ( .A(\mem<8><14> ), .B(n1721), .Y(n376) );
  INVX1 U497 ( .A(n376), .Y(n377) );
  AND2X2 U498 ( .A(\mem<8><15> ), .B(n1721), .Y(n378) );
  INVX1 U499 ( .A(n378), .Y(n379) );
  BUFX2 U500 ( .A(n591), .Y(n1721) );
  BUFX2 U501 ( .A(n595), .Y(n1722) );
  AND2X2 U502 ( .A(\mem<7><11> ), .B(n1723), .Y(n380) );
  INVX1 U503 ( .A(n380), .Y(n381) );
  AND2X2 U504 ( .A(\mem<7><12> ), .B(n1723), .Y(n382) );
  INVX1 U505 ( .A(n382), .Y(n383) );
  AND2X2 U506 ( .A(\mem<7><13> ), .B(n1723), .Y(n384) );
  INVX1 U507 ( .A(n384), .Y(n385) );
  AND2X2 U508 ( .A(\mem<7><14> ), .B(n1723), .Y(n386) );
  INVX1 U509 ( .A(n386), .Y(n387) );
  AND2X2 U510 ( .A(\mem<7><15> ), .B(n1723), .Y(n388) );
  INVX1 U511 ( .A(n388), .Y(n389) );
  BUFX2 U512 ( .A(n595), .Y(n1723) );
  BUFX2 U513 ( .A(n599), .Y(n1724) );
  AND2X2 U514 ( .A(\mem<6><11> ), .B(n1725), .Y(n390) );
  INVX1 U515 ( .A(n390), .Y(n391) );
  AND2X2 U516 ( .A(\mem<6><12> ), .B(n1725), .Y(n392) );
  INVX1 U517 ( .A(n392), .Y(n393) );
  AND2X2 U518 ( .A(\mem<6><13> ), .B(n1725), .Y(n394) );
  INVX1 U519 ( .A(n394), .Y(n395) );
  AND2X2 U520 ( .A(\mem<6><14> ), .B(n1725), .Y(n396) );
  INVX1 U521 ( .A(n396), .Y(n397) );
  AND2X2 U522 ( .A(\mem<6><15> ), .B(n1725), .Y(n398) );
  INVX1 U523 ( .A(n398), .Y(n399) );
  BUFX2 U524 ( .A(n599), .Y(n1725) );
  BUFX2 U525 ( .A(n603), .Y(n1726) );
  AND2X2 U526 ( .A(\mem<5><11> ), .B(n1727), .Y(n400) );
  INVX1 U527 ( .A(n400), .Y(n401) );
  AND2X2 U528 ( .A(\mem<5><12> ), .B(n1727), .Y(n402) );
  INVX1 U529 ( .A(n402), .Y(n403) );
  AND2X2 U530 ( .A(\mem<5><13> ), .B(n1727), .Y(n404) );
  INVX1 U531 ( .A(n404), .Y(n405) );
  AND2X2 U532 ( .A(\mem<5><14> ), .B(n1727), .Y(n406) );
  INVX1 U533 ( .A(n406), .Y(n407) );
  AND2X2 U534 ( .A(\mem<5><15> ), .B(n1727), .Y(n408) );
  INVX1 U535 ( .A(n408), .Y(n409) );
  BUFX2 U536 ( .A(n603), .Y(n1727) );
  BUFX2 U537 ( .A(n607), .Y(n1728) );
  AND2X2 U538 ( .A(\mem<4><11> ), .B(n1729), .Y(n410) );
  INVX1 U539 ( .A(n410), .Y(n411) );
  AND2X2 U540 ( .A(\mem<4><12> ), .B(n1729), .Y(n412) );
  INVX1 U541 ( .A(n412), .Y(n413) );
  AND2X2 U542 ( .A(\mem<4><13> ), .B(n1729), .Y(n414) );
  INVX1 U543 ( .A(n414), .Y(n415) );
  AND2X2 U544 ( .A(\mem<4><14> ), .B(n1729), .Y(n416) );
  INVX1 U545 ( .A(n416), .Y(n417) );
  AND2X2 U546 ( .A(\mem<4><15> ), .B(n1729), .Y(n418) );
  INVX1 U547 ( .A(n418), .Y(n419) );
  BUFX2 U548 ( .A(n607), .Y(n1729) );
  BUFX2 U549 ( .A(n611), .Y(n1730) );
  AND2X2 U550 ( .A(\mem<3><11> ), .B(n1731), .Y(n420) );
  INVX1 U551 ( .A(n420), .Y(n421) );
  AND2X2 U552 ( .A(\mem<3><12> ), .B(n1731), .Y(n422) );
  INVX1 U553 ( .A(n422), .Y(n423) );
  AND2X2 U554 ( .A(\mem<3><13> ), .B(n1731), .Y(n424) );
  INVX1 U555 ( .A(n424), .Y(n425) );
  AND2X2 U556 ( .A(\mem<3><14> ), .B(n1731), .Y(n426) );
  INVX1 U557 ( .A(n426), .Y(n427) );
  AND2X2 U558 ( .A(\mem<3><15> ), .B(n1731), .Y(n428) );
  INVX1 U559 ( .A(n428), .Y(n429) );
  BUFX2 U560 ( .A(n611), .Y(n1731) );
  BUFX2 U561 ( .A(n615), .Y(n1732) );
  AND2X2 U562 ( .A(\mem<2><11> ), .B(n1733), .Y(n430) );
  INVX1 U563 ( .A(n430), .Y(n431) );
  AND2X2 U564 ( .A(\mem<2><12> ), .B(n1733), .Y(n432) );
  INVX1 U565 ( .A(n432), .Y(n433) );
  AND2X2 U566 ( .A(\mem<2><13> ), .B(n1733), .Y(n434) );
  INVX1 U567 ( .A(n434), .Y(n435) );
  AND2X2 U568 ( .A(\mem<2><14> ), .B(n1733), .Y(n436) );
  INVX1 U569 ( .A(n436), .Y(n437) );
  AND2X2 U570 ( .A(\mem<2><15> ), .B(n1733), .Y(n438) );
  INVX1 U571 ( .A(n438), .Y(n439) );
  BUFX2 U572 ( .A(n615), .Y(n1733) );
  BUFX2 U573 ( .A(n619), .Y(n1734) );
  AND2X2 U574 ( .A(\mem<1><11> ), .B(n1735), .Y(n440) );
  INVX1 U575 ( .A(n440), .Y(n441) );
  AND2X2 U576 ( .A(\mem<1><12> ), .B(n1735), .Y(n442) );
  INVX1 U577 ( .A(n442), .Y(n443) );
  AND2X2 U578 ( .A(\mem<1><13> ), .B(n1735), .Y(n444) );
  INVX1 U579 ( .A(n444), .Y(n445) );
  AND2X2 U580 ( .A(\mem<1><14> ), .B(n1735), .Y(n446) );
  INVX1 U581 ( .A(n446), .Y(n447) );
  AND2X2 U582 ( .A(\mem<1><15> ), .B(n1735), .Y(n448) );
  INVX1 U583 ( .A(n448), .Y(n449) );
  BUFX2 U584 ( .A(n619), .Y(n1735) );
  BUFX2 U585 ( .A(n621), .Y(n1736) );
  AND2X2 U586 ( .A(\mem<0><8> ), .B(n1737), .Y(n450) );
  INVX1 U587 ( .A(n450), .Y(n451) );
  AND2X2 U588 ( .A(\mem<0><9> ), .B(n1737), .Y(n452) );
  INVX1 U589 ( .A(n452), .Y(n453) );
  AND2X2 U590 ( .A(\mem<0><10> ), .B(n1737), .Y(n454) );
  INVX1 U591 ( .A(n454), .Y(n455) );
  AND2X2 U592 ( .A(\mem<0><11> ), .B(n1737), .Y(n456) );
  INVX1 U593 ( .A(n456), .Y(n457) );
  AND2X2 U594 ( .A(\mem<0><12> ), .B(n1737), .Y(n458) );
  INVX1 U595 ( .A(n458), .Y(n459) );
  AND2X2 U596 ( .A(\mem<0><13> ), .B(n1737), .Y(n460) );
  INVX1 U597 ( .A(n460), .Y(n461) );
  AND2X2 U598 ( .A(\mem<0><14> ), .B(n1737), .Y(n462) );
  INVX1 U599 ( .A(n462), .Y(n463) );
  AND2X2 U600 ( .A(\mem<0><15> ), .B(n1737), .Y(n464) );
  INVX1 U601 ( .A(n464), .Y(n465) );
  BUFX2 U602 ( .A(n621), .Y(n1737) );
  INVX1 U603 ( .A(n1769), .Y(n1768) );
  AND2X1 U604 ( .A(n1636), .B(n1765), .Y(n477) );
  INVX1 U605 ( .A(n1766), .Y(n1765) );
  AND2X1 U606 ( .A(n2582), .B(n1770), .Y(n478) );
  INVX1 U607 ( .A(n1771), .Y(n1770) );
  BUFX2 U608 ( .A(n1791), .Y(n479) );
  INVX1 U609 ( .A(n479), .Y(n2000) );
  BUFX2 U610 ( .A(n1800), .Y(n480) );
  INVX1 U611 ( .A(n480), .Y(n2012) );
  BUFX2 U612 ( .A(n1809), .Y(n481) );
  INVX1 U613 ( .A(n481), .Y(n2024) );
  BUFX2 U614 ( .A(n1818), .Y(n482) );
  INVX1 U615 ( .A(n482), .Y(n2036) );
  BUFX2 U616 ( .A(n1827), .Y(n483) );
  INVX1 U617 ( .A(n483), .Y(n2048) );
  BUFX2 U618 ( .A(n1908), .Y(n484) );
  INVX1 U619 ( .A(n484), .Y(n1965) );
  BUFX2 U620 ( .A(n1977), .Y(n485) );
  INVX1 U621 ( .A(n485), .Y(n2060) );
  AND2X1 U622 ( .A(n1667), .B(n477), .Y(n486) );
  AND2X1 U623 ( .A(n1768), .B(n478), .Y(n487) );
  AND2X2 U624 ( .A(write), .B(n1772), .Y(n488) );
  AND2X1 U625 ( .A(n1764), .B(n477), .Y(n489) );
  AND2X1 U626 ( .A(n1769), .B(n478), .Y(n490) );
  AND2X2 U627 ( .A(\data_in<11> ), .B(n1739), .Y(n491) );
  AND2X2 U628 ( .A(\data_in<13> ), .B(n1739), .Y(n493) );
  AND2X2 U629 ( .A(\data_in<15> ), .B(n1739), .Y(n495) );
  AND2X1 U630 ( .A(n487), .B(n2061), .Y(n496) );
  AND2X1 U631 ( .A(n2061), .B(n490), .Y(n497) );
  AND2X1 U632 ( .A(n2061), .B(n1965), .Y(n498) );
  INVX1 U633 ( .A(n498), .Y(n499) );
  AND2X1 U634 ( .A(n2061), .B(n2060), .Y(n500) );
  INVX1 U635 ( .A(n500), .Y(n501) );
  AND2X1 U636 ( .A(n486), .B(n487), .Y(n502) );
  INVX1 U637 ( .A(n502), .Y(n503) );
  AND2X1 U638 ( .A(n1740), .B(n502), .Y(n504) );
  INVX1 U639 ( .A(n504), .Y(n505) );
  AND2X1 U640 ( .A(n487), .B(n489), .Y(n506) );
  INVX1 U641 ( .A(n506), .Y(n507) );
  AND2X1 U642 ( .A(n1738), .B(n506), .Y(n508) );
  INVX1 U643 ( .A(n508), .Y(n509) );
  AND2X1 U644 ( .A(n487), .B(n2000), .Y(n510) );
  INVX1 U645 ( .A(n510), .Y(n511) );
  AND2X1 U646 ( .A(n1740), .B(n510), .Y(n512) );
  INVX1 U647 ( .A(n512), .Y(n513) );
  AND2X1 U648 ( .A(n487), .B(n2012), .Y(n514) );
  INVX1 U649 ( .A(n514), .Y(n515) );
  AND2X1 U650 ( .A(n1738), .B(n514), .Y(n516) );
  INVX1 U651 ( .A(n516), .Y(n517) );
  AND2X1 U652 ( .A(n487), .B(n2024), .Y(n518) );
  INVX1 U653 ( .A(n518), .Y(n519) );
  AND2X1 U654 ( .A(n1740), .B(n518), .Y(n520) );
  INVX1 U655 ( .A(n520), .Y(n521) );
  AND2X1 U656 ( .A(n487), .B(n2036), .Y(n522) );
  INVX1 U657 ( .A(n522), .Y(n523) );
  AND2X1 U658 ( .A(n1738), .B(n522), .Y(n524) );
  INVX1 U659 ( .A(n524), .Y(n525) );
  AND2X1 U660 ( .A(n487), .B(n2048), .Y(n526) );
  INVX1 U661 ( .A(n526), .Y(n527) );
  AND2X1 U662 ( .A(n1740), .B(n526), .Y(n528) );
  INVX1 U663 ( .A(n528), .Y(n529) );
  AND2X1 U664 ( .A(n1738), .B(n496), .Y(n530) );
  INVX1 U665 ( .A(n530), .Y(n531) );
  AND2X1 U666 ( .A(n486), .B(n490), .Y(n532) );
  INVX1 U667 ( .A(n532), .Y(n533) );
  AND2X1 U668 ( .A(n1738), .B(n532), .Y(n534) );
  INVX1 U669 ( .A(n534), .Y(n535) );
  AND2X1 U670 ( .A(n489), .B(n490), .Y(n536) );
  INVX1 U671 ( .A(n536), .Y(n537) );
  AND2X1 U672 ( .A(n1740), .B(n536), .Y(n538) );
  INVX1 U673 ( .A(n538), .Y(n539) );
  AND2X1 U674 ( .A(n2000), .B(n490), .Y(n540) );
  INVX1 U675 ( .A(n540), .Y(n541) );
  AND2X1 U676 ( .A(n1738), .B(n540), .Y(n542) );
  INVX1 U677 ( .A(n542), .Y(n543) );
  AND2X1 U678 ( .A(n2012), .B(n490), .Y(n544) );
  INVX1 U679 ( .A(n544), .Y(n545) );
  AND2X1 U680 ( .A(n1740), .B(n544), .Y(n546) );
  INVX1 U681 ( .A(n546), .Y(n547) );
  AND2X1 U682 ( .A(n2024), .B(n490), .Y(n548) );
  INVX1 U683 ( .A(n548), .Y(n549) );
  AND2X1 U684 ( .A(n1738), .B(n548), .Y(n550) );
  INVX1 U685 ( .A(n550), .Y(n551) );
  AND2X1 U686 ( .A(n2036), .B(n490), .Y(n552) );
  INVX1 U687 ( .A(n552), .Y(n553) );
  AND2X1 U688 ( .A(n1738), .B(n552), .Y(n554) );
  INVX1 U689 ( .A(n554), .Y(n555) );
  AND2X1 U690 ( .A(n2048), .B(n490), .Y(n556) );
  INVX1 U691 ( .A(n556), .Y(n557) );
  AND2X1 U692 ( .A(n1738), .B(n556), .Y(n558) );
  INVX1 U693 ( .A(n558), .Y(n559) );
  AND2X1 U694 ( .A(n1738), .B(n497), .Y(n560) );
  INVX1 U695 ( .A(n560), .Y(n561) );
  AND2X1 U696 ( .A(n486), .B(n1965), .Y(n562) );
  INVX1 U697 ( .A(n562), .Y(n563) );
  AND2X1 U698 ( .A(n1738), .B(n562), .Y(n564) );
  INVX1 U699 ( .A(n564), .Y(n565) );
  AND2X1 U700 ( .A(n489), .B(n1965), .Y(n566) );
  INVX1 U701 ( .A(n566), .Y(n567) );
  AND2X1 U702 ( .A(n1738), .B(n566), .Y(n568) );
  INVX1 U703 ( .A(n568), .Y(n569) );
  AND2X1 U704 ( .A(n2000), .B(n1965), .Y(n570) );
  INVX1 U705 ( .A(n570), .Y(n571) );
  AND2X1 U706 ( .A(n1738), .B(n570), .Y(n572) );
  INVX1 U707 ( .A(n572), .Y(n573) );
  AND2X1 U708 ( .A(n2012), .B(n1965), .Y(n574) );
  INVX1 U709 ( .A(n574), .Y(n575) );
  AND2X1 U710 ( .A(n1738), .B(n574), .Y(n576) );
  INVX1 U711 ( .A(n576), .Y(n577) );
  AND2X1 U712 ( .A(n2024), .B(n1965), .Y(n578) );
  INVX1 U713 ( .A(n578), .Y(n579) );
  AND2X1 U714 ( .A(n1738), .B(n578), .Y(n580) );
  INVX1 U715 ( .A(n580), .Y(n581) );
  AND2X1 U716 ( .A(n2036), .B(n1965), .Y(n582) );
  INVX1 U717 ( .A(n582), .Y(n583) );
  AND2X1 U718 ( .A(n1738), .B(n582), .Y(n584) );
  INVX1 U719 ( .A(n584), .Y(n585) );
  AND2X1 U720 ( .A(n2048), .B(n1965), .Y(n586) );
  INVX1 U721 ( .A(n586), .Y(n587) );
  AND2X1 U722 ( .A(n1738), .B(n586), .Y(n588) );
  INVX1 U723 ( .A(n588), .Y(n589) );
  AND2X1 U724 ( .A(n1739), .B(n498), .Y(n590) );
  INVX1 U725 ( .A(n590), .Y(n591) );
  AND2X1 U726 ( .A(n486), .B(n2060), .Y(n592) );
  INVX1 U727 ( .A(n592), .Y(n593) );
  AND2X1 U728 ( .A(n1739), .B(n592), .Y(n594) );
  INVX1 U729 ( .A(n594), .Y(n595) );
  AND2X1 U730 ( .A(n489), .B(n2060), .Y(n596) );
  INVX1 U731 ( .A(n596), .Y(n597) );
  AND2X1 U732 ( .A(n1739), .B(n596), .Y(n598) );
  INVX1 U733 ( .A(n598), .Y(n599) );
  AND2X1 U734 ( .A(n2000), .B(n2060), .Y(n600) );
  INVX1 U735 ( .A(n600), .Y(n601) );
  AND2X1 U736 ( .A(n1739), .B(n600), .Y(n602) );
  INVX1 U737 ( .A(n602), .Y(n603) );
  AND2X1 U738 ( .A(n2012), .B(n2060), .Y(n604) );
  INVX1 U739 ( .A(n604), .Y(n605) );
  AND2X1 U740 ( .A(n1739), .B(n604), .Y(n606) );
  INVX1 U741 ( .A(n606), .Y(n607) );
  AND2X1 U742 ( .A(n2024), .B(n2060), .Y(n608) );
  INVX1 U743 ( .A(n608), .Y(n609) );
  AND2X1 U744 ( .A(n1739), .B(n608), .Y(n610) );
  INVX1 U745 ( .A(n610), .Y(n611) );
  AND2X1 U746 ( .A(n2036), .B(n2060), .Y(n612) );
  INVX1 U747 ( .A(n612), .Y(n613) );
  AND2X1 U748 ( .A(n1739), .B(n612), .Y(n614) );
  INVX1 U749 ( .A(n614), .Y(n615) );
  AND2X1 U750 ( .A(n2048), .B(n2060), .Y(n616) );
  INVX1 U751 ( .A(n616), .Y(n617) );
  AND2X1 U752 ( .A(n1739), .B(n616), .Y(n618) );
  INVX1 U753 ( .A(n618), .Y(n619) );
  AND2X1 U754 ( .A(n1738), .B(n500), .Y(n620) );
  INVX1 U755 ( .A(n620), .Y(n621) );
  MUX2X1 U756 ( .B(n623), .A(n624), .S(n1640), .Y(n622) );
  MUX2X1 U757 ( .B(n626), .A(n627), .S(n1640), .Y(n625) );
  MUX2X1 U758 ( .B(n629), .A(n630), .S(n1640), .Y(n628) );
  MUX2X1 U759 ( .B(n632), .A(n633), .S(n1640), .Y(n631) );
  MUX2X1 U760 ( .B(n635), .A(n636), .S(n1633), .Y(n634) );
  MUX2X1 U761 ( .B(n638), .A(n639), .S(n1640), .Y(n637) );
  MUX2X1 U762 ( .B(n641), .A(n642), .S(n1640), .Y(n640) );
  MUX2X1 U763 ( .B(n644), .A(n645), .S(n1640), .Y(n643) );
  MUX2X1 U764 ( .B(n647), .A(n648), .S(n1640), .Y(n646) );
  MUX2X1 U765 ( .B(n650), .A(n1163), .S(n1633), .Y(n649) );
  MUX2X1 U766 ( .B(n1165), .A(n1166), .S(n1641), .Y(n1164) );
  MUX2X1 U767 ( .B(n1168), .A(n1169), .S(n1641), .Y(n1167) );
  MUX2X1 U768 ( .B(n1171), .A(n1172), .S(n1641), .Y(n1170) );
  MUX2X1 U769 ( .B(n1174), .A(n1175), .S(n1641), .Y(n1173) );
  MUX2X1 U770 ( .B(n1177), .A(n1178), .S(n1633), .Y(n1176) );
  MUX2X1 U771 ( .B(n1180), .A(n1181), .S(n1641), .Y(n1179) );
  MUX2X1 U772 ( .B(n1183), .A(n1184), .S(n1641), .Y(n1182) );
  MUX2X1 U773 ( .B(n1186), .A(n1187), .S(n1641), .Y(n1185) );
  MUX2X1 U774 ( .B(n1189), .A(n1190), .S(n1641), .Y(n1188) );
  MUX2X1 U775 ( .B(n1192), .A(n1193), .S(n1633), .Y(n1191) );
  MUX2X1 U776 ( .B(n1195), .A(n1196), .S(n1641), .Y(n1194) );
  MUX2X1 U777 ( .B(n1198), .A(n1199), .S(n1641), .Y(n1197) );
  MUX2X1 U778 ( .B(n1201), .A(n1202), .S(n1641), .Y(n1200) );
  MUX2X1 U779 ( .B(n1204), .A(n1205), .S(n1641), .Y(n1203) );
  MUX2X1 U780 ( .B(n1207), .A(n1208), .S(n1633), .Y(n1206) );
  MUX2X1 U781 ( .B(n1210), .A(n1211), .S(n1642), .Y(n1209) );
  MUX2X1 U782 ( .B(n1213), .A(n1214), .S(n1642), .Y(n1212) );
  MUX2X1 U783 ( .B(n1216), .A(n1217), .S(n1642), .Y(n1215) );
  MUX2X1 U784 ( .B(n1219), .A(n1220), .S(n1642), .Y(n1218) );
  MUX2X1 U785 ( .B(n1222), .A(n1223), .S(n1633), .Y(n1221) );
  MUX2X1 U786 ( .B(n1225), .A(n1226), .S(n1642), .Y(n1224) );
  MUX2X1 U787 ( .B(n1228), .A(n1229), .S(n1642), .Y(n1227) );
  MUX2X1 U788 ( .B(n1231), .A(n1232), .S(n1642), .Y(n1230) );
  MUX2X1 U789 ( .B(n1234), .A(n1235), .S(n1642), .Y(n1233) );
  MUX2X1 U790 ( .B(n1237), .A(n1238), .S(n1633), .Y(n1236) );
  MUX2X1 U791 ( .B(n1240), .A(n1241), .S(n1642), .Y(n1239) );
  MUX2X1 U792 ( .B(n1243), .A(n1244), .S(n1642), .Y(n1242) );
  MUX2X1 U793 ( .B(n1246), .A(n1247), .S(n1642), .Y(n1245) );
  MUX2X1 U794 ( .B(n1249), .A(n1250), .S(n1642), .Y(n1248) );
  MUX2X1 U795 ( .B(n1252), .A(n1253), .S(n1633), .Y(n1251) );
  MUX2X1 U796 ( .B(n1255), .A(n1256), .S(n1643), .Y(n1254) );
  MUX2X1 U797 ( .B(n1258), .A(n1259), .S(n1643), .Y(n1257) );
  MUX2X1 U798 ( .B(n1261), .A(n1262), .S(n1643), .Y(n1260) );
  MUX2X1 U799 ( .B(n1264), .A(n1265), .S(n1643), .Y(n1263) );
  MUX2X1 U800 ( .B(n1267), .A(n1268), .S(n1633), .Y(n1266) );
  MUX2X1 U801 ( .B(n1270), .A(n1271), .S(n1643), .Y(n1269) );
  MUX2X1 U802 ( .B(n1273), .A(n1274), .S(n1643), .Y(n1272) );
  MUX2X1 U803 ( .B(n1276), .A(n1277), .S(n1643), .Y(n1275) );
  MUX2X1 U804 ( .B(n1279), .A(n1280), .S(n1643), .Y(n1278) );
  MUX2X1 U805 ( .B(n1282), .A(n1283), .S(n1633), .Y(n1281) );
  MUX2X1 U806 ( .B(n1285), .A(n1286), .S(n1643), .Y(n1284) );
  MUX2X1 U807 ( .B(n1288), .A(n1289), .S(n1643), .Y(n1287) );
  MUX2X1 U808 ( .B(n1291), .A(n1292), .S(n1643), .Y(n1290) );
  MUX2X1 U809 ( .B(n1294), .A(n1295), .S(n1643), .Y(n1293) );
  MUX2X1 U810 ( .B(n1297), .A(n1298), .S(n1633), .Y(n1296) );
  MUX2X1 U811 ( .B(n1300), .A(n1301), .S(n1644), .Y(n1299) );
  MUX2X1 U812 ( .B(n1303), .A(n1304), .S(n1644), .Y(n1302) );
  MUX2X1 U813 ( .B(n1306), .A(n1307), .S(n1644), .Y(n1305) );
  MUX2X1 U814 ( .B(n1309), .A(n1310), .S(n1644), .Y(n1308) );
  MUX2X1 U815 ( .B(n1312), .A(n1313), .S(n1633), .Y(n1311) );
  MUX2X1 U816 ( .B(n1315), .A(n1316), .S(n1644), .Y(n1314) );
  MUX2X1 U817 ( .B(n1318), .A(n1319), .S(n1644), .Y(n1317) );
  MUX2X1 U818 ( .B(n1321), .A(n1322), .S(n1644), .Y(n1320) );
  MUX2X1 U819 ( .B(n1324), .A(n1325), .S(n1644), .Y(n1323) );
  MUX2X1 U820 ( .B(n1327), .A(n1328), .S(n1632), .Y(n1326) );
  MUX2X1 U821 ( .B(n1330), .A(n1331), .S(n1644), .Y(n1329) );
  MUX2X1 U822 ( .B(n1333), .A(n1334), .S(n1644), .Y(n1332) );
  MUX2X1 U823 ( .B(n1336), .A(n1337), .S(n1644), .Y(n1335) );
  MUX2X1 U824 ( .B(n1339), .A(n1340), .S(n1644), .Y(n1338) );
  MUX2X1 U825 ( .B(n1342), .A(n1343), .S(n1632), .Y(n1341) );
  MUX2X1 U826 ( .B(n1345), .A(n1346), .S(n1645), .Y(n1344) );
  MUX2X1 U827 ( .B(n1348), .A(n1349), .S(n1645), .Y(n1347) );
  MUX2X1 U828 ( .B(n1351), .A(n1352), .S(n1645), .Y(n1350) );
  MUX2X1 U829 ( .B(n1354), .A(n1355), .S(n1645), .Y(n1353) );
  MUX2X1 U830 ( .B(n1357), .A(n1358), .S(n1632), .Y(n1356) );
  MUX2X1 U831 ( .B(n1360), .A(n1361), .S(n1645), .Y(n1359) );
  MUX2X1 U832 ( .B(n1363), .A(n1364), .S(n1645), .Y(n1362) );
  MUX2X1 U833 ( .B(n1366), .A(n1367), .S(n1645), .Y(n1365) );
  MUX2X1 U834 ( .B(n1369), .A(n1370), .S(n1645), .Y(n1368) );
  MUX2X1 U835 ( .B(n1372), .A(n1373), .S(n1632), .Y(n1371) );
  MUX2X1 U836 ( .B(n1375), .A(n1376), .S(n1645), .Y(n1374) );
  MUX2X1 U837 ( .B(n1378), .A(n1379), .S(n1645), .Y(n1377) );
  MUX2X1 U838 ( .B(n1381), .A(n1382), .S(n1645), .Y(n1380) );
  MUX2X1 U839 ( .B(n1384), .A(n1385), .S(n1645), .Y(n1383) );
  MUX2X1 U840 ( .B(n1387), .A(n1388), .S(n1632), .Y(n1386) );
  MUX2X1 U841 ( .B(n1390), .A(n1391), .S(n1646), .Y(n1389) );
  MUX2X1 U842 ( .B(n1393), .A(n1394), .S(n1646), .Y(n1392) );
  MUX2X1 U843 ( .B(n1396), .A(n1397), .S(n1646), .Y(n1395) );
  MUX2X1 U844 ( .B(n1399), .A(n1400), .S(n1646), .Y(n1398) );
  MUX2X1 U845 ( .B(n1402), .A(n1403), .S(n1632), .Y(n1401) );
  MUX2X1 U846 ( .B(n1405), .A(n1406), .S(n1646), .Y(n1404) );
  MUX2X1 U847 ( .B(n1408), .A(n1409), .S(n1646), .Y(n1407) );
  MUX2X1 U848 ( .B(n1411), .A(n1412), .S(n1646), .Y(n1410) );
  MUX2X1 U849 ( .B(n1414), .A(n1415), .S(n1646), .Y(n1413) );
  MUX2X1 U850 ( .B(n1417), .A(n1418), .S(n1632), .Y(n1416) );
  MUX2X1 U851 ( .B(n1420), .A(n1421), .S(n1646), .Y(n1419) );
  MUX2X1 U852 ( .B(n1423), .A(n1424), .S(n1646), .Y(n1422) );
  MUX2X1 U853 ( .B(n1426), .A(n1427), .S(n1646), .Y(n1425) );
  MUX2X1 U854 ( .B(n1429), .A(n1430), .S(n1646), .Y(n1428) );
  MUX2X1 U855 ( .B(n1432), .A(n1433), .S(n1632), .Y(n1431) );
  MUX2X1 U856 ( .B(n1435), .A(n1436), .S(n1647), .Y(n1434) );
  MUX2X1 U857 ( .B(n1438), .A(n1439), .S(n1647), .Y(n1437) );
  MUX2X1 U858 ( .B(n1441), .A(n1442), .S(n1647), .Y(n1440) );
  MUX2X1 U859 ( .B(n1444), .A(n1445), .S(n1647), .Y(n1443) );
  MUX2X1 U860 ( .B(n1447), .A(n1448), .S(n1632), .Y(n1446) );
  MUX2X1 U861 ( .B(n1450), .A(n1451), .S(n1647), .Y(n1449) );
  MUX2X1 U862 ( .B(n1453), .A(n1454), .S(n1647), .Y(n1452) );
  MUX2X1 U863 ( .B(n1456), .A(n1457), .S(n1647), .Y(n1455) );
  MUX2X1 U864 ( .B(n1459), .A(n1460), .S(n1647), .Y(n1458) );
  MUX2X1 U865 ( .B(n1462), .A(n1463), .S(n1632), .Y(n1461) );
  MUX2X1 U866 ( .B(n1465), .A(n1466), .S(n1647), .Y(n1464) );
  MUX2X1 U867 ( .B(n1468), .A(n1469), .S(n1647), .Y(n1467) );
  MUX2X1 U868 ( .B(n1471), .A(n1472), .S(n1647), .Y(n1470) );
  MUX2X1 U869 ( .B(n1474), .A(n1475), .S(n1647), .Y(n1473) );
  MUX2X1 U870 ( .B(n1477), .A(n1478), .S(n1632), .Y(n1476) );
  MUX2X1 U871 ( .B(n1480), .A(n1481), .S(n1648), .Y(n1479) );
  MUX2X1 U872 ( .B(n1483), .A(n1484), .S(n1648), .Y(n1482) );
  MUX2X1 U873 ( .B(n1486), .A(n1487), .S(n1648), .Y(n1485) );
  MUX2X1 U874 ( .B(n1489), .A(n1490), .S(n1648), .Y(n1488) );
  MUX2X1 U875 ( .B(n1492), .A(n1493), .S(n1632), .Y(n1491) );
  MUX2X1 U876 ( .B(n1495), .A(n1496), .S(n1648), .Y(n1494) );
  MUX2X1 U877 ( .B(n1498), .A(n1499), .S(n1648), .Y(n1497) );
  MUX2X1 U878 ( .B(n1501), .A(n1502), .S(n1648), .Y(n1500) );
  MUX2X1 U879 ( .B(n1504), .A(n1505), .S(n1648), .Y(n1503) );
  MUX2X1 U880 ( .B(n1507), .A(n1508), .S(n1631), .Y(n1506) );
  MUX2X1 U881 ( .B(n1510), .A(n1511), .S(n1648), .Y(n1509) );
  MUX2X1 U882 ( .B(n1513), .A(n1514), .S(n1648), .Y(n1512) );
  MUX2X1 U883 ( .B(n1516), .A(n1517), .S(n1648), .Y(n1515) );
  MUX2X1 U884 ( .B(n1519), .A(n1520), .S(n1648), .Y(n1518) );
  MUX2X1 U885 ( .B(n1522), .A(n1523), .S(n1631), .Y(n1521) );
  MUX2X1 U886 ( .B(n1525), .A(n1526), .S(n1649), .Y(n1524) );
  MUX2X1 U887 ( .B(n1528), .A(n1529), .S(n1649), .Y(n1527) );
  MUX2X1 U888 ( .B(n1531), .A(n1532), .S(n1649), .Y(n1530) );
  MUX2X1 U889 ( .B(n1534), .A(n1535), .S(n1649), .Y(n1533) );
  MUX2X1 U890 ( .B(n1537), .A(n1538), .S(n1631), .Y(n1536) );
  MUX2X1 U891 ( .B(n1540), .A(n1541), .S(n1649), .Y(n1539) );
  MUX2X1 U892 ( .B(n1543), .A(n1544), .S(n1649), .Y(n1542) );
  MUX2X1 U893 ( .B(n1546), .A(n1547), .S(n1649), .Y(n1545) );
  MUX2X1 U894 ( .B(n1549), .A(n1550), .S(n1649), .Y(n1548) );
  MUX2X1 U895 ( .B(n1552), .A(n1553), .S(n1631), .Y(n1551) );
  MUX2X1 U896 ( .B(n1555), .A(n1556), .S(n1649), .Y(n1554) );
  MUX2X1 U897 ( .B(n1558), .A(n1559), .S(n1649), .Y(n1557) );
  MUX2X1 U898 ( .B(n1561), .A(n1562), .S(n1649), .Y(n1560) );
  MUX2X1 U899 ( .B(n1564), .A(n1565), .S(n1649), .Y(n1563) );
  MUX2X1 U900 ( .B(n1567), .A(n1568), .S(n1631), .Y(n1566) );
  MUX2X1 U901 ( .B(n1570), .A(n1571), .S(n1650), .Y(n1569) );
  MUX2X1 U902 ( .B(n1573), .A(n1574), .S(n1650), .Y(n1572) );
  MUX2X1 U903 ( .B(n1576), .A(n1577), .S(n1650), .Y(n1575) );
  MUX2X1 U904 ( .B(n1579), .A(n1580), .S(n1650), .Y(n1578) );
  MUX2X1 U905 ( .B(n1582), .A(n1583), .S(n1631), .Y(n1581) );
  MUX2X1 U906 ( .B(n1585), .A(n1586), .S(n1650), .Y(n1584) );
  MUX2X1 U907 ( .B(n1588), .A(n1589), .S(n1650), .Y(n1587) );
  MUX2X1 U908 ( .B(n1591), .A(n1592), .S(n1650), .Y(n1590) );
  MUX2X1 U909 ( .B(n1594), .A(n1595), .S(n1650), .Y(n1593) );
  MUX2X1 U910 ( .B(n1597), .A(n1598), .S(n1631), .Y(n1596) );
  MUX2X1 U911 ( .B(n1600), .A(n1601), .S(n1650), .Y(n1599) );
  MUX2X1 U912 ( .B(n1603), .A(n1604), .S(n1650), .Y(n1602) );
  MUX2X1 U913 ( .B(n1606), .A(n1607), .S(n1650), .Y(n1605) );
  MUX2X1 U914 ( .B(n1609), .A(n1610), .S(n1650), .Y(n1608) );
  MUX2X1 U915 ( .B(n1612), .A(n1613), .S(n1631), .Y(n1611) );
  MUX2X1 U916 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1663), .Y(n624) );
  MUX2X1 U917 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1662), .Y(n623) );
  MUX2X1 U918 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1658), .Y(n627) );
  MUX2X1 U919 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1657), .Y(n626) );
  MUX2X1 U920 ( .B(n625), .A(n622), .S(n1637), .Y(n636) );
  MUX2X1 U921 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1655), .Y(n630) );
  MUX2X1 U922 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1655), .Y(n629) );
  MUX2X1 U923 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1655), .Y(n633) );
  MUX2X1 U924 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1655), .Y(n632) );
  MUX2X1 U925 ( .B(n631), .A(n628), .S(n1637), .Y(n635) );
  MUX2X1 U926 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1655), .Y(n639) );
  MUX2X1 U927 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1655), .Y(n638) );
  MUX2X1 U928 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1655), .Y(n642) );
  MUX2X1 U929 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1655), .Y(n641) );
  MUX2X1 U930 ( .B(n640), .A(n637), .S(n1637), .Y(n1163) );
  MUX2X1 U931 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1655), .Y(n645) );
  MUX2X1 U932 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1655), .Y(n644) );
  MUX2X1 U933 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1655), .Y(n648) );
  MUX2X1 U934 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1655), .Y(n647) );
  MUX2X1 U935 ( .B(n646), .A(n643), .S(n1637), .Y(n650) );
  MUX2X1 U936 ( .B(n649), .A(n634), .S(n1630), .Y(n1614) );
  MUX2X1 U937 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1656), .Y(n1166) );
  MUX2X1 U938 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1656), .Y(n1165) );
  MUX2X1 U939 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1656), .Y(n1169) );
  MUX2X1 U940 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1656), .Y(n1168) );
  MUX2X1 U941 ( .B(n1167), .A(n1164), .S(n1637), .Y(n1178) );
  MUX2X1 U942 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1656), .Y(n1172) );
  MUX2X1 U943 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1656), .Y(n1171) );
  MUX2X1 U944 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1656), .Y(n1175) );
  MUX2X1 U945 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1656), .Y(n1174) );
  MUX2X1 U946 ( .B(n1173), .A(n1170), .S(n1637), .Y(n1177) );
  MUX2X1 U947 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1656), .Y(n1181) );
  MUX2X1 U948 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1656), .Y(n1180) );
  MUX2X1 U949 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1656), .Y(n1184) );
  MUX2X1 U950 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1656), .Y(n1183) );
  MUX2X1 U951 ( .B(n1182), .A(n1179), .S(n1637), .Y(n1193) );
  MUX2X1 U952 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1657), .Y(n1187) );
  MUX2X1 U953 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1657), .Y(n1186) );
  MUX2X1 U954 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1657), .Y(n1190) );
  MUX2X1 U955 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1657), .Y(n1189) );
  MUX2X1 U956 ( .B(n1188), .A(n1185), .S(n1637), .Y(n1192) );
  MUX2X1 U957 ( .B(n1191), .A(n1176), .S(n1630), .Y(n1615) );
  MUX2X1 U958 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1657), .Y(n1196) );
  MUX2X1 U959 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1657), .Y(n1195) );
  MUX2X1 U960 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1657), .Y(n1199) );
  MUX2X1 U961 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1657), .Y(n1198) );
  MUX2X1 U962 ( .B(n1197), .A(n1194), .S(n1637), .Y(n1208) );
  MUX2X1 U963 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1657), .Y(n1202) );
  MUX2X1 U964 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1657), .Y(n1201) );
  MUX2X1 U965 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1657), .Y(n1205) );
  MUX2X1 U966 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1657), .Y(n1204) );
  MUX2X1 U967 ( .B(n1203), .A(n1200), .S(n1637), .Y(n1207) );
  MUX2X1 U968 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1658), .Y(n1211) );
  MUX2X1 U969 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1658), .Y(n1210) );
  MUX2X1 U970 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1658), .Y(n1214) );
  MUX2X1 U971 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1658), .Y(n1213) );
  MUX2X1 U972 ( .B(n1212), .A(n1209), .S(n1637), .Y(n1223) );
  MUX2X1 U973 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1658), .Y(n1217) );
  MUX2X1 U974 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1658), .Y(n1216) );
  MUX2X1 U975 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1658), .Y(n1220) );
  MUX2X1 U976 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1658), .Y(n1219) );
  MUX2X1 U977 ( .B(n1218), .A(n1215), .S(n1637), .Y(n1222) );
  MUX2X1 U978 ( .B(n1221), .A(n1206), .S(n1630), .Y(n1616) );
  MUX2X1 U979 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1658), .Y(n1226) );
  MUX2X1 U980 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1658), .Y(n1225) );
  MUX2X1 U981 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1658), .Y(n1229) );
  MUX2X1 U982 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1658), .Y(n1228) );
  MUX2X1 U983 ( .B(n1227), .A(n1224), .S(n1636), .Y(n1238) );
  MUX2X1 U984 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1658), .Y(n1232) );
  MUX2X1 U985 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1657), .Y(n1231) );
  MUX2X1 U986 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1670), .Y(n1235) );
  MUX2X1 U987 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1670), .Y(n1234) );
  MUX2X1 U988 ( .B(n1233), .A(n1230), .S(n1636), .Y(n1237) );
  MUX2X1 U989 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1669), .Y(n1241) );
  MUX2X1 U990 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1663), .Y(n1240) );
  MUX2X1 U991 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1670), .Y(n1244) );
  MUX2X1 U992 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1669), .Y(n1243) );
  MUX2X1 U993 ( .B(n1242), .A(n1239), .S(n1636), .Y(n1253) );
  MUX2X1 U994 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1669), .Y(n1247) );
  MUX2X1 U995 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1658), .Y(n1246) );
  MUX2X1 U996 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1657), .Y(n1250) );
  MUX2X1 U997 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1670), .Y(n1249) );
  MUX2X1 U998 ( .B(n1248), .A(n1245), .S(n1636), .Y(n1252) );
  MUX2X1 U999 ( .B(n1251), .A(n1236), .S(n1630), .Y(n1617) );
  MUX2X1 U1000 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1659), .Y(n1256) );
  MUX2X1 U1001 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1659), .Y(n1255) );
  MUX2X1 U1002 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1659), .Y(n1259) );
  MUX2X1 U1003 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1659), .Y(n1258) );
  MUX2X1 U1004 ( .B(n1257), .A(n1254), .S(n1636), .Y(n1268) );
  MUX2X1 U1005 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1659), .Y(n1262) );
  MUX2X1 U1006 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1659), .Y(n1261) );
  MUX2X1 U1007 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1659), .Y(n1265) );
  MUX2X1 U1008 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1659), .Y(n1264) );
  MUX2X1 U1009 ( .B(n1263), .A(n1260), .S(n1636), .Y(n1267) );
  MUX2X1 U1010 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1659), .Y(n1271) );
  MUX2X1 U1011 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1659), .Y(n1270) );
  MUX2X1 U1012 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1659), .Y(n1274) );
  MUX2X1 U1013 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1659), .Y(n1273) );
  MUX2X1 U1014 ( .B(n1272), .A(n1269), .S(n1636), .Y(n1283) );
  MUX2X1 U1015 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1660), .Y(n1277) );
  MUX2X1 U1016 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1660), .Y(n1276) );
  MUX2X1 U1017 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1660), .Y(n1280) );
  MUX2X1 U1018 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1660), .Y(n1279) );
  MUX2X1 U1019 ( .B(n1278), .A(n1275), .S(n1636), .Y(n1282) );
  MUX2X1 U1020 ( .B(n1281), .A(n1266), .S(n1630), .Y(n1618) );
  MUX2X1 U1021 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1660), .Y(n1286) );
  MUX2X1 U1022 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1660), .Y(n1285) );
  MUX2X1 U1023 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1660), .Y(n1289) );
  MUX2X1 U1024 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1660), .Y(n1288) );
  MUX2X1 U1025 ( .B(n1287), .A(n1284), .S(n1636), .Y(n1298) );
  MUX2X1 U1026 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1660), .Y(n1292) );
  MUX2X1 U1027 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1660), .Y(n1291) );
  MUX2X1 U1028 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1660), .Y(n1295) );
  MUX2X1 U1029 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1660), .Y(n1294) );
  MUX2X1 U1030 ( .B(n1293), .A(n1290), .S(n1636), .Y(n1297) );
  MUX2X1 U1031 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1661), .Y(n1301) );
  MUX2X1 U1032 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1661), .Y(n1300) );
  MUX2X1 U1033 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1661), .Y(n1304) );
  MUX2X1 U1034 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1661), .Y(n1303) );
  MUX2X1 U1035 ( .B(n1302), .A(n1299), .S(n1636), .Y(n1313) );
  MUX2X1 U1036 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1661), .Y(n1307) );
  MUX2X1 U1037 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1661), .Y(n1306) );
  MUX2X1 U1038 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1661), .Y(n1310) );
  MUX2X1 U1039 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1661), .Y(n1309) );
  MUX2X1 U1040 ( .B(n1308), .A(n1305), .S(n1636), .Y(n1312) );
  MUX2X1 U1041 ( .B(n1311), .A(n1296), .S(n1630), .Y(n1619) );
  MUX2X1 U1042 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1661), .Y(n1316) );
  MUX2X1 U1043 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1661), .Y(n1315) );
  MUX2X1 U1044 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1661), .Y(n1319) );
  MUX2X1 U1045 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1661), .Y(n1318) );
  MUX2X1 U1046 ( .B(n1317), .A(n1314), .S(n1635), .Y(n1328) );
  MUX2X1 U1047 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1661), .Y(n1322) );
  MUX2X1 U1048 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1661), .Y(n1321) );
  MUX2X1 U1049 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1661), .Y(n1325) );
  MUX2X1 U1050 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1661), .Y(n1324) );
  MUX2X1 U1051 ( .B(n1323), .A(n1320), .S(n1635), .Y(n1327) );
  MUX2X1 U1052 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1661), .Y(n1331) );
  MUX2X1 U1053 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1661), .Y(n1330) );
  MUX2X1 U1054 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1661), .Y(n1334) );
  MUX2X1 U1055 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1661), .Y(n1333) );
  MUX2X1 U1056 ( .B(n1332), .A(n1329), .S(n1635), .Y(n1343) );
  MUX2X1 U1057 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1661), .Y(n1337) );
  MUX2X1 U1058 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1661), .Y(n1336) );
  MUX2X1 U1059 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1661), .Y(n1340) );
  MUX2X1 U1060 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1661), .Y(n1339) );
  MUX2X1 U1061 ( .B(n1338), .A(n1335), .S(n1635), .Y(n1342) );
  MUX2X1 U1062 ( .B(n1341), .A(n1326), .S(n1630), .Y(n1620) );
  MUX2X1 U1063 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1662), .Y(n1346) );
  MUX2X1 U1064 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1662), .Y(n1345) );
  MUX2X1 U1065 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1662), .Y(n1349) );
  MUX2X1 U1066 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1662), .Y(n1348) );
  MUX2X1 U1067 ( .B(n1347), .A(n1344), .S(n1635), .Y(n1358) );
  MUX2X1 U1068 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1662), .Y(n1352) );
  MUX2X1 U1069 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1662), .Y(n1351) );
  MUX2X1 U1070 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1662), .Y(n1355) );
  MUX2X1 U1071 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1662), .Y(n1354) );
  MUX2X1 U1072 ( .B(n1353), .A(n1350), .S(n1635), .Y(n1357) );
  MUX2X1 U1073 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1662), .Y(n1361) );
  MUX2X1 U1074 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1662), .Y(n1360) );
  MUX2X1 U1075 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1662), .Y(n1364) );
  MUX2X1 U1076 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1662), .Y(n1363) );
  MUX2X1 U1077 ( .B(n1362), .A(n1359), .S(n1635), .Y(n1373) );
  MUX2X1 U1078 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1663), .Y(n1367) );
  MUX2X1 U1079 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1663), .Y(n1366) );
  MUX2X1 U1080 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1663), .Y(n1370) );
  MUX2X1 U1081 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1663), .Y(n1369) );
  MUX2X1 U1082 ( .B(n1368), .A(n1365), .S(n1635), .Y(n1372) );
  MUX2X1 U1083 ( .B(n1371), .A(n1356), .S(n1630), .Y(n1621) );
  MUX2X1 U1084 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1663), .Y(n1376) );
  MUX2X1 U1085 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1663), .Y(n1375) );
  MUX2X1 U1086 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1663), .Y(n1379) );
  MUX2X1 U1087 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1663), .Y(n1378) );
  MUX2X1 U1088 ( .B(n1377), .A(n1374), .S(n1635), .Y(n1388) );
  MUX2X1 U1089 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1663), .Y(n1382) );
  MUX2X1 U1090 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1663), .Y(n1381) );
  MUX2X1 U1091 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1663), .Y(n1385) );
  MUX2X1 U1092 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1663), .Y(n1384) );
  MUX2X1 U1093 ( .B(n1383), .A(n1380), .S(n1635), .Y(n1387) );
  MUX2X1 U1094 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1664), .Y(n1391) );
  MUX2X1 U1095 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1664), .Y(n1390) );
  MUX2X1 U1096 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1664), .Y(n1394) );
  MUX2X1 U1097 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1664), .Y(n1393) );
  MUX2X1 U1098 ( .B(n1392), .A(n1389), .S(n1635), .Y(n1403) );
  MUX2X1 U1099 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1664), .Y(n1397) );
  MUX2X1 U1100 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1664), .Y(n1396) );
  MUX2X1 U1101 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1664), .Y(n1400) );
  MUX2X1 U1102 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1664), .Y(n1399) );
  MUX2X1 U1103 ( .B(n1398), .A(n1395), .S(n1635), .Y(n1402) );
  MUX2X1 U1104 ( .B(n1401), .A(n1386), .S(n1630), .Y(n1622) );
  MUX2X1 U1105 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1664), .Y(n1406) );
  MUX2X1 U1106 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1664), .Y(n1405) );
  MUX2X1 U1107 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1664), .Y(n1409) );
  MUX2X1 U1108 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1664), .Y(n1408) );
  MUX2X1 U1109 ( .B(n1407), .A(n1404), .S(n1634), .Y(n1418) );
  MUX2X1 U1110 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1665), .Y(n1412) );
  MUX2X1 U1111 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1665), .Y(n1411) );
  MUX2X1 U1112 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1665), .Y(n1415) );
  MUX2X1 U1113 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1665), .Y(n1414) );
  MUX2X1 U1114 ( .B(n1413), .A(n1410), .S(n1634), .Y(n1417) );
  MUX2X1 U1115 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1665), .Y(n1421) );
  MUX2X1 U1116 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1665), .Y(n1420) );
  MUX2X1 U1117 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1665), .Y(n1424) );
  MUX2X1 U1118 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1665), .Y(n1423) );
  MUX2X1 U1119 ( .B(n1422), .A(n1419), .S(n1634), .Y(n1433) );
  MUX2X1 U1120 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1665), .Y(n1427) );
  MUX2X1 U1121 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1665), .Y(n1426) );
  MUX2X1 U1122 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1665), .Y(n1430) );
  MUX2X1 U1123 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1665), .Y(n1429) );
  MUX2X1 U1124 ( .B(n1428), .A(n1425), .S(n1634), .Y(n1432) );
  MUX2X1 U1125 ( .B(n1431), .A(n1416), .S(n1630), .Y(n1623) );
  MUX2X1 U1126 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1655), .Y(n1436) );
  MUX2X1 U1127 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1656), .Y(n1435) );
  MUX2X1 U1128 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1656), .Y(n1439) );
  MUX2X1 U1129 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1655), .Y(n1438) );
  MUX2X1 U1130 ( .B(n1437), .A(n1434), .S(n1634), .Y(n1448) );
  MUX2X1 U1131 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1655), .Y(n1442) );
  MUX2X1 U1132 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1656), .Y(n1441) );
  MUX2X1 U1133 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1656), .Y(n1445) );
  MUX2X1 U1134 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1656), .Y(n1444) );
  MUX2X1 U1135 ( .B(n1443), .A(n1440), .S(n1634), .Y(n1447) );
  MUX2X1 U1136 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1655), .Y(n1451) );
  MUX2X1 U1137 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1655), .Y(n1450) );
  MUX2X1 U1138 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1655), .Y(n1454) );
  MUX2X1 U1139 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1655), .Y(n1453) );
  MUX2X1 U1140 ( .B(n1452), .A(n1449), .S(n1634), .Y(n1463) );
  MUX2X1 U1141 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1666), .Y(n1457) );
  MUX2X1 U1142 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1666), .Y(n1456) );
  MUX2X1 U1143 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1666), .Y(n1460) );
  MUX2X1 U1144 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1666), .Y(n1459) );
  MUX2X1 U1145 ( .B(n1458), .A(n1455), .S(n1634), .Y(n1462) );
  MUX2X1 U1146 ( .B(n1461), .A(n1446), .S(n1630), .Y(n1624) );
  MUX2X1 U1147 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1666), .Y(n1466) );
  MUX2X1 U1148 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1666), .Y(n1465) );
  MUX2X1 U1149 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1666), .Y(n1469) );
  MUX2X1 U1150 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1666), .Y(n1468) );
  MUX2X1 U1151 ( .B(n1467), .A(n1464), .S(n1634), .Y(n1478) );
  MUX2X1 U1152 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1666), .Y(n1472) );
  MUX2X1 U1153 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1666), .Y(n1471) );
  MUX2X1 U1154 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1666), .Y(n1475) );
  MUX2X1 U1155 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1666), .Y(n1474) );
  MUX2X1 U1156 ( .B(n1473), .A(n1470), .S(n1634), .Y(n1477) );
  MUX2X1 U1157 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1667), .Y(n1481) );
  MUX2X1 U1158 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1667), .Y(n1480) );
  MUX2X1 U1159 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1667), .Y(n1484) );
  MUX2X1 U1160 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1667), .Y(n1483) );
  MUX2X1 U1161 ( .B(n1482), .A(n1479), .S(n1634), .Y(n1493) );
  MUX2X1 U1162 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1667), .Y(n1487) );
  MUX2X1 U1163 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1667), .Y(n1486) );
  MUX2X1 U1164 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1667), .Y(n1490) );
  MUX2X1 U1165 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1667), .Y(n1489) );
  MUX2X1 U1166 ( .B(n1488), .A(n1485), .S(n1634), .Y(n1492) );
  MUX2X1 U1167 ( .B(n1491), .A(n1476), .S(n1630), .Y(n1625) );
  MUX2X1 U1168 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1667), .Y(n1496) );
  MUX2X1 U1169 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1667), .Y(n1495) );
  MUX2X1 U1170 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1667), .Y(n1499) );
  MUX2X1 U1171 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1667), .Y(n1498) );
  MUX2X1 U1172 ( .B(n1497), .A(n1494), .S(n1634), .Y(n1508) );
  MUX2X1 U1173 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1668), .Y(n1502) );
  MUX2X1 U1174 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1668), .Y(n1501) );
  MUX2X1 U1175 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1668), .Y(n1505) );
  MUX2X1 U1177 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1668), .Y(n1504) );
  MUX2X1 U1178 ( .B(n1503), .A(n1500), .S(n1634), .Y(n1507) );
  MUX2X1 U1179 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1668), .Y(n1511) );
  MUX2X1 U1180 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1668), .Y(n1510) );
  MUX2X1 U1181 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1668), .Y(n1514) );
  MUX2X1 U1182 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1668), .Y(n1513) );
  MUX2X1 U1183 ( .B(n1512), .A(n1509), .S(n1634), .Y(n1523) );
  MUX2X1 U1184 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1668), .Y(n1517) );
  MUX2X1 U1185 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1668), .Y(n1516) );
  MUX2X1 U1186 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1668), .Y(n1520) );
  MUX2X1 U1187 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1668), .Y(n1519) );
  MUX2X1 U1188 ( .B(n1518), .A(n1515), .S(n1634), .Y(n1522) );
  MUX2X1 U1189 ( .B(n1521), .A(n1506), .S(n1630), .Y(n1626) );
  MUX2X1 U1190 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1669), .Y(n1526) );
  MUX2X1 U1191 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1669), .Y(n1525) );
  MUX2X1 U1192 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1669), .Y(n1529) );
  MUX2X1 U1193 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1669), .Y(n1528) );
  MUX2X1 U1194 ( .B(n1527), .A(n1524), .S(n1634), .Y(n1538) );
  MUX2X1 U1195 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1669), .Y(n1532) );
  MUX2X1 U1196 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1669), .Y(n1531) );
  MUX2X1 U1197 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1669), .Y(n1535) );
  MUX2X1 U1198 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1669), .Y(n1534) );
  MUX2X1 U1199 ( .B(n1533), .A(n1530), .S(n1634), .Y(n1537) );
  MUX2X1 U1200 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1669), .Y(n1541) );
  MUX2X1 U1201 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1669), .Y(n1540) );
  MUX2X1 U1202 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1669), .Y(n1544) );
  MUX2X1 U1203 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1669), .Y(n1543) );
  MUX2X1 U1204 ( .B(n1542), .A(n1539), .S(n1634), .Y(n1553) );
  MUX2X1 U1205 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1670), .Y(n1547) );
  MUX2X1 U1206 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1670), .Y(n1546) );
  MUX2X1 U1207 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1670), .Y(n1550) );
  MUX2X1 U1208 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1670), .Y(n1549) );
  MUX2X1 U1209 ( .B(n1548), .A(n1545), .S(n1634), .Y(n1552) );
  MUX2X1 U1210 ( .B(n1551), .A(n1536), .S(n1630), .Y(n1627) );
  MUX2X1 U1211 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1670), .Y(n1556) );
  MUX2X1 U1212 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1670), .Y(n1555) );
  MUX2X1 U1213 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1670), .Y(n1559) );
  MUX2X1 U1214 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1670), .Y(n1558) );
  MUX2X1 U1215 ( .B(n1557), .A(n1554), .S(n1634), .Y(n1568) );
  MUX2X1 U1216 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1670), .Y(n1562) );
  MUX2X1 U1217 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1670), .Y(n1561) );
  MUX2X1 U1218 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1670), .Y(n1565) );
  MUX2X1 U1219 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1670), .Y(n1564) );
  MUX2X1 U1220 ( .B(n1563), .A(n1560), .S(n1634), .Y(n1567) );
  MUX2X1 U1221 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1657), .Y(n1571) );
  MUX2X1 U1222 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1661), .Y(n1570) );
  MUX2X1 U1223 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1657), .Y(n1574) );
  MUX2X1 U1224 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1657), .Y(n1573) );
  MUX2X1 U1225 ( .B(n1572), .A(n1569), .S(n1634), .Y(n1583) );
  MUX2X1 U1226 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1662), .Y(n1577) );
  MUX2X1 U1227 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1663), .Y(n1576) );
  MUX2X1 U1228 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1657), .Y(n1580) );
  MUX2X1 U1229 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1657), .Y(n1579) );
  MUX2X1 U1230 ( .B(n1578), .A(n1575), .S(n1634), .Y(n1582) );
  MUX2X1 U1231 ( .B(n1581), .A(n1566), .S(n1630), .Y(n1628) );
  MUX2X1 U1232 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1663), .Y(n1586) );
  MUX2X1 U1233 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1665), .Y(n1585) );
  MUX2X1 U1234 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1665), .Y(n1589) );
  MUX2X1 U1235 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1661), .Y(n1588) );
  MUX2X1 U1236 ( .B(n1587), .A(n1584), .S(n1634), .Y(n1598) );
  MUX2X1 U1237 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1663), .Y(n1592) );
  MUX2X1 U1238 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1665), .Y(n1591) );
  MUX2X1 U1239 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1657), .Y(n1595) );
  MUX2X1 U1240 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1667), .Y(n1594) );
  MUX2X1 U1241 ( .B(n1593), .A(n1590), .S(n1634), .Y(n1597) );
  MUX2X1 U1242 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1661), .Y(n1601) );
  MUX2X1 U1243 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1657), .Y(n1600) );
  MUX2X1 U1244 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1671), .Y(n1604) );
  MUX2X1 U1245 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1658), .Y(n1603) );
  MUX2X1 U1246 ( .B(n1602), .A(n1599), .S(n1634), .Y(n1613) );
  MUX2X1 U1247 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1657), .Y(n1607) );
  MUX2X1 U1248 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1666), .Y(n1606) );
  MUX2X1 U1249 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1659), .Y(n1610) );
  MUX2X1 U1250 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1660), .Y(n1609) );
  MUX2X1 U1251 ( .B(n1608), .A(n1605), .S(n1634), .Y(n1612) );
  MUX2X1 U1252 ( .B(n1611), .A(n1596), .S(n1630), .Y(n1629) );
  INVX8 U1253 ( .A(n1652), .Y(n1659) );
  INVX8 U1254 ( .A(n1652), .Y(n1660) );
  INVX8 U1255 ( .A(n1652), .Y(n1664) );
  INVX8 U1256 ( .A(n1652), .Y(n1668) );
  INVX1 U1257 ( .A(N11), .Y(n1766) );
  INVX1 U1258 ( .A(N10), .Y(n1764) );
  INVX4 U1259 ( .A(n1773), .Y(n1774) );
  INVX8 U1260 ( .A(n1741), .Y(n1738) );
  INVX8 U1261 ( .A(n1741), .Y(n1739) );
  INVX8 U1262 ( .A(n1741), .Y(n1740) );
  INVX8 U1263 ( .A(n488), .Y(n1741) );
  INVX8 U1264 ( .A(n466), .Y(n1742) );
  INVX8 U1265 ( .A(n466), .Y(n1743) );
  INVX8 U1266 ( .A(n467), .Y(n1744) );
  INVX8 U1267 ( .A(n467), .Y(n1745) );
  INVX8 U1268 ( .A(n468), .Y(n1746) );
  INVX8 U1269 ( .A(n469), .Y(n1747) );
  INVX8 U1270 ( .A(n470), .Y(n1748) );
  INVX8 U1271 ( .A(n470), .Y(n1749) );
  INVX8 U1272 ( .A(n471), .Y(n1750) );
  INVX8 U1273 ( .A(n471), .Y(n1751) );
  INVX8 U1274 ( .A(n472), .Y(n1752) );
  INVX8 U1275 ( .A(n473), .Y(n1753) );
  INVX8 U1276 ( .A(n474), .Y(n1754) );
  INVX8 U1277 ( .A(n474), .Y(n1755) );
  INVX8 U1278 ( .A(n475), .Y(n1756) );
  INVX8 U1279 ( .A(n475), .Y(n1757) );
  INVX8 U1280 ( .A(n476), .Y(n1758) );
  INVX8 U1281 ( .A(n491), .Y(n1759) );
  INVX8 U1282 ( .A(n492), .Y(n1760) );
  INVX8 U1283 ( .A(n493), .Y(n1761) );
  INVX8 U1284 ( .A(n494), .Y(n1762) );
  INVX8 U1285 ( .A(n495), .Y(n1763) );
  OR2X2 U1286 ( .A(rst), .B(write), .Y(n1773) );
  AND2X2 U1287 ( .A(N32), .B(n1774), .Y(\data_out<0> ) );
  AND2X2 U1288 ( .A(N31), .B(n1774), .Y(\data_out<1> ) );
  AND2X2 U1289 ( .A(N30), .B(n1774), .Y(\data_out<2> ) );
  AND2X2 U1290 ( .A(N29), .B(n1774), .Y(\data_out<3> ) );
  AND2X2 U1291 ( .A(N28), .B(n1774), .Y(\data_out<4> ) );
  AND2X2 U1292 ( .A(N27), .B(n1774), .Y(\data_out<5> ) );
  AND2X2 U1293 ( .A(N26), .B(n1774), .Y(\data_out<6> ) );
  AND2X2 U1294 ( .A(N25), .B(n1774), .Y(\data_out<7> ) );
  AND2X2 U1295 ( .A(N24), .B(n1774), .Y(\data_out<8> ) );
  AND2X2 U1296 ( .A(N23), .B(n1774), .Y(\data_out<9> ) );
  AND2X2 U1297 ( .A(N22), .B(n1774), .Y(\data_out<10> ) );
  AND2X2 U1298 ( .A(N21), .B(n1774), .Y(\data_out<11> ) );
  AND2X2 U1299 ( .A(N20), .B(n1774), .Y(\data_out<12> ) );
  AND2X2 U1300 ( .A(N19), .B(n1774), .Y(\data_out<13> ) );
  AND2X2 U1301 ( .A(N18), .B(n1774), .Y(\data_out<14> ) );
  AND2X2 U1302 ( .A(N17), .B(n1774), .Y(\data_out<15> ) );
  NAND2X1 U1303 ( .A(\mem<31><0> ), .B(n1672), .Y(n1775) );
  OAI21X1 U1304 ( .A(n503), .B(n1742), .C(n1775), .Y(n2581) );
  NAND2X1 U1305 ( .A(\mem<31><1> ), .B(n1672), .Y(n1776) );
  OAI21X1 U1306 ( .A(n1745), .B(n503), .C(n1776), .Y(n2580) );
  NAND2X1 U1307 ( .A(\mem<31><2> ), .B(n1672), .Y(n1777) );
  OAI21X1 U1308 ( .A(n1746), .B(n503), .C(n1777), .Y(n2579) );
  NAND2X1 U1309 ( .A(\mem<31><3> ), .B(n1672), .Y(n1778) );
  OAI21X1 U1310 ( .A(n1747), .B(n503), .C(n1778), .Y(n2578) );
  NAND2X1 U1311 ( .A(\mem<31><4> ), .B(n1672), .Y(n1779) );
  OAI21X1 U1312 ( .A(n1749), .B(n503), .C(n1779), .Y(n2577) );
  NAND2X1 U1313 ( .A(\mem<31><5> ), .B(n1672), .Y(n1780) );
  OAI21X1 U1314 ( .A(n1751), .B(n503), .C(n1780), .Y(n2576) );
  NAND2X1 U1315 ( .A(\mem<31><6> ), .B(n1672), .Y(n1781) );
  OAI21X1 U1316 ( .A(n1752), .B(n503), .C(n1781), .Y(n2575) );
  NAND2X1 U1317 ( .A(\mem<31><7> ), .B(n1672), .Y(n1782) );
  OAI21X1 U1318 ( .A(n1753), .B(n503), .C(n1782), .Y(n2574) );
  OAI21X1 U1319 ( .A(n1755), .B(n503), .C(n2), .Y(n2573) );
  OAI21X1 U1320 ( .A(n1756), .B(n503), .C(n4), .Y(n2572) );
  OAI21X1 U1321 ( .A(n1758), .B(n503), .C(n6), .Y(n2571) );
  OAI21X1 U1322 ( .A(n1759), .B(n503), .C(n8), .Y(n2570) );
  OAI21X1 U1323 ( .A(n1760), .B(n503), .C(n10), .Y(n2569) );
  OAI21X1 U1324 ( .A(n1761), .B(n503), .C(n12), .Y(n2568) );
  OAI21X1 U1325 ( .A(n1762), .B(n503), .C(n14), .Y(n2567) );
  OAI21X1 U1326 ( .A(n1763), .B(n503), .C(n16), .Y(n2566) );
  NAND2X1 U1327 ( .A(\mem<30><0> ), .B(n1674), .Y(n1783) );
  OAI21X1 U1328 ( .A(n507), .B(n1742), .C(n1783), .Y(n2565) );
  NAND2X1 U1329 ( .A(\mem<30><1> ), .B(n1674), .Y(n1784) );
  OAI21X1 U1330 ( .A(n507), .B(n1745), .C(n1784), .Y(n2564) );
  NAND2X1 U1331 ( .A(\mem<30><2> ), .B(n1674), .Y(n1785) );
  OAI21X1 U1332 ( .A(n507), .B(n1746), .C(n1785), .Y(n2563) );
  NAND2X1 U1333 ( .A(\mem<30><3> ), .B(n1674), .Y(n1786) );
  OAI21X1 U1334 ( .A(n507), .B(n1747), .C(n1786), .Y(n2562) );
  NAND2X1 U1335 ( .A(\mem<30><4> ), .B(n1674), .Y(n1787) );
  OAI21X1 U1336 ( .A(n507), .B(n1749), .C(n1787), .Y(n2561) );
  NAND2X1 U1337 ( .A(\mem<30><5> ), .B(n1674), .Y(n1788) );
  OAI21X1 U1338 ( .A(n507), .B(n1751), .C(n1788), .Y(n2560) );
  NAND2X1 U1339 ( .A(\mem<30><6> ), .B(n1674), .Y(n1789) );
  OAI21X1 U1340 ( .A(n507), .B(n1752), .C(n1789), .Y(n2559) );
  NAND2X1 U1341 ( .A(\mem<30><7> ), .B(n1674), .Y(n1790) );
  OAI21X1 U1342 ( .A(n507), .B(n1753), .C(n1790), .Y(n2558) );
  OAI21X1 U1343 ( .A(n507), .B(n1754), .C(n18), .Y(n2557) );
  OAI21X1 U1344 ( .A(n507), .B(n1757), .C(n20), .Y(n2556) );
  OAI21X1 U1345 ( .A(n507), .B(n1758), .C(n22), .Y(n2555) );
  OAI21X1 U1346 ( .A(n507), .B(n1759), .C(n24), .Y(n2554) );
  OAI21X1 U1347 ( .A(n507), .B(n1760), .C(n26), .Y(n2553) );
  OAI21X1 U1348 ( .A(n507), .B(n1761), .C(n28), .Y(n2552) );
  OAI21X1 U1349 ( .A(n507), .B(n1762), .C(n30), .Y(n2551) );
  OAI21X1 U1350 ( .A(n507), .B(n1763), .C(n32), .Y(n2550) );
  NAND3X1 U1351 ( .A(n1666), .B(n1636), .C(n1766), .Y(n1791) );
  NAND2X1 U1352 ( .A(\mem<29><0> ), .B(n1676), .Y(n1792) );
  OAI21X1 U1353 ( .A(n511), .B(n1742), .C(n1792), .Y(n2549) );
  NAND2X1 U1354 ( .A(\mem<29><1> ), .B(n1676), .Y(n1793) );
  OAI21X1 U1355 ( .A(n511), .B(n1744), .C(n1793), .Y(n2548) );
  NAND2X1 U1356 ( .A(\mem<29><2> ), .B(n1676), .Y(n1794) );
  OAI21X1 U1357 ( .A(n511), .B(n1746), .C(n1794), .Y(n2547) );
  NAND2X1 U1358 ( .A(\mem<29><3> ), .B(n1676), .Y(n1795) );
  OAI21X1 U1359 ( .A(n511), .B(n1747), .C(n1795), .Y(n2546) );
  NAND2X1 U1360 ( .A(\mem<29><4> ), .B(n1676), .Y(n1796) );
  OAI21X1 U1361 ( .A(n511), .B(n1748), .C(n1796), .Y(n2545) );
  NAND2X1 U1362 ( .A(\mem<29><5> ), .B(n1676), .Y(n1797) );
  OAI21X1 U1363 ( .A(n511), .B(n1750), .C(n1797), .Y(n2544) );
  NAND2X1 U1364 ( .A(\mem<29><6> ), .B(n1676), .Y(n1798) );
  OAI21X1 U1365 ( .A(n511), .B(n1752), .C(n1798), .Y(n2543) );
  NAND2X1 U1366 ( .A(\mem<29><7> ), .B(n1676), .Y(n1799) );
  OAI21X1 U1367 ( .A(n511), .B(n1753), .C(n1799), .Y(n2542) );
  OAI21X1 U1368 ( .A(n511), .B(n1755), .C(n34), .Y(n2541) );
  OAI21X1 U1369 ( .A(n511), .B(n1756), .C(n36), .Y(n2540) );
  OAI21X1 U1370 ( .A(n511), .B(n1758), .C(n38), .Y(n2539) );
  OAI21X1 U1371 ( .A(n511), .B(n1759), .C(n40), .Y(n2538) );
  OAI21X1 U1372 ( .A(n511), .B(n1760), .C(n42), .Y(n2537) );
  OAI21X1 U1373 ( .A(n511), .B(n1761), .C(n44), .Y(n2536) );
  OAI21X1 U1374 ( .A(n511), .B(n1762), .C(n46), .Y(n2535) );
  OAI21X1 U1375 ( .A(n511), .B(n1763), .C(n48), .Y(n2534) );
  NAND3X1 U1376 ( .A(n1635), .B(n1766), .C(n1764), .Y(n1800) );
  NAND2X1 U1377 ( .A(\mem<28><0> ), .B(n1678), .Y(n1801) );
  OAI21X1 U1378 ( .A(n515), .B(n1742), .C(n1801), .Y(n2533) );
  NAND2X1 U1379 ( .A(\mem<28><1> ), .B(n1678), .Y(n1802) );
  OAI21X1 U1380 ( .A(n515), .B(n1745), .C(n1802), .Y(n2532) );
  NAND2X1 U1381 ( .A(\mem<28><2> ), .B(n1678), .Y(n1803) );
  OAI21X1 U1382 ( .A(n515), .B(n1746), .C(n1803), .Y(n2531) );
  NAND2X1 U1383 ( .A(\mem<28><3> ), .B(n1678), .Y(n1804) );
  OAI21X1 U1384 ( .A(n515), .B(n1747), .C(n1804), .Y(n2530) );
  NAND2X1 U1385 ( .A(\mem<28><4> ), .B(n1678), .Y(n1805) );
  OAI21X1 U1386 ( .A(n515), .B(n1749), .C(n1805), .Y(n2529) );
  NAND2X1 U1387 ( .A(\mem<28><5> ), .B(n1678), .Y(n1806) );
  OAI21X1 U1388 ( .A(n515), .B(n1751), .C(n1806), .Y(n2528) );
  NAND2X1 U1389 ( .A(\mem<28><6> ), .B(n1678), .Y(n1807) );
  OAI21X1 U1390 ( .A(n515), .B(n1752), .C(n1807), .Y(n2527) );
  NAND2X1 U1391 ( .A(\mem<28><7> ), .B(n1678), .Y(n1808) );
  OAI21X1 U1392 ( .A(n515), .B(n1753), .C(n1808), .Y(n2526) );
  OAI21X1 U1393 ( .A(n515), .B(n1754), .C(n50), .Y(n2525) );
  OAI21X1 U1394 ( .A(n515), .B(n1757), .C(n52), .Y(n2524) );
  OAI21X1 U1395 ( .A(n515), .B(n1758), .C(n54), .Y(n2523) );
  OAI21X1 U1396 ( .A(n515), .B(n1759), .C(n56), .Y(n2522) );
  OAI21X1 U1397 ( .A(n515), .B(n1760), .C(n58), .Y(n2521) );
  OAI21X1 U1398 ( .A(n515), .B(n1761), .C(n60), .Y(n2520) );
  OAI21X1 U1399 ( .A(n515), .B(n1762), .C(n62), .Y(n2519) );
  OAI21X1 U1400 ( .A(n515), .B(n1763), .C(n64), .Y(n2518) );
  NAND3X1 U1401 ( .A(n1666), .B(n1765), .C(n1767), .Y(n1809) );
  NAND2X1 U1402 ( .A(\mem<27><0> ), .B(n1680), .Y(n1810) );
  OAI21X1 U1403 ( .A(n519), .B(n1742), .C(n1810), .Y(n2517) );
  NAND2X1 U1404 ( .A(\mem<27><1> ), .B(n1680), .Y(n1811) );
  OAI21X1 U1405 ( .A(n519), .B(n1744), .C(n1811), .Y(n2516) );
  NAND2X1 U1406 ( .A(\mem<27><2> ), .B(n1680), .Y(n1812) );
  OAI21X1 U1407 ( .A(n519), .B(n1746), .C(n1812), .Y(n2515) );
  NAND2X1 U1408 ( .A(\mem<27><3> ), .B(n1680), .Y(n1813) );
  OAI21X1 U1409 ( .A(n519), .B(n1747), .C(n1813), .Y(n2514) );
  NAND2X1 U1410 ( .A(\mem<27><4> ), .B(n1680), .Y(n1814) );
  OAI21X1 U1411 ( .A(n519), .B(n1748), .C(n1814), .Y(n2513) );
  NAND2X1 U1412 ( .A(\mem<27><5> ), .B(n1680), .Y(n1815) );
  OAI21X1 U1413 ( .A(n519), .B(n1750), .C(n1815), .Y(n2512) );
  NAND2X1 U1414 ( .A(\mem<27><6> ), .B(n1680), .Y(n1816) );
  OAI21X1 U1415 ( .A(n519), .B(n1752), .C(n1816), .Y(n2511) );
  NAND2X1 U1416 ( .A(\mem<27><7> ), .B(n1680), .Y(n1817) );
  OAI21X1 U1417 ( .A(n519), .B(n1753), .C(n1817), .Y(n2510) );
  OAI21X1 U1418 ( .A(n519), .B(n1755), .C(n66), .Y(n2509) );
  OAI21X1 U1419 ( .A(n519), .B(n1756), .C(n68), .Y(n2508) );
  OAI21X1 U1420 ( .A(n519), .B(n1758), .C(n70), .Y(n2507) );
  OAI21X1 U1421 ( .A(n519), .B(n1759), .C(n72), .Y(n2506) );
  OAI21X1 U1422 ( .A(n519), .B(n1760), .C(n74), .Y(n2505) );
  OAI21X1 U1423 ( .A(n519), .B(n1761), .C(n76), .Y(n2504) );
  OAI21X1 U1424 ( .A(n519), .B(n1762), .C(n78), .Y(n2503) );
  OAI21X1 U1425 ( .A(n519), .B(n1763), .C(n80), .Y(n2502) );
  NAND3X1 U1426 ( .A(n1767), .B(n1765), .C(n1764), .Y(n1818) );
  NAND2X1 U1427 ( .A(\mem<26><0> ), .B(n1682), .Y(n1819) );
  OAI21X1 U1428 ( .A(n523), .B(n1742), .C(n1819), .Y(n2501) );
  NAND2X1 U1429 ( .A(\mem<26><1> ), .B(n1682), .Y(n1820) );
  OAI21X1 U1430 ( .A(n523), .B(n1745), .C(n1820), .Y(n2500) );
  NAND2X1 U1431 ( .A(\mem<26><2> ), .B(n1682), .Y(n1821) );
  OAI21X1 U1432 ( .A(n523), .B(n1746), .C(n1821), .Y(n2499) );
  NAND2X1 U1433 ( .A(\mem<26><3> ), .B(n1682), .Y(n1822) );
  OAI21X1 U1434 ( .A(n523), .B(n1747), .C(n1822), .Y(n2498) );
  NAND2X1 U1435 ( .A(\mem<26><4> ), .B(n1682), .Y(n1823) );
  OAI21X1 U1436 ( .A(n523), .B(n1749), .C(n1823), .Y(n2497) );
  NAND2X1 U1437 ( .A(\mem<26><5> ), .B(n1682), .Y(n1824) );
  OAI21X1 U1438 ( .A(n523), .B(n1751), .C(n1824), .Y(n2496) );
  NAND2X1 U1439 ( .A(\mem<26><6> ), .B(n1682), .Y(n1825) );
  OAI21X1 U1440 ( .A(n523), .B(n1752), .C(n1825), .Y(n2495) );
  NAND2X1 U1441 ( .A(\mem<26><7> ), .B(n1682), .Y(n1826) );
  OAI21X1 U1442 ( .A(n523), .B(n1753), .C(n1826), .Y(n2494) );
  OAI21X1 U1443 ( .A(n523), .B(n1754), .C(n82), .Y(n2493) );
  OAI21X1 U1444 ( .A(n523), .B(n1757), .C(n84), .Y(n2492) );
  OAI21X1 U1445 ( .A(n523), .B(n1758), .C(n86), .Y(n2491) );
  OAI21X1 U1446 ( .A(n523), .B(n1759), .C(n88), .Y(n2490) );
  OAI21X1 U1447 ( .A(n523), .B(n1760), .C(n90), .Y(n2489) );
  OAI21X1 U1448 ( .A(n523), .B(n1761), .C(n92), .Y(n2488) );
  OAI21X1 U1449 ( .A(n523), .B(n1762), .C(n94), .Y(n2487) );
  OAI21X1 U1450 ( .A(n523), .B(n1763), .C(n96), .Y(n2486) );
  NAND3X1 U1451 ( .A(n1667), .B(n1767), .C(n1766), .Y(n1827) );
  NAND2X1 U1452 ( .A(\mem<25><0> ), .B(n1684), .Y(n1828) );
  OAI21X1 U1453 ( .A(n527), .B(n1742), .C(n1828), .Y(n2485) );
  NAND2X1 U1454 ( .A(\mem<25><1> ), .B(n1684), .Y(n1829) );
  OAI21X1 U1455 ( .A(n527), .B(n1744), .C(n1829), .Y(n2484) );
  NAND2X1 U1456 ( .A(\mem<25><2> ), .B(n1684), .Y(n1830) );
  OAI21X1 U1457 ( .A(n527), .B(n1746), .C(n1830), .Y(n2483) );
  NAND2X1 U1458 ( .A(\mem<25><3> ), .B(n1684), .Y(n1831) );
  OAI21X1 U1459 ( .A(n527), .B(n1747), .C(n1831), .Y(n2482) );
  NAND2X1 U1460 ( .A(\mem<25><4> ), .B(n1684), .Y(n1832) );
  OAI21X1 U1461 ( .A(n527), .B(n1748), .C(n1832), .Y(n2481) );
  NAND2X1 U1462 ( .A(\mem<25><5> ), .B(n1684), .Y(n1833) );
  OAI21X1 U1463 ( .A(n527), .B(n1750), .C(n1833), .Y(n2480) );
  NAND2X1 U1464 ( .A(\mem<25><6> ), .B(n1684), .Y(n1834) );
  OAI21X1 U1465 ( .A(n527), .B(n1752), .C(n1834), .Y(n2479) );
  NAND2X1 U1466 ( .A(\mem<25><7> ), .B(n1684), .Y(n1835) );
  OAI21X1 U1467 ( .A(n527), .B(n1753), .C(n1835), .Y(n2478) );
  OAI21X1 U1468 ( .A(n527), .B(n1755), .C(n98), .Y(n2477) );
  OAI21X1 U1469 ( .A(n527), .B(n1756), .C(n100), .Y(n2476) );
  OAI21X1 U1470 ( .A(n527), .B(n1758), .C(n102), .Y(n2475) );
  OAI21X1 U1471 ( .A(n527), .B(n1759), .C(n104), .Y(n2474) );
  OAI21X1 U1472 ( .A(n527), .B(n1760), .C(n106), .Y(n2473) );
  OAI21X1 U1473 ( .A(n527), .B(n1761), .C(n108), .Y(n2472) );
  OAI21X1 U1474 ( .A(n527), .B(n1762), .C(n110), .Y(n2471) );
  OAI21X1 U1475 ( .A(n527), .B(n1763), .C(n112), .Y(n2470) );
  NOR3X1 U1476 ( .A(n1667), .B(n1765), .C(n1637), .Y(n2061) );
  NAND2X1 U1477 ( .A(\mem<24><0> ), .B(n1687), .Y(n1836) );
  OAI21X1 U1478 ( .A(n1686), .B(n1742), .C(n1836), .Y(n2469) );
  NAND2X1 U1479 ( .A(\mem<24><1> ), .B(n1687), .Y(n1837) );
  OAI21X1 U1480 ( .A(n1686), .B(n1744), .C(n1837), .Y(n2468) );
  NAND2X1 U1481 ( .A(\mem<24><2> ), .B(n1687), .Y(n1838) );
  OAI21X1 U1482 ( .A(n1686), .B(n1746), .C(n1838), .Y(n2467) );
  NAND2X1 U1483 ( .A(\mem<24><3> ), .B(n1687), .Y(n1839) );
  OAI21X1 U1484 ( .A(n1686), .B(n1747), .C(n1839), .Y(n2466) );
  NAND2X1 U1485 ( .A(\mem<24><4> ), .B(n1687), .Y(n1840) );
  OAI21X1 U1486 ( .A(n1686), .B(n1748), .C(n1840), .Y(n2465) );
  NAND2X1 U1487 ( .A(\mem<24><5> ), .B(n1687), .Y(n1841) );
  OAI21X1 U1488 ( .A(n1686), .B(n1750), .C(n1841), .Y(n2464) );
  NAND2X1 U1489 ( .A(\mem<24><6> ), .B(n1687), .Y(n1842) );
  OAI21X1 U1490 ( .A(n1686), .B(n1752), .C(n1842), .Y(n2463) );
  NAND2X1 U1491 ( .A(\mem<24><7> ), .B(n1687), .Y(n1843) );
  OAI21X1 U1492 ( .A(n1686), .B(n1753), .C(n1843), .Y(n2462) );
  OAI21X1 U1493 ( .A(n1686), .B(n1754), .C(n114), .Y(n2461) );
  OAI21X1 U1494 ( .A(n1686), .B(n1757), .C(n116), .Y(n2460) );
  OAI21X1 U1495 ( .A(n1686), .B(n1758), .C(n118), .Y(n2459) );
  OAI21X1 U1496 ( .A(n1686), .B(n1759), .C(n120), .Y(n2458) );
  OAI21X1 U1497 ( .A(n1686), .B(n1760), .C(n122), .Y(n2457) );
  OAI21X1 U1498 ( .A(n1686), .B(n1761), .C(n124), .Y(n2456) );
  OAI21X1 U1499 ( .A(n1686), .B(n1762), .C(n126), .Y(n2455) );
  OAI21X1 U1500 ( .A(n1686), .B(n1763), .C(n128), .Y(n2454) );
  NAND2X1 U1501 ( .A(\mem<23><0> ), .B(n1689), .Y(n1844) );
  OAI21X1 U1502 ( .A(n533), .B(n1742), .C(n1844), .Y(n2453) );
  NAND2X1 U1503 ( .A(\mem<23><1> ), .B(n1689), .Y(n1845) );
  OAI21X1 U1504 ( .A(n533), .B(n1745), .C(n1845), .Y(n2452) );
  NAND2X1 U1505 ( .A(\mem<23><2> ), .B(n1689), .Y(n1846) );
  OAI21X1 U1506 ( .A(n533), .B(n1746), .C(n1846), .Y(n2451) );
  NAND2X1 U1507 ( .A(\mem<23><3> ), .B(n1689), .Y(n1847) );
  OAI21X1 U1508 ( .A(n533), .B(n1747), .C(n1847), .Y(n2450) );
  NAND2X1 U1509 ( .A(\mem<23><4> ), .B(n1689), .Y(n1848) );
  OAI21X1 U1510 ( .A(n533), .B(n1749), .C(n1848), .Y(n2449) );
  NAND2X1 U1511 ( .A(\mem<23><5> ), .B(n1689), .Y(n1849) );
  OAI21X1 U1512 ( .A(n533), .B(n1751), .C(n1849), .Y(n2448) );
  NAND2X1 U1513 ( .A(\mem<23><6> ), .B(n1689), .Y(n1850) );
  OAI21X1 U1514 ( .A(n533), .B(n1752), .C(n1850), .Y(n2447) );
  NAND2X1 U1515 ( .A(\mem<23><7> ), .B(n1689), .Y(n1851) );
  OAI21X1 U1516 ( .A(n533), .B(n1753), .C(n1851), .Y(n2446) );
  OAI21X1 U1517 ( .A(n533), .B(n1755), .C(n130), .Y(n2445) );
  OAI21X1 U1518 ( .A(n533), .B(n1757), .C(n132), .Y(n2444) );
  OAI21X1 U1519 ( .A(n533), .B(n1758), .C(n134), .Y(n2443) );
  OAI21X1 U1520 ( .A(n533), .B(n1759), .C(n136), .Y(n2442) );
  OAI21X1 U1521 ( .A(n533), .B(n1760), .C(n138), .Y(n2441) );
  OAI21X1 U1522 ( .A(n533), .B(n1761), .C(n140), .Y(n2440) );
  OAI21X1 U1523 ( .A(n533), .B(n1762), .C(n142), .Y(n2439) );
  OAI21X1 U1524 ( .A(n533), .B(n1763), .C(n144), .Y(n2438) );
  NAND2X1 U1525 ( .A(\mem<22><0> ), .B(n1691), .Y(n1852) );
  OAI21X1 U1526 ( .A(n537), .B(n1742), .C(n1852), .Y(n2437) );
  NAND2X1 U1527 ( .A(\mem<22><1> ), .B(n1691), .Y(n1853) );
  OAI21X1 U1528 ( .A(n537), .B(n1745), .C(n1853), .Y(n2436) );
  NAND2X1 U1529 ( .A(\mem<22><2> ), .B(n1691), .Y(n1854) );
  OAI21X1 U1530 ( .A(n537), .B(n1746), .C(n1854), .Y(n2435) );
  NAND2X1 U1531 ( .A(\mem<22><3> ), .B(n1691), .Y(n1855) );
  OAI21X1 U1532 ( .A(n537), .B(n1747), .C(n1855), .Y(n2434) );
  NAND2X1 U1533 ( .A(\mem<22><4> ), .B(n1691), .Y(n1856) );
  OAI21X1 U1534 ( .A(n537), .B(n1749), .C(n1856), .Y(n2433) );
  NAND2X1 U1535 ( .A(\mem<22><5> ), .B(n1691), .Y(n1857) );
  OAI21X1 U1536 ( .A(n537), .B(n1751), .C(n1857), .Y(n2432) );
  NAND2X1 U1537 ( .A(\mem<22><6> ), .B(n1691), .Y(n1858) );
  OAI21X1 U1538 ( .A(n537), .B(n1752), .C(n1858), .Y(n2431) );
  NAND2X1 U1539 ( .A(\mem<22><7> ), .B(n1691), .Y(n1859) );
  OAI21X1 U1540 ( .A(n537), .B(n1753), .C(n1859), .Y(n2430) );
  OAI21X1 U1541 ( .A(n537), .B(n1755), .C(n146), .Y(n2429) );
  OAI21X1 U1542 ( .A(n537), .B(n1757), .C(n148), .Y(n2428) );
  OAI21X1 U1543 ( .A(n537), .B(n1758), .C(n150), .Y(n2427) );
  OAI21X1 U1544 ( .A(n537), .B(n1759), .C(n152), .Y(n2426) );
  OAI21X1 U1545 ( .A(n537), .B(n1760), .C(n154), .Y(n2425) );
  OAI21X1 U1546 ( .A(n537), .B(n1761), .C(n156), .Y(n2424) );
  OAI21X1 U1547 ( .A(n537), .B(n1762), .C(n158), .Y(n2423) );
  OAI21X1 U1548 ( .A(n537), .B(n1763), .C(n160), .Y(n2422) );
  NAND2X1 U1549 ( .A(\mem<21><0> ), .B(n1693), .Y(n1860) );
  OAI21X1 U1550 ( .A(n541), .B(n1742), .C(n1860), .Y(n2421) );
  NAND2X1 U1551 ( .A(\mem<21><1> ), .B(n1693), .Y(n1861) );
  OAI21X1 U1552 ( .A(n541), .B(n1745), .C(n1861), .Y(n2420) );
  NAND2X1 U1553 ( .A(\mem<21><2> ), .B(n1693), .Y(n1862) );
  OAI21X1 U1554 ( .A(n541), .B(n1746), .C(n1862), .Y(n2419) );
  NAND2X1 U1555 ( .A(\mem<21><3> ), .B(n1693), .Y(n1863) );
  OAI21X1 U1556 ( .A(n541), .B(n1747), .C(n1863), .Y(n2418) );
  NAND2X1 U1557 ( .A(\mem<21><4> ), .B(n1693), .Y(n1864) );
  OAI21X1 U1558 ( .A(n541), .B(n1749), .C(n1864), .Y(n2417) );
  NAND2X1 U1559 ( .A(\mem<21><5> ), .B(n1693), .Y(n1865) );
  OAI21X1 U1560 ( .A(n541), .B(n1751), .C(n1865), .Y(n2416) );
  NAND2X1 U1561 ( .A(\mem<21><6> ), .B(n1693), .Y(n1866) );
  OAI21X1 U1562 ( .A(n541), .B(n1752), .C(n1866), .Y(n2415) );
  NAND2X1 U1563 ( .A(\mem<21><7> ), .B(n1693), .Y(n1867) );
  OAI21X1 U1564 ( .A(n541), .B(n1753), .C(n1867), .Y(n2414) );
  OAI21X1 U1565 ( .A(n541), .B(n1755), .C(n162), .Y(n2413) );
  OAI21X1 U1566 ( .A(n541), .B(n1757), .C(n164), .Y(n2412) );
  OAI21X1 U1567 ( .A(n541), .B(n1758), .C(n166), .Y(n2411) );
  OAI21X1 U1568 ( .A(n541), .B(n1759), .C(n168), .Y(n2410) );
  OAI21X1 U1569 ( .A(n541), .B(n1760), .C(n170), .Y(n2409) );
  OAI21X1 U1570 ( .A(n541), .B(n1761), .C(n172), .Y(n2408) );
  OAI21X1 U1571 ( .A(n541), .B(n1762), .C(n174), .Y(n2407) );
  OAI21X1 U1572 ( .A(n541), .B(n1763), .C(n176), .Y(n2406) );
  NAND2X1 U1573 ( .A(\mem<20><0> ), .B(n1695), .Y(n1868) );
  OAI21X1 U1574 ( .A(n545), .B(n1742), .C(n1868), .Y(n2405) );
  NAND2X1 U1575 ( .A(\mem<20><1> ), .B(n1695), .Y(n1869) );
  OAI21X1 U1576 ( .A(n545), .B(n1745), .C(n1869), .Y(n2404) );
  NAND2X1 U1577 ( .A(\mem<20><2> ), .B(n1695), .Y(n1870) );
  OAI21X1 U1578 ( .A(n545), .B(n1746), .C(n1870), .Y(n2403) );
  NAND2X1 U1579 ( .A(\mem<20><3> ), .B(n1695), .Y(n1871) );
  OAI21X1 U1580 ( .A(n545), .B(n1747), .C(n1871), .Y(n2402) );
  NAND2X1 U1581 ( .A(\mem<20><4> ), .B(n1695), .Y(n1872) );
  OAI21X1 U1582 ( .A(n545), .B(n1749), .C(n1872), .Y(n2401) );
  NAND2X1 U1583 ( .A(\mem<20><5> ), .B(n1695), .Y(n1873) );
  OAI21X1 U1584 ( .A(n545), .B(n1751), .C(n1873), .Y(n2400) );
  NAND2X1 U1585 ( .A(\mem<20><6> ), .B(n1695), .Y(n1874) );
  OAI21X1 U1586 ( .A(n545), .B(n1752), .C(n1874), .Y(n2399) );
  NAND2X1 U1587 ( .A(\mem<20><7> ), .B(n1695), .Y(n1875) );
  OAI21X1 U1588 ( .A(n545), .B(n1753), .C(n1875), .Y(n2398) );
  OAI21X1 U1589 ( .A(n545), .B(n1755), .C(n178), .Y(n2397) );
  OAI21X1 U1590 ( .A(n545), .B(n1757), .C(n180), .Y(n2396) );
  OAI21X1 U1591 ( .A(n545), .B(n1758), .C(n182), .Y(n2395) );
  OAI21X1 U1592 ( .A(n545), .B(n1759), .C(n184), .Y(n2394) );
  OAI21X1 U1593 ( .A(n545), .B(n1760), .C(n186), .Y(n2393) );
  OAI21X1 U1594 ( .A(n545), .B(n1761), .C(n188), .Y(n2392) );
  OAI21X1 U1595 ( .A(n545), .B(n1762), .C(n190), .Y(n2391) );
  OAI21X1 U1596 ( .A(n545), .B(n1763), .C(n192), .Y(n2390) );
  NAND2X1 U1597 ( .A(\mem<19><0> ), .B(n1697), .Y(n1876) );
  OAI21X1 U1598 ( .A(n549), .B(n1743), .C(n1876), .Y(n2389) );
  NAND2X1 U1599 ( .A(\mem<19><1> ), .B(n1697), .Y(n1877) );
  OAI21X1 U1600 ( .A(n549), .B(n1745), .C(n1877), .Y(n2388) );
  NAND2X1 U1601 ( .A(\mem<19><2> ), .B(n1697), .Y(n1878) );
  OAI21X1 U1602 ( .A(n549), .B(n1746), .C(n1878), .Y(n2387) );
  NAND2X1 U1603 ( .A(\mem<19><3> ), .B(n1697), .Y(n1879) );
  OAI21X1 U1604 ( .A(n549), .B(n1747), .C(n1879), .Y(n2386) );
  NAND2X1 U1605 ( .A(\mem<19><4> ), .B(n1697), .Y(n1880) );
  OAI21X1 U1606 ( .A(n549), .B(n1749), .C(n1880), .Y(n2385) );
  NAND2X1 U1607 ( .A(\mem<19><5> ), .B(n1697), .Y(n1881) );
  OAI21X1 U1608 ( .A(n549), .B(n1751), .C(n1881), .Y(n2384) );
  NAND2X1 U1609 ( .A(\mem<19><6> ), .B(n1697), .Y(n1882) );
  OAI21X1 U1610 ( .A(n549), .B(n1752), .C(n1882), .Y(n2383) );
  NAND2X1 U1611 ( .A(\mem<19><7> ), .B(n1697), .Y(n1883) );
  OAI21X1 U1612 ( .A(n549), .B(n1753), .C(n1883), .Y(n2382) );
  OAI21X1 U1613 ( .A(n549), .B(n1755), .C(n194), .Y(n2381) );
  OAI21X1 U1614 ( .A(n549), .B(n1757), .C(n196), .Y(n2380) );
  OAI21X1 U1615 ( .A(n549), .B(n1758), .C(n198), .Y(n2379) );
  OAI21X1 U1616 ( .A(n549), .B(n1759), .C(n200), .Y(n2378) );
  OAI21X1 U1617 ( .A(n549), .B(n1760), .C(n202), .Y(n2377) );
  OAI21X1 U1618 ( .A(n549), .B(n1761), .C(n204), .Y(n2376) );
  OAI21X1 U1619 ( .A(n549), .B(n1762), .C(n206), .Y(n2375) );
  OAI21X1 U1620 ( .A(n549), .B(n1763), .C(n208), .Y(n2374) );
  NAND2X1 U1621 ( .A(\mem<18><0> ), .B(n1699), .Y(n1884) );
  OAI21X1 U1622 ( .A(n553), .B(n1743), .C(n1884), .Y(n2373) );
  NAND2X1 U1623 ( .A(\mem<18><1> ), .B(n1699), .Y(n1885) );
  OAI21X1 U1624 ( .A(n553), .B(n1745), .C(n1885), .Y(n2372) );
  NAND2X1 U1625 ( .A(\mem<18><2> ), .B(n1699), .Y(n1886) );
  OAI21X1 U1626 ( .A(n553), .B(n1746), .C(n1886), .Y(n2371) );
  NAND2X1 U1627 ( .A(\mem<18><3> ), .B(n1699), .Y(n1887) );
  OAI21X1 U1628 ( .A(n553), .B(n1747), .C(n1887), .Y(n2370) );
  NAND2X1 U1629 ( .A(\mem<18><4> ), .B(n1699), .Y(n1888) );
  OAI21X1 U1630 ( .A(n553), .B(n1749), .C(n1888), .Y(n2369) );
  NAND2X1 U1631 ( .A(\mem<18><5> ), .B(n1699), .Y(n1889) );
  OAI21X1 U1632 ( .A(n553), .B(n1751), .C(n1889), .Y(n2368) );
  NAND2X1 U1633 ( .A(\mem<18><6> ), .B(n1699), .Y(n1890) );
  OAI21X1 U1634 ( .A(n553), .B(n1752), .C(n1890), .Y(n2367) );
  NAND2X1 U1635 ( .A(\mem<18><7> ), .B(n1699), .Y(n1891) );
  OAI21X1 U1636 ( .A(n553), .B(n1753), .C(n1891), .Y(n2366) );
  OAI21X1 U1637 ( .A(n553), .B(n1755), .C(n210), .Y(n2365) );
  OAI21X1 U1638 ( .A(n553), .B(n1757), .C(n212), .Y(n2364) );
  OAI21X1 U1639 ( .A(n553), .B(n1758), .C(n215), .Y(n2363) );
  OAI21X1 U1640 ( .A(n553), .B(n1759), .C(n217), .Y(n2362) );
  OAI21X1 U1641 ( .A(n553), .B(n1760), .C(n219), .Y(n2361) );
  OAI21X1 U1642 ( .A(n553), .B(n1761), .C(n221), .Y(n2360) );
  OAI21X1 U1643 ( .A(n553), .B(n1762), .C(n223), .Y(n2359) );
  OAI21X1 U1644 ( .A(n553), .B(n1763), .C(n225), .Y(n2358) );
  NAND2X1 U1645 ( .A(\mem<17><0> ), .B(n1701), .Y(n1892) );
  OAI21X1 U1646 ( .A(n557), .B(n1743), .C(n1892), .Y(n2357) );
  NAND2X1 U1647 ( .A(\mem<17><1> ), .B(n1701), .Y(n1893) );
  OAI21X1 U1648 ( .A(n557), .B(n1745), .C(n1893), .Y(n2356) );
  NAND2X1 U1649 ( .A(\mem<17><2> ), .B(n1701), .Y(n1894) );
  OAI21X1 U1650 ( .A(n557), .B(n1746), .C(n1894), .Y(n2355) );
  NAND2X1 U1651 ( .A(\mem<17><3> ), .B(n1701), .Y(n1895) );
  OAI21X1 U1652 ( .A(n557), .B(n1747), .C(n1895), .Y(n2354) );
  NAND2X1 U1653 ( .A(\mem<17><4> ), .B(n1701), .Y(n1896) );
  OAI21X1 U1654 ( .A(n557), .B(n1749), .C(n1896), .Y(n2353) );
  NAND2X1 U1655 ( .A(\mem<17><5> ), .B(n1701), .Y(n1897) );
  OAI21X1 U1656 ( .A(n557), .B(n1751), .C(n1897), .Y(n2352) );
  NAND2X1 U1657 ( .A(\mem<17><6> ), .B(n1701), .Y(n1898) );
  OAI21X1 U1658 ( .A(n557), .B(n1752), .C(n1898), .Y(n2351) );
  NAND2X1 U1659 ( .A(\mem<17><7> ), .B(n1701), .Y(n1899) );
  OAI21X1 U1660 ( .A(n557), .B(n1753), .C(n1899), .Y(n2350) );
  OAI21X1 U1661 ( .A(n557), .B(n1755), .C(n227), .Y(n2349) );
  OAI21X1 U1662 ( .A(n557), .B(n1757), .C(n229), .Y(n2348) );
  OAI21X1 U1663 ( .A(n557), .B(n1758), .C(n231), .Y(n2347) );
  OAI21X1 U1664 ( .A(n557), .B(n1759), .C(n233), .Y(n2346) );
  OAI21X1 U1665 ( .A(n557), .B(n1760), .C(n235), .Y(n2345) );
  OAI21X1 U1666 ( .A(n557), .B(n1761), .C(n237), .Y(n2344) );
  OAI21X1 U1667 ( .A(n557), .B(n1762), .C(n239), .Y(n2343) );
  OAI21X1 U1668 ( .A(n557), .B(n1763), .C(n241), .Y(n2342) );
  NAND2X1 U1669 ( .A(\mem<16><0> ), .B(n1704), .Y(n1900) );
  OAI21X1 U1670 ( .A(n1703), .B(n1743), .C(n1900), .Y(n2341) );
  NAND2X1 U1671 ( .A(\mem<16><1> ), .B(n1704), .Y(n1901) );
  OAI21X1 U1672 ( .A(n1703), .B(n1745), .C(n1901), .Y(n2340) );
  NAND2X1 U1673 ( .A(\mem<16><2> ), .B(n1704), .Y(n1902) );
  OAI21X1 U1674 ( .A(n1703), .B(n1746), .C(n1902), .Y(n2339) );
  NAND2X1 U1675 ( .A(\mem<16><3> ), .B(n1704), .Y(n1903) );
  OAI21X1 U1676 ( .A(n1703), .B(n1747), .C(n1903), .Y(n2338) );
  NAND2X1 U1677 ( .A(\mem<16><4> ), .B(n1704), .Y(n1904) );
  OAI21X1 U1678 ( .A(n1703), .B(n1749), .C(n1904), .Y(n2337) );
  NAND2X1 U1679 ( .A(\mem<16><5> ), .B(n1704), .Y(n1905) );
  OAI21X1 U1680 ( .A(n1703), .B(n1751), .C(n1905), .Y(n2336) );
  NAND2X1 U1681 ( .A(\mem<16><6> ), .B(n1704), .Y(n1906) );
  OAI21X1 U1682 ( .A(n1703), .B(n1752), .C(n1906), .Y(n2335) );
  NAND2X1 U1683 ( .A(\mem<16><7> ), .B(n1704), .Y(n1907) );
  OAI21X1 U1684 ( .A(n1703), .B(n1753), .C(n1907), .Y(n2334) );
  OAI21X1 U1685 ( .A(n1703), .B(n1755), .C(n243), .Y(n2333) );
  OAI21X1 U1686 ( .A(n1703), .B(n1757), .C(n245), .Y(n2332) );
  OAI21X1 U1687 ( .A(n1703), .B(n1758), .C(n247), .Y(n2331) );
  OAI21X1 U1688 ( .A(n1703), .B(n1759), .C(n249), .Y(n2330) );
  OAI21X1 U1689 ( .A(n1703), .B(n1760), .C(n251), .Y(n2329) );
  OAI21X1 U1690 ( .A(n1703), .B(n1761), .C(n253), .Y(n2328) );
  OAI21X1 U1691 ( .A(n1703), .B(n1762), .C(n255), .Y(n2327) );
  OAI21X1 U1692 ( .A(n1703), .B(n1763), .C(n257), .Y(n2326) );
  NAND3X1 U1693 ( .A(n1768), .B(n2582), .C(n1771), .Y(n1908) );
  NAND2X1 U1694 ( .A(\mem<15><0> ), .B(n1706), .Y(n1909) );
  OAI21X1 U1695 ( .A(n563), .B(n1743), .C(n1909), .Y(n2325) );
  NAND2X1 U1696 ( .A(\mem<15><1> ), .B(n1706), .Y(n1910) );
  OAI21X1 U1697 ( .A(n563), .B(n1745), .C(n1910), .Y(n2324) );
  NAND2X1 U1698 ( .A(\mem<15><2> ), .B(n1706), .Y(n1911) );
  OAI21X1 U1699 ( .A(n563), .B(n1746), .C(n1911), .Y(n2323) );
  NAND2X1 U1700 ( .A(\mem<15><3> ), .B(n1706), .Y(n1912) );
  OAI21X1 U1701 ( .A(n563), .B(n1747), .C(n1912), .Y(n2322) );
  NAND2X1 U1702 ( .A(\mem<15><4> ), .B(n1706), .Y(n1913) );
  OAI21X1 U1703 ( .A(n563), .B(n1749), .C(n1913), .Y(n2321) );
  NAND2X1 U1704 ( .A(\mem<15><5> ), .B(n1706), .Y(n1914) );
  OAI21X1 U1705 ( .A(n563), .B(n1751), .C(n1914), .Y(n2320) );
  NAND2X1 U1706 ( .A(\mem<15><6> ), .B(n1706), .Y(n1915) );
  OAI21X1 U1707 ( .A(n563), .B(n1752), .C(n1915), .Y(n2319) );
  NAND2X1 U1708 ( .A(\mem<15><7> ), .B(n1706), .Y(n1916) );
  OAI21X1 U1709 ( .A(n563), .B(n1753), .C(n1916), .Y(n2318) );
  OAI21X1 U1710 ( .A(n563), .B(n1755), .C(n259), .Y(n2317) );
  OAI21X1 U1711 ( .A(n563), .B(n1757), .C(n261), .Y(n2316) );
  OAI21X1 U1712 ( .A(n563), .B(n1758), .C(n263), .Y(n2315) );
  OAI21X1 U1713 ( .A(n563), .B(n1759), .C(n265), .Y(n2314) );
  OAI21X1 U1714 ( .A(n563), .B(n1760), .C(n267), .Y(n2313) );
  OAI21X1 U1715 ( .A(n563), .B(n1761), .C(n269), .Y(n2312) );
  OAI21X1 U1716 ( .A(n563), .B(n1762), .C(n271), .Y(n2311) );
  OAI21X1 U1717 ( .A(n563), .B(n1763), .C(n273), .Y(n2310) );
  NAND2X1 U1718 ( .A(\mem<14><0> ), .B(n1708), .Y(n1917) );
  OAI21X1 U1719 ( .A(n567), .B(n1743), .C(n1917), .Y(n2309) );
  NAND2X1 U1720 ( .A(\mem<14><1> ), .B(n1708), .Y(n1918) );
  OAI21X1 U1721 ( .A(n567), .B(n1745), .C(n1918), .Y(n2308) );
  NAND2X1 U1722 ( .A(\mem<14><2> ), .B(n1708), .Y(n1919) );
  OAI21X1 U1723 ( .A(n567), .B(n1746), .C(n1919), .Y(n2307) );
  NAND2X1 U1724 ( .A(\mem<14><3> ), .B(n1708), .Y(n1920) );
  OAI21X1 U1725 ( .A(n567), .B(n1747), .C(n1920), .Y(n2306) );
  NAND2X1 U1726 ( .A(\mem<14><4> ), .B(n1708), .Y(n1921) );
  OAI21X1 U1727 ( .A(n567), .B(n1749), .C(n1921), .Y(n2305) );
  NAND2X1 U1728 ( .A(\mem<14><5> ), .B(n1708), .Y(n1922) );
  OAI21X1 U1729 ( .A(n567), .B(n1751), .C(n1922), .Y(n2304) );
  NAND2X1 U1730 ( .A(\mem<14><6> ), .B(n1708), .Y(n1923) );
  OAI21X1 U1731 ( .A(n567), .B(n1752), .C(n1923), .Y(n2303) );
  NAND2X1 U1732 ( .A(\mem<14><7> ), .B(n1708), .Y(n1924) );
  OAI21X1 U1733 ( .A(n567), .B(n1753), .C(n1924), .Y(n2302) );
  OAI21X1 U1734 ( .A(n567), .B(n1755), .C(n275), .Y(n2301) );
  OAI21X1 U1735 ( .A(n567), .B(n1757), .C(n277), .Y(n2300) );
  OAI21X1 U1736 ( .A(n567), .B(n1758), .C(n279), .Y(n2299) );
  OAI21X1 U1737 ( .A(n567), .B(n1759), .C(n281), .Y(n2298) );
  OAI21X1 U1738 ( .A(n567), .B(n1760), .C(n283), .Y(n2297) );
  OAI21X1 U1739 ( .A(n567), .B(n1761), .C(n285), .Y(n2296) );
  OAI21X1 U1740 ( .A(n567), .B(n1762), .C(n287), .Y(n2295) );
  OAI21X1 U1741 ( .A(n567), .B(n1763), .C(n289), .Y(n2294) );
  NAND2X1 U1742 ( .A(\mem<13><0> ), .B(n1710), .Y(n1925) );
  OAI21X1 U1743 ( .A(n571), .B(n1743), .C(n1925), .Y(n2293) );
  NAND2X1 U1744 ( .A(\mem<13><1> ), .B(n1710), .Y(n1926) );
  OAI21X1 U1745 ( .A(n571), .B(n1745), .C(n1926), .Y(n2292) );
  NAND2X1 U1746 ( .A(\mem<13><2> ), .B(n1710), .Y(n1927) );
  OAI21X1 U1747 ( .A(n571), .B(n1746), .C(n1927), .Y(n2291) );
  NAND2X1 U1748 ( .A(\mem<13><3> ), .B(n1710), .Y(n1928) );
  OAI21X1 U1749 ( .A(n571), .B(n1747), .C(n1928), .Y(n2290) );
  NAND2X1 U1750 ( .A(\mem<13><4> ), .B(n1710), .Y(n1929) );
  OAI21X1 U1751 ( .A(n571), .B(n1749), .C(n1929), .Y(n2289) );
  NAND2X1 U1752 ( .A(\mem<13><5> ), .B(n1710), .Y(n1930) );
  OAI21X1 U1753 ( .A(n571), .B(n1751), .C(n1930), .Y(n2288) );
  NAND2X1 U1754 ( .A(\mem<13><6> ), .B(n1710), .Y(n1931) );
  OAI21X1 U1755 ( .A(n571), .B(n1752), .C(n1931), .Y(n2287) );
  NAND2X1 U1756 ( .A(\mem<13><7> ), .B(n1710), .Y(n1932) );
  OAI21X1 U1757 ( .A(n571), .B(n1753), .C(n1932), .Y(n2286) );
  OAI21X1 U1758 ( .A(n571), .B(n1755), .C(n291), .Y(n2285) );
  OAI21X1 U1759 ( .A(n571), .B(n1757), .C(n293), .Y(n2284) );
  OAI21X1 U1760 ( .A(n571), .B(n1758), .C(n295), .Y(n2283) );
  OAI21X1 U1761 ( .A(n571), .B(n1759), .C(n297), .Y(n2282) );
  OAI21X1 U1762 ( .A(n571), .B(n1760), .C(n299), .Y(n2281) );
  OAI21X1 U1763 ( .A(n571), .B(n1761), .C(n301), .Y(n2280) );
  OAI21X1 U1764 ( .A(n571), .B(n1762), .C(n303), .Y(n2279) );
  OAI21X1 U1765 ( .A(n571), .B(n1763), .C(n305), .Y(n2278) );
  NAND2X1 U1766 ( .A(\mem<12><0> ), .B(n1712), .Y(n1933) );
  OAI21X1 U1767 ( .A(n575), .B(n1743), .C(n1933), .Y(n2277) );
  NAND2X1 U1768 ( .A(\mem<12><1> ), .B(n1712), .Y(n1934) );
  OAI21X1 U1769 ( .A(n575), .B(n1745), .C(n1934), .Y(n2276) );
  NAND2X1 U1770 ( .A(\mem<12><2> ), .B(n1712), .Y(n1935) );
  OAI21X1 U1771 ( .A(n575), .B(n1746), .C(n1935), .Y(n2275) );
  NAND2X1 U1772 ( .A(\mem<12><3> ), .B(n1712), .Y(n1936) );
  OAI21X1 U1773 ( .A(n575), .B(n1747), .C(n1936), .Y(n2274) );
  NAND2X1 U1774 ( .A(\mem<12><4> ), .B(n1712), .Y(n1937) );
  OAI21X1 U1775 ( .A(n575), .B(n1749), .C(n1937), .Y(n2273) );
  NAND2X1 U1776 ( .A(\mem<12><5> ), .B(n1712), .Y(n1938) );
  OAI21X1 U1777 ( .A(n575), .B(n1751), .C(n1938), .Y(n2272) );
  NAND2X1 U1778 ( .A(\mem<12><6> ), .B(n1712), .Y(n1939) );
  OAI21X1 U1779 ( .A(n575), .B(n1752), .C(n1939), .Y(n2271) );
  NAND2X1 U1780 ( .A(\mem<12><7> ), .B(n1712), .Y(n1940) );
  OAI21X1 U1781 ( .A(n575), .B(n1753), .C(n1940), .Y(n2270) );
  OAI21X1 U1782 ( .A(n575), .B(n1755), .C(n307), .Y(n2269) );
  OAI21X1 U1783 ( .A(n575), .B(n1757), .C(n309), .Y(n2268) );
  OAI21X1 U1784 ( .A(n575), .B(n1758), .C(n311), .Y(n2267) );
  OAI21X1 U1785 ( .A(n575), .B(n1759), .C(n313), .Y(n2266) );
  OAI21X1 U1786 ( .A(n575), .B(n1760), .C(n315), .Y(n2265) );
  OAI21X1 U1787 ( .A(n575), .B(n1761), .C(n317), .Y(n2264) );
  OAI21X1 U1788 ( .A(n575), .B(n1762), .C(n319), .Y(n2263) );
  OAI21X1 U1789 ( .A(n575), .B(n1763), .C(n321), .Y(n2262) );
  NAND2X1 U1790 ( .A(\mem<11><0> ), .B(n1714), .Y(n1941) );
  OAI21X1 U1791 ( .A(n579), .B(n1743), .C(n1941), .Y(n2261) );
  NAND2X1 U1792 ( .A(\mem<11><1> ), .B(n1714), .Y(n1942) );
  OAI21X1 U1793 ( .A(n579), .B(n1744), .C(n1942), .Y(n2260) );
  NAND2X1 U1794 ( .A(\mem<11><2> ), .B(n1714), .Y(n1943) );
  OAI21X1 U1795 ( .A(n579), .B(n1746), .C(n1943), .Y(n2259) );
  NAND2X1 U1796 ( .A(\mem<11><3> ), .B(n1714), .Y(n1944) );
  OAI21X1 U1797 ( .A(n579), .B(n1747), .C(n1944), .Y(n2258) );
  NAND2X1 U1798 ( .A(\mem<11><4> ), .B(n1714), .Y(n1945) );
  OAI21X1 U1799 ( .A(n579), .B(n1748), .C(n1945), .Y(n2257) );
  NAND2X1 U1800 ( .A(\mem<11><5> ), .B(n1714), .Y(n1946) );
  OAI21X1 U1801 ( .A(n579), .B(n1750), .C(n1946), .Y(n2256) );
  NAND2X1 U1802 ( .A(\mem<11><6> ), .B(n1714), .Y(n1947) );
  OAI21X1 U1803 ( .A(n579), .B(n1752), .C(n1947), .Y(n2255) );
  NAND2X1 U1804 ( .A(\mem<11><7> ), .B(n1714), .Y(n1948) );
  OAI21X1 U1805 ( .A(n579), .B(n1753), .C(n1948), .Y(n2254) );
  OAI21X1 U1806 ( .A(n579), .B(n1754), .C(n323), .Y(n2253) );
  OAI21X1 U1807 ( .A(n579), .B(n1756), .C(n325), .Y(n2252) );
  OAI21X1 U1808 ( .A(n579), .B(n1758), .C(n327), .Y(n2251) );
  OAI21X1 U1809 ( .A(n579), .B(n1759), .C(n329), .Y(n2250) );
  OAI21X1 U1810 ( .A(n579), .B(n1760), .C(n331), .Y(n2249) );
  OAI21X1 U1811 ( .A(n579), .B(n1761), .C(n333), .Y(n2248) );
  OAI21X1 U1812 ( .A(n579), .B(n1762), .C(n335), .Y(n2247) );
  OAI21X1 U1813 ( .A(n579), .B(n1763), .C(n337), .Y(n2246) );
  NAND2X1 U1814 ( .A(\mem<10><0> ), .B(n1716), .Y(n1949) );
  OAI21X1 U1815 ( .A(n583), .B(n1743), .C(n1949), .Y(n2245) );
  NAND2X1 U1816 ( .A(\mem<10><1> ), .B(n1716), .Y(n1950) );
  OAI21X1 U1817 ( .A(n583), .B(n1744), .C(n1950), .Y(n2244) );
  NAND2X1 U1818 ( .A(\mem<10><2> ), .B(n1716), .Y(n1951) );
  OAI21X1 U1819 ( .A(n583), .B(n1746), .C(n1951), .Y(n2243) );
  NAND2X1 U1820 ( .A(\mem<10><3> ), .B(n1716), .Y(n1952) );
  OAI21X1 U1821 ( .A(n583), .B(n1747), .C(n1952), .Y(n2242) );
  NAND2X1 U1822 ( .A(\mem<10><4> ), .B(n1716), .Y(n1953) );
  OAI21X1 U1823 ( .A(n583), .B(n1748), .C(n1953), .Y(n2241) );
  NAND2X1 U1824 ( .A(\mem<10><5> ), .B(n1716), .Y(n1954) );
  OAI21X1 U1825 ( .A(n583), .B(n1750), .C(n1954), .Y(n2240) );
  NAND2X1 U1826 ( .A(\mem<10><6> ), .B(n1716), .Y(n1955) );
  OAI21X1 U1827 ( .A(n583), .B(n1752), .C(n1955), .Y(n2239) );
  NAND2X1 U1828 ( .A(\mem<10><7> ), .B(n1716), .Y(n1956) );
  OAI21X1 U1829 ( .A(n583), .B(n1753), .C(n1956), .Y(n2238) );
  OAI21X1 U1830 ( .A(n583), .B(n1754), .C(n339), .Y(n2237) );
  OAI21X1 U1831 ( .A(n583), .B(n1756), .C(n341), .Y(n2236) );
  OAI21X1 U1832 ( .A(n583), .B(n1758), .C(n343), .Y(n2235) );
  OAI21X1 U1833 ( .A(n583), .B(n1759), .C(n345), .Y(n2234) );
  OAI21X1 U1834 ( .A(n583), .B(n1760), .C(n347), .Y(n2233) );
  OAI21X1 U1835 ( .A(n583), .B(n1761), .C(n349), .Y(n2232) );
  OAI21X1 U1836 ( .A(n583), .B(n1762), .C(n351), .Y(n2231) );
  OAI21X1 U1837 ( .A(n583), .B(n1763), .C(n353), .Y(n2230) );
  NAND2X1 U1838 ( .A(\mem<9><0> ), .B(n1718), .Y(n1957) );
  OAI21X1 U1839 ( .A(n587), .B(n1743), .C(n1957), .Y(n2229) );
  NAND2X1 U1840 ( .A(\mem<9><1> ), .B(n1718), .Y(n1958) );
  OAI21X1 U1841 ( .A(n587), .B(n1744), .C(n1958), .Y(n2228) );
  NAND2X1 U1842 ( .A(\mem<9><2> ), .B(n1718), .Y(n1959) );
  OAI21X1 U1843 ( .A(n587), .B(n1746), .C(n1959), .Y(n2227) );
  NAND2X1 U1844 ( .A(\mem<9><3> ), .B(n1718), .Y(n1960) );
  OAI21X1 U1845 ( .A(n587), .B(n1747), .C(n1960), .Y(n2226) );
  NAND2X1 U1846 ( .A(\mem<9><4> ), .B(n1718), .Y(n1961) );
  OAI21X1 U1847 ( .A(n587), .B(n1748), .C(n1961), .Y(n2225) );
  NAND2X1 U1848 ( .A(\mem<9><5> ), .B(n1718), .Y(n1962) );
  OAI21X1 U1849 ( .A(n587), .B(n1750), .C(n1962), .Y(n2224) );
  NAND2X1 U1850 ( .A(\mem<9><6> ), .B(n1718), .Y(n1963) );
  OAI21X1 U1851 ( .A(n587), .B(n1752), .C(n1963), .Y(n2223) );
  NAND2X1 U1852 ( .A(\mem<9><7> ), .B(n1718), .Y(n1964) );
  OAI21X1 U1853 ( .A(n587), .B(n1753), .C(n1964), .Y(n2222) );
  OAI21X1 U1854 ( .A(n587), .B(n1754), .C(n355), .Y(n2221) );
  OAI21X1 U1855 ( .A(n587), .B(n1756), .C(n357), .Y(n2220) );
  OAI21X1 U1856 ( .A(n587), .B(n1758), .C(n359), .Y(n2219) );
  OAI21X1 U1857 ( .A(n587), .B(n1759), .C(n361), .Y(n2218) );
  OAI21X1 U1858 ( .A(n587), .B(n1760), .C(n363), .Y(n2217) );
  OAI21X1 U1859 ( .A(n587), .B(n1761), .C(n365), .Y(n2216) );
  OAI21X1 U1860 ( .A(n587), .B(n1762), .C(n367), .Y(n2215) );
  OAI21X1 U1861 ( .A(n587), .B(n1763), .C(n369), .Y(n2214) );
  NAND2X1 U1862 ( .A(\mem<8><0> ), .B(n1720), .Y(n1966) );
  OAI21X1 U1863 ( .A(n499), .B(n1743), .C(n1966), .Y(n2213) );
  NAND2X1 U1864 ( .A(\mem<8><1> ), .B(n1720), .Y(n1967) );
  OAI21X1 U1865 ( .A(n499), .B(n1744), .C(n1967), .Y(n2212) );
  NAND2X1 U1866 ( .A(\mem<8><2> ), .B(n1720), .Y(n1968) );
  OAI21X1 U1867 ( .A(n499), .B(n1746), .C(n1968), .Y(n2211) );
  NAND2X1 U1868 ( .A(\mem<8><3> ), .B(n1720), .Y(n1969) );
  OAI21X1 U1869 ( .A(n499), .B(n1747), .C(n1969), .Y(n2210) );
  NAND2X1 U1870 ( .A(\mem<8><4> ), .B(n1720), .Y(n1970) );
  OAI21X1 U1871 ( .A(n499), .B(n1748), .C(n1970), .Y(n2209) );
  NAND2X1 U1872 ( .A(\mem<8><5> ), .B(n1720), .Y(n1971) );
  OAI21X1 U1873 ( .A(n499), .B(n1750), .C(n1971), .Y(n2208) );
  NAND2X1 U1874 ( .A(\mem<8><6> ), .B(n1720), .Y(n1972) );
  OAI21X1 U1875 ( .A(n499), .B(n1752), .C(n1972), .Y(n2207) );
  NAND2X1 U1876 ( .A(\mem<8><7> ), .B(n1720), .Y(n1973) );
  OAI21X1 U1877 ( .A(n499), .B(n1753), .C(n1973), .Y(n2206) );
  NAND2X1 U1878 ( .A(\mem<8><8> ), .B(n1721), .Y(n1974) );
  OAI21X1 U1879 ( .A(n499), .B(n1754), .C(n1974), .Y(n2205) );
  NAND2X1 U1880 ( .A(\mem<8><9> ), .B(n1721), .Y(n1975) );
  OAI21X1 U1881 ( .A(n499), .B(n1756), .C(n1975), .Y(n2204) );
  NAND2X1 U1882 ( .A(\mem<8><10> ), .B(n1721), .Y(n1976) );
  OAI21X1 U1883 ( .A(n499), .B(n1758), .C(n1976), .Y(n2203) );
  OAI21X1 U1884 ( .A(n499), .B(n1759), .C(n371), .Y(n2202) );
  OAI21X1 U1885 ( .A(n499), .B(n1760), .C(n373), .Y(n2201) );
  OAI21X1 U1886 ( .A(n499), .B(n1761), .C(n375), .Y(n2200) );
  OAI21X1 U1887 ( .A(n499), .B(n1762), .C(n377), .Y(n2199) );
  OAI21X1 U1888 ( .A(n499), .B(n1763), .C(n379), .Y(n2198) );
  NAND3X1 U1889 ( .A(n1769), .B(n2582), .C(n1771), .Y(n1977) );
  NAND2X1 U1890 ( .A(\mem<7><0> ), .B(n1722), .Y(n1978) );
  OAI21X1 U1891 ( .A(n593), .B(n1742), .C(n1978), .Y(n2197) );
  NAND2X1 U1892 ( .A(\mem<7><1> ), .B(n1722), .Y(n1979) );
  OAI21X1 U1893 ( .A(n593), .B(n1744), .C(n1979), .Y(n2196) );
  NAND2X1 U1894 ( .A(\mem<7><2> ), .B(n1722), .Y(n1980) );
  OAI21X1 U1895 ( .A(n593), .B(n1746), .C(n1980), .Y(n2195) );
  NAND2X1 U1896 ( .A(\mem<7><3> ), .B(n1722), .Y(n1981) );
  OAI21X1 U1897 ( .A(n593), .B(n1747), .C(n1981), .Y(n2194) );
  NAND2X1 U1898 ( .A(\mem<7><4> ), .B(n1722), .Y(n1982) );
  OAI21X1 U1899 ( .A(n593), .B(n1748), .C(n1982), .Y(n2193) );
  NAND2X1 U1900 ( .A(\mem<7><5> ), .B(n1722), .Y(n1983) );
  OAI21X1 U1901 ( .A(n593), .B(n1750), .C(n1983), .Y(n2192) );
  NAND2X1 U1902 ( .A(\mem<7><6> ), .B(n1722), .Y(n1984) );
  OAI21X1 U1903 ( .A(n593), .B(n1752), .C(n1984), .Y(n2191) );
  NAND2X1 U1904 ( .A(\mem<7><7> ), .B(n1722), .Y(n1985) );
  OAI21X1 U1905 ( .A(n593), .B(n1753), .C(n1985), .Y(n2190) );
  NAND2X1 U1906 ( .A(\mem<7><8> ), .B(n1723), .Y(n1986) );
  OAI21X1 U1907 ( .A(n593), .B(n1754), .C(n1986), .Y(n2189) );
  NAND2X1 U1908 ( .A(\mem<7><9> ), .B(n1723), .Y(n1987) );
  OAI21X1 U1909 ( .A(n593), .B(n1756), .C(n1987), .Y(n2188) );
  NAND2X1 U1910 ( .A(\mem<7><10> ), .B(n1723), .Y(n1988) );
  OAI21X1 U1911 ( .A(n593), .B(n1758), .C(n1988), .Y(n2187) );
  OAI21X1 U1912 ( .A(n593), .B(n1759), .C(n381), .Y(n2186) );
  OAI21X1 U1913 ( .A(n593), .B(n1760), .C(n383), .Y(n2185) );
  OAI21X1 U1914 ( .A(n593), .B(n1761), .C(n385), .Y(n2184) );
  OAI21X1 U1915 ( .A(n593), .B(n1762), .C(n387), .Y(n2183) );
  OAI21X1 U1916 ( .A(n593), .B(n1763), .C(n389), .Y(n2182) );
  NAND2X1 U1917 ( .A(\mem<6><0> ), .B(n1724), .Y(n1989) );
  OAI21X1 U1918 ( .A(n597), .B(n1743), .C(n1989), .Y(n2181) );
  NAND2X1 U1919 ( .A(\mem<6><1> ), .B(n1724), .Y(n1990) );
  OAI21X1 U1920 ( .A(n597), .B(n1744), .C(n1990), .Y(n2180) );
  NAND2X1 U1921 ( .A(\mem<6><2> ), .B(n1724), .Y(n1991) );
  OAI21X1 U1922 ( .A(n597), .B(n1746), .C(n1991), .Y(n2179) );
  NAND2X1 U1923 ( .A(\mem<6><3> ), .B(n1724), .Y(n1992) );
  OAI21X1 U1924 ( .A(n597), .B(n1747), .C(n1992), .Y(n2178) );
  NAND2X1 U1925 ( .A(\mem<6><4> ), .B(n1724), .Y(n1993) );
  OAI21X1 U1926 ( .A(n597), .B(n1748), .C(n1993), .Y(n2177) );
  NAND2X1 U1927 ( .A(\mem<6><5> ), .B(n1724), .Y(n1994) );
  OAI21X1 U1928 ( .A(n597), .B(n1750), .C(n1994), .Y(n2176) );
  NAND2X1 U1929 ( .A(\mem<6><6> ), .B(n1724), .Y(n1995) );
  OAI21X1 U1930 ( .A(n597), .B(n1752), .C(n1995), .Y(n2175) );
  NAND2X1 U1931 ( .A(\mem<6><7> ), .B(n1724), .Y(n1996) );
  OAI21X1 U1932 ( .A(n597), .B(n1753), .C(n1996), .Y(n2174) );
  NAND2X1 U1933 ( .A(\mem<6><8> ), .B(n1725), .Y(n1997) );
  OAI21X1 U1934 ( .A(n597), .B(n1754), .C(n1997), .Y(n2173) );
  NAND2X1 U1935 ( .A(\mem<6><9> ), .B(n1725), .Y(n1998) );
  OAI21X1 U1936 ( .A(n597), .B(n1756), .C(n1998), .Y(n2172) );
  NAND2X1 U1937 ( .A(\mem<6><10> ), .B(n1725), .Y(n1999) );
  OAI21X1 U1938 ( .A(n597), .B(n1758), .C(n1999), .Y(n2171) );
  OAI21X1 U1939 ( .A(n597), .B(n1759), .C(n391), .Y(n2170) );
  OAI21X1 U1940 ( .A(n597), .B(n1760), .C(n393), .Y(n2169) );
  OAI21X1 U1941 ( .A(n597), .B(n1761), .C(n395), .Y(n2168) );
  OAI21X1 U1942 ( .A(n597), .B(n1762), .C(n397), .Y(n2167) );
  OAI21X1 U1943 ( .A(n597), .B(n1763), .C(n399), .Y(n2166) );
  NAND2X1 U1944 ( .A(\mem<5><0> ), .B(n1726), .Y(n2001) );
  OAI21X1 U1945 ( .A(n601), .B(n1742), .C(n2001), .Y(n2165) );
  NAND2X1 U1946 ( .A(\mem<5><1> ), .B(n1726), .Y(n2002) );
  OAI21X1 U1947 ( .A(n601), .B(n1744), .C(n2002), .Y(n2164) );
  NAND2X1 U1948 ( .A(\mem<5><2> ), .B(n1726), .Y(n2003) );
  OAI21X1 U1949 ( .A(n601), .B(n1746), .C(n2003), .Y(n2163) );
  NAND2X1 U1950 ( .A(\mem<5><3> ), .B(n1726), .Y(n2004) );
  OAI21X1 U1951 ( .A(n601), .B(n1747), .C(n2004), .Y(n2162) );
  NAND2X1 U1952 ( .A(\mem<5><4> ), .B(n1726), .Y(n2005) );
  OAI21X1 U1953 ( .A(n601), .B(n1748), .C(n2005), .Y(n2161) );
  NAND2X1 U1954 ( .A(\mem<5><5> ), .B(n1726), .Y(n2006) );
  OAI21X1 U1955 ( .A(n601), .B(n1750), .C(n2006), .Y(n2160) );
  NAND2X1 U1956 ( .A(\mem<5><6> ), .B(n1726), .Y(n2007) );
  OAI21X1 U1957 ( .A(n601), .B(n1752), .C(n2007), .Y(n2159) );
  NAND2X1 U1958 ( .A(\mem<5><7> ), .B(n1726), .Y(n2008) );
  OAI21X1 U1959 ( .A(n601), .B(n1753), .C(n2008), .Y(n2158) );
  NAND2X1 U1960 ( .A(\mem<5><8> ), .B(n1727), .Y(n2009) );
  OAI21X1 U1961 ( .A(n601), .B(n1754), .C(n2009), .Y(n2157) );
  NAND2X1 U1962 ( .A(\mem<5><9> ), .B(n1727), .Y(n2010) );
  OAI21X1 U1963 ( .A(n601), .B(n1756), .C(n2010), .Y(n2156) );
  NAND2X1 U1964 ( .A(\mem<5><10> ), .B(n1727), .Y(n2011) );
  OAI21X1 U1965 ( .A(n601), .B(n1758), .C(n2011), .Y(n2155) );
  OAI21X1 U1966 ( .A(n601), .B(n1759), .C(n401), .Y(n2154) );
  OAI21X1 U1967 ( .A(n601), .B(n1760), .C(n403), .Y(n2153) );
  OAI21X1 U1968 ( .A(n601), .B(n1761), .C(n405), .Y(n2152) );
  OAI21X1 U1969 ( .A(n601), .B(n1762), .C(n407), .Y(n2151) );
  OAI21X1 U1970 ( .A(n601), .B(n1763), .C(n409), .Y(n2150) );
  NAND2X1 U1971 ( .A(\mem<4><0> ), .B(n1728), .Y(n2013) );
  OAI21X1 U1972 ( .A(n605), .B(n1743), .C(n2013), .Y(n2149) );
  NAND2X1 U1973 ( .A(\mem<4><1> ), .B(n1728), .Y(n2014) );
  OAI21X1 U1974 ( .A(n605), .B(n1744), .C(n2014), .Y(n2148) );
  NAND2X1 U1975 ( .A(\mem<4><2> ), .B(n1728), .Y(n2015) );
  OAI21X1 U1976 ( .A(n605), .B(n1746), .C(n2015), .Y(n2147) );
  NAND2X1 U1977 ( .A(\mem<4><3> ), .B(n1728), .Y(n2016) );
  OAI21X1 U1978 ( .A(n605), .B(n1747), .C(n2016), .Y(n2146) );
  NAND2X1 U1979 ( .A(\mem<4><4> ), .B(n1728), .Y(n2017) );
  OAI21X1 U1980 ( .A(n605), .B(n1748), .C(n2017), .Y(n2145) );
  NAND2X1 U1981 ( .A(\mem<4><5> ), .B(n1728), .Y(n2018) );
  OAI21X1 U1982 ( .A(n605), .B(n1750), .C(n2018), .Y(n2144) );
  NAND2X1 U1983 ( .A(\mem<4><6> ), .B(n1728), .Y(n2019) );
  OAI21X1 U1984 ( .A(n605), .B(n1752), .C(n2019), .Y(n2143) );
  NAND2X1 U1985 ( .A(\mem<4><7> ), .B(n1728), .Y(n2020) );
  OAI21X1 U1986 ( .A(n605), .B(n1753), .C(n2020), .Y(n2142) );
  NAND2X1 U1987 ( .A(\mem<4><8> ), .B(n1729), .Y(n2021) );
  OAI21X1 U1988 ( .A(n605), .B(n1754), .C(n2021), .Y(n2141) );
  NAND2X1 U1989 ( .A(\mem<4><9> ), .B(n1729), .Y(n2022) );
  OAI21X1 U1990 ( .A(n605), .B(n1756), .C(n2022), .Y(n2140) );
  NAND2X1 U1991 ( .A(\mem<4><10> ), .B(n1729), .Y(n2023) );
  OAI21X1 U1992 ( .A(n605), .B(n1758), .C(n2023), .Y(n2139) );
  OAI21X1 U1993 ( .A(n605), .B(n1759), .C(n411), .Y(n2138) );
  OAI21X1 U1994 ( .A(n605), .B(n1760), .C(n413), .Y(n2137) );
  OAI21X1 U1995 ( .A(n605), .B(n1761), .C(n415), .Y(n2136) );
  OAI21X1 U1996 ( .A(n605), .B(n1762), .C(n417), .Y(n2135) );
  OAI21X1 U1997 ( .A(n605), .B(n1763), .C(n419), .Y(n2134) );
  NAND2X1 U1998 ( .A(\mem<3><0> ), .B(n1730), .Y(n2025) );
  OAI21X1 U1999 ( .A(n609), .B(n1742), .C(n2025), .Y(n2133) );
  NAND2X1 U2000 ( .A(\mem<3><1> ), .B(n1730), .Y(n2026) );
  OAI21X1 U2001 ( .A(n609), .B(n1744), .C(n2026), .Y(n2132) );
  NAND2X1 U2002 ( .A(\mem<3><2> ), .B(n1730), .Y(n2027) );
  OAI21X1 U2003 ( .A(n609), .B(n1746), .C(n2027), .Y(n2131) );
  NAND2X1 U2004 ( .A(\mem<3><3> ), .B(n1730), .Y(n2028) );
  OAI21X1 U2005 ( .A(n609), .B(n1747), .C(n2028), .Y(n2130) );
  NAND2X1 U2006 ( .A(\mem<3><4> ), .B(n1730), .Y(n2029) );
  OAI21X1 U2007 ( .A(n609), .B(n1748), .C(n2029), .Y(n2129) );
  NAND2X1 U2008 ( .A(\mem<3><5> ), .B(n1730), .Y(n2030) );
  OAI21X1 U2009 ( .A(n609), .B(n1750), .C(n2030), .Y(n2128) );
  NAND2X1 U2010 ( .A(\mem<3><6> ), .B(n1730), .Y(n2031) );
  OAI21X1 U2011 ( .A(n609), .B(n1752), .C(n2031), .Y(n2127) );
  NAND2X1 U2012 ( .A(\mem<3><7> ), .B(n1730), .Y(n2032) );
  OAI21X1 U2013 ( .A(n609), .B(n1753), .C(n2032), .Y(n2126) );
  NAND2X1 U2014 ( .A(\mem<3><8> ), .B(n1731), .Y(n2033) );
  OAI21X1 U2015 ( .A(n609), .B(n1754), .C(n2033), .Y(n2125) );
  NAND2X1 U2016 ( .A(\mem<3><9> ), .B(n1731), .Y(n2034) );
  OAI21X1 U2017 ( .A(n609), .B(n1756), .C(n2034), .Y(n2124) );
  NAND2X1 U2018 ( .A(\mem<3><10> ), .B(n1731), .Y(n2035) );
  OAI21X1 U2019 ( .A(n609), .B(n1758), .C(n2035), .Y(n2123) );
  OAI21X1 U2020 ( .A(n609), .B(n1759), .C(n421), .Y(n2122) );
  OAI21X1 U2021 ( .A(n609), .B(n1760), .C(n423), .Y(n2121) );
  OAI21X1 U2022 ( .A(n609), .B(n1761), .C(n425), .Y(n2120) );
  OAI21X1 U2023 ( .A(n609), .B(n1762), .C(n427), .Y(n2119) );
  OAI21X1 U2024 ( .A(n609), .B(n1763), .C(n429), .Y(n2118) );
  NAND2X1 U2025 ( .A(\mem<2><0> ), .B(n1732), .Y(n2037) );
  OAI21X1 U2026 ( .A(n613), .B(n1743), .C(n2037), .Y(n2117) );
  NAND2X1 U2027 ( .A(\mem<2><1> ), .B(n1732), .Y(n2038) );
  OAI21X1 U2028 ( .A(n613), .B(n1744), .C(n2038), .Y(n2116) );
  NAND2X1 U2029 ( .A(\mem<2><2> ), .B(n1732), .Y(n2039) );
  OAI21X1 U2030 ( .A(n613), .B(n1746), .C(n2039), .Y(n2115) );
  NAND2X1 U2031 ( .A(\mem<2><3> ), .B(n1732), .Y(n2040) );
  OAI21X1 U2032 ( .A(n613), .B(n1747), .C(n2040), .Y(n2114) );
  NAND2X1 U2033 ( .A(\mem<2><4> ), .B(n1732), .Y(n2041) );
  OAI21X1 U2034 ( .A(n613), .B(n1748), .C(n2041), .Y(n2113) );
  NAND2X1 U2035 ( .A(\mem<2><5> ), .B(n1732), .Y(n2042) );
  OAI21X1 U2036 ( .A(n613), .B(n1750), .C(n2042), .Y(n2112) );
  NAND2X1 U2037 ( .A(\mem<2><6> ), .B(n1732), .Y(n2043) );
  OAI21X1 U2038 ( .A(n613), .B(n1752), .C(n2043), .Y(n2111) );
  NAND2X1 U2039 ( .A(\mem<2><7> ), .B(n1732), .Y(n2044) );
  OAI21X1 U2040 ( .A(n613), .B(n1753), .C(n2044), .Y(n2110) );
  NAND2X1 U2041 ( .A(\mem<2><8> ), .B(n1733), .Y(n2045) );
  OAI21X1 U2042 ( .A(n613), .B(n1754), .C(n2045), .Y(n2109) );
  NAND2X1 U2043 ( .A(\mem<2><9> ), .B(n1733), .Y(n2046) );
  OAI21X1 U2044 ( .A(n613), .B(n1756), .C(n2046), .Y(n2108) );
  NAND2X1 U2045 ( .A(\mem<2><10> ), .B(n1733), .Y(n2047) );
  OAI21X1 U2046 ( .A(n613), .B(n1758), .C(n2047), .Y(n2107) );
  OAI21X1 U2047 ( .A(n613), .B(n1759), .C(n431), .Y(n2106) );
  OAI21X1 U2048 ( .A(n613), .B(n1760), .C(n433), .Y(n2105) );
  OAI21X1 U2049 ( .A(n613), .B(n1761), .C(n435), .Y(n2104) );
  OAI21X1 U2050 ( .A(n613), .B(n1762), .C(n437), .Y(n2103) );
  OAI21X1 U2051 ( .A(n613), .B(n1763), .C(n439), .Y(n2102) );
  NAND2X1 U2052 ( .A(\mem<1><0> ), .B(n1734), .Y(n2049) );
  OAI21X1 U2053 ( .A(n617), .B(n1742), .C(n2049), .Y(n2101) );
  NAND2X1 U2054 ( .A(\mem<1><1> ), .B(n1734), .Y(n2050) );
  OAI21X1 U2055 ( .A(n617), .B(n1744), .C(n2050), .Y(n2100) );
  NAND2X1 U2056 ( .A(\mem<1><2> ), .B(n1734), .Y(n2051) );
  OAI21X1 U2057 ( .A(n617), .B(n1746), .C(n2051), .Y(n2099) );
  NAND2X1 U2058 ( .A(\mem<1><3> ), .B(n1734), .Y(n2052) );
  OAI21X1 U2059 ( .A(n617), .B(n1747), .C(n2052), .Y(n2098) );
  NAND2X1 U2060 ( .A(\mem<1><4> ), .B(n1734), .Y(n2053) );
  OAI21X1 U2061 ( .A(n617), .B(n1748), .C(n2053), .Y(n2097) );
  NAND2X1 U2062 ( .A(\mem<1><5> ), .B(n1734), .Y(n2054) );
  OAI21X1 U2063 ( .A(n617), .B(n1750), .C(n2054), .Y(n2096) );
  NAND2X1 U2064 ( .A(\mem<1><6> ), .B(n1734), .Y(n2055) );
  OAI21X1 U2065 ( .A(n617), .B(n1752), .C(n2055), .Y(n2095) );
  NAND2X1 U2066 ( .A(\mem<1><7> ), .B(n1734), .Y(n2056) );
  OAI21X1 U2067 ( .A(n617), .B(n1753), .C(n2056), .Y(n2094) );
  NAND2X1 U2068 ( .A(\mem<1><8> ), .B(n1735), .Y(n2057) );
  OAI21X1 U2069 ( .A(n617), .B(n1754), .C(n2057), .Y(n2093) );
  NAND2X1 U2070 ( .A(\mem<1><9> ), .B(n1735), .Y(n2058) );
  OAI21X1 U2071 ( .A(n617), .B(n1756), .C(n2058), .Y(n2092) );
  NAND2X1 U2072 ( .A(\mem<1><10> ), .B(n1735), .Y(n2059) );
  OAI21X1 U2073 ( .A(n617), .B(n1758), .C(n2059), .Y(n2091) );
  OAI21X1 U2074 ( .A(n617), .B(n1759), .C(n441), .Y(n2090) );
  OAI21X1 U2075 ( .A(n617), .B(n1760), .C(n443), .Y(n2089) );
  OAI21X1 U2076 ( .A(n617), .B(n1761), .C(n445), .Y(n2088) );
  OAI21X1 U2077 ( .A(n617), .B(n1762), .C(n447), .Y(n2087) );
  OAI21X1 U2078 ( .A(n617), .B(n1763), .C(n449), .Y(n2086) );
  NAND2X1 U2079 ( .A(\mem<0><0> ), .B(n1736), .Y(n2062) );
  OAI21X1 U2080 ( .A(n501), .B(n1743), .C(n2062), .Y(n2085) );
  NAND2X1 U2081 ( .A(\mem<0><1> ), .B(n1736), .Y(n2063) );
  OAI21X1 U2082 ( .A(n501), .B(n1744), .C(n2063), .Y(n2084) );
  NAND2X1 U2083 ( .A(\mem<0><2> ), .B(n1736), .Y(n2064) );
  OAI21X1 U2084 ( .A(n501), .B(n1746), .C(n2064), .Y(n2083) );
  NAND2X1 U2085 ( .A(\mem<0><3> ), .B(n1736), .Y(n2065) );
  OAI21X1 U2086 ( .A(n501), .B(n1747), .C(n2065), .Y(n2082) );
  NAND2X1 U2087 ( .A(\mem<0><4> ), .B(n1736), .Y(n2066) );
  OAI21X1 U2088 ( .A(n501), .B(n1748), .C(n2066), .Y(n2081) );
  NAND2X1 U2089 ( .A(\mem<0><5> ), .B(n1736), .Y(n2067) );
  OAI21X1 U2090 ( .A(n501), .B(n1750), .C(n2067), .Y(n2080) );
  NAND2X1 U2091 ( .A(\mem<0><6> ), .B(n1736), .Y(n2068) );
  OAI21X1 U2092 ( .A(n501), .B(n1752), .C(n2068), .Y(n2079) );
  NAND2X1 U2093 ( .A(\mem<0><7> ), .B(n1736), .Y(n2069) );
  OAI21X1 U2094 ( .A(n501), .B(n1753), .C(n2069), .Y(n2078) );
  OAI21X1 U2095 ( .A(n501), .B(n1754), .C(n451), .Y(n2077) );
  OAI21X1 U2096 ( .A(n501), .B(n1756), .C(n453), .Y(n2076) );
  OAI21X1 U2097 ( .A(n501), .B(n1758), .C(n455), .Y(n2075) );
  OAI21X1 U2098 ( .A(n501), .B(n1759), .C(n457), .Y(n2074) );
  OAI21X1 U2099 ( .A(n501), .B(n1760), .C(n459), .Y(n2073) );
  OAI21X1 U2100 ( .A(n501), .B(n1761), .C(n461), .Y(n2072) );
  OAI21X1 U2101 ( .A(n501), .B(n1762), .C(n463), .Y(n2071) );
  OAI21X1 U2102 ( .A(n501), .B(n1763), .C(n465), .Y(n2070) );
endmodule


module memc_Size16_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N31, n2, n3, n4, n5, n6, n7, n9, n11, n13, n15, n17,
         n19, n21, n23, n25, n27, n29, n31, n33, n35, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n47, n48, n50, n52, n54, n56, n58, n60, n62, n64,
         n66, n68, n70, n72, n74, n76, n80, n82, n99, n101, n118, n120, n137,
         n139, n156, n158, n175, n177, n194, n196, n215, n217, n233, n235,
         n251, n253, n269, n271, n287, n289, n305, n307, n323, n325, n341,
         n343, n360, n362, n378, n380, n396, n398, n414, n416, n432, n434,
         n450, n452, n468, n470, n486, n488, n505, n507, n523, n525, n541,
         n543, n559, n561, n577, n579, n595, n597, n613, n615, n631, n633,
         n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1864), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1865), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1866), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1867), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1868), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1869), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1870), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1871), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1872), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1873), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1874), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1875), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1876), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1877), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1878), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1879), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1880), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1881), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1882), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1883), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1884), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1885), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1886), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1887), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1888), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1889), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1890), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1891), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1892), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1893), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1894), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1895), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1896), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1897), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1898), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1899), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1900), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1901), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1902), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1903), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1904), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1905), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1906), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1907), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1908), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1909), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1910), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1911), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1912), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1913), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1914), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1915), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1916), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1917), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1918), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1919), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1920), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1921), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1922), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1923), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1924), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1925), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1926), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1927), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1928), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1929), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1930), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1931), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1932), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1933), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1934), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1935), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1936), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1937), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1938), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1939), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1940), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1941), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1942), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1943), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1944), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1945), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1946), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1947), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1948), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1949), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1950), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1951), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1952), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1953), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1954), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1955), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1956), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1957), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1958), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1959), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1960), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1961), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1962), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1963), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1964), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1965), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1966), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1967), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1968), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1969), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1970), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1971), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1972), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1973), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1974), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1975), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1976), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1977), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1978), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1979), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1980), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1981), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1982), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1983), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1984), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1985), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1986), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1987), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1988), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1989), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1990), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1991), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1992), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1993), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1994), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1995), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1996), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1997), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1998), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1999), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2000), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2001), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2002), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2003), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2004), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2005), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2006), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2007), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2008), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2009), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2010), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2011), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2012), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2013), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2014), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2015), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2016), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2017), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2018), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2019), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2020), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2021), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2022), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2023), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2024), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2025), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2026), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2027), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2028), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2029), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2030), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2031), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2032), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2033), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2034), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2035), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2036), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2037), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2038), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2039), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2040), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2041), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2042), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2043), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2044), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2045), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2046), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2047), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2048), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2049), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2050), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2051), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2052), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2053), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2054), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2055), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2056), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2057), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2058), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2059), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2060), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2061), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2062), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2063), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2064), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2065), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2066), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2067), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2068), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2069), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2070), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2071), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2072), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2073), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2074), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2075), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2076), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2077), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2078), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2079), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2080), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2081), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2082), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2083), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2084), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2085), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2086), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2087), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2088), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2089), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2090), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2091), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2092), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2093), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2094), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2095), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2096), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2097), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2098), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2099), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2100), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2101), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2102), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2103), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2104), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2105), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2106), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2107), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2108), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2109), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2110), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2111), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2112), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2113), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2114), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2115), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2116), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2117), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2118), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2119), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2120), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2121), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2122), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2123), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2124), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2125), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2126), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2127), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2128), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2129), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2130), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2131), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2132), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2133), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2134), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2135), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2136), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2137), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2138), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2139), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2140), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2141), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2142), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2143), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2144), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2145), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2146), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2147), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2148), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2149), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2150), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2151), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2152), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2153), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2154), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2155), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2156), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2157), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2158), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2159), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2160), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2161), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2162), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2163), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2164), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2165), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2166), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2167), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2168), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2169), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2170), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2171), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2172), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2173), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2174), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2175), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2176), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2177), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2178), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2179), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2180), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2181), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2182), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2183), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2184), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2185), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2186), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2187), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2188), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2189), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2190), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2191), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2192), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2193), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2194), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2195), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2196), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2197), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2198), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2199), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2200), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2201), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2202), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2203), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2204), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2205), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2206), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2207), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2208), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2209), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2210), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2211), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2212), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2213), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2214), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2215), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2216), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2217), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2218), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2219), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2220), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2221), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2222), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2223), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2224), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2225), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2226), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2227), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2228), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2229), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2230), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2231), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2232), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2233), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2234), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2235), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2236), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2237), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2238), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2239), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2240), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2241), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2242), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2243), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2244), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2245), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2246), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2247), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2248), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2249), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2250), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2251), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2252), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2253), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2254), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2255), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2256), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2257), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2258), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2259), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2260), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2261), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2262), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2263), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2264), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2265), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2266), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2267), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2268), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2269), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2270), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2271), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2272), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2273), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2274), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2275), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2276), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2277), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2278), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2279), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2280), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2281), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2282), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2283), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2284), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2285), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2286), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2287), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2288), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2289), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2290), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2291), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2292), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2293), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2294), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2295), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2296), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2297), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2298), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2299), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2300), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2301), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2302), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2303), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2304), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2305), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2306), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2307), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2308), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2309), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2310), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2311), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2312), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2313), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2314), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2315), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2316), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2317), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2318), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2319), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2320), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2321), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2322), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2323), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2324), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2325), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2326), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2327), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2328), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2329), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2330), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2331), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2332), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2333), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2334), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2335), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2336), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2337), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2338), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2339), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2340), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2341), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2342), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2343), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2344), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2345), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2346), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2347), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2348), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2349), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2350), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2351), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2352), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2353), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2354), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2355), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2356), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2357), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2358), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2359), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2360), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2361), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2362), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2363), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2364), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2365), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2366), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2367), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2368), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2369), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2370), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2371), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2372), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2373), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2374), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2375), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(n1859), .B(write), .Y(n2885) );
  OAI21X1 U61 ( .A(n1819), .B(n1851), .C(n2901), .Y(n2375) );
  NAND2X1 U62 ( .A(\mem<31><0> ), .B(n1821), .Y(n2901) );
  OAI21X1 U63 ( .A(n1819), .B(n1849), .C(n2900), .Y(n2374) );
  NAND2X1 U64 ( .A(\mem<31><1> ), .B(n1821), .Y(n2900) );
  OAI21X1 U65 ( .A(n1819), .B(n1847), .C(n2899), .Y(n2373) );
  NAND2X1 U66 ( .A(\mem<31><2> ), .B(n1821), .Y(n2899) );
  OAI21X1 U67 ( .A(n1819), .B(n1846), .C(n2898), .Y(n2372) );
  NAND2X1 U68 ( .A(\mem<31><3> ), .B(n1821), .Y(n2898) );
  OAI21X1 U69 ( .A(n1819), .B(n1845), .C(n2897), .Y(n2371) );
  NAND2X1 U70 ( .A(\mem<31><4> ), .B(n1821), .Y(n2897) );
  OAI21X1 U71 ( .A(n1819), .B(n1843), .C(n2896), .Y(n2370) );
  NAND2X1 U72 ( .A(\mem<31><5> ), .B(n1821), .Y(n2896) );
  OAI21X1 U73 ( .A(n1819), .B(n1841), .C(n2895), .Y(n2369) );
  NAND2X1 U74 ( .A(\mem<31><6> ), .B(n1821), .Y(n2895) );
  OAI21X1 U75 ( .A(n1819), .B(n1840), .C(n2894), .Y(n2368) );
  NAND2X1 U76 ( .A(\mem<31><7> ), .B(n1821), .Y(n2894) );
  OAI21X1 U77 ( .A(n1819), .B(n1839), .C(n2893), .Y(n2367) );
  NAND2X1 U78 ( .A(\mem<31><8> ), .B(n1820), .Y(n2893) );
  OAI21X1 U79 ( .A(n1819), .B(n1837), .C(n2892), .Y(n2366) );
  NAND2X1 U80 ( .A(\mem<31><9> ), .B(n1820), .Y(n2892) );
  OAI21X1 U81 ( .A(n1819), .B(n1835), .C(n2891), .Y(n2365) );
  NAND2X1 U82 ( .A(\mem<31><10> ), .B(n1820), .Y(n2891) );
  OAI21X1 U83 ( .A(n1819), .B(n1834), .C(n2890), .Y(n2364) );
  NAND2X1 U84 ( .A(\mem<31><11> ), .B(n1820), .Y(n2890) );
  OAI21X1 U85 ( .A(n1819), .B(n1832), .C(n2889), .Y(n2363) );
  NAND2X1 U86 ( .A(\mem<31><12> ), .B(n1820), .Y(n2889) );
  OAI21X1 U87 ( .A(n1819), .B(n1830), .C(n2888), .Y(n2362) );
  NAND2X1 U88 ( .A(\mem<31><13> ), .B(n1820), .Y(n2888) );
  OAI21X1 U89 ( .A(n1819), .B(n1828), .C(n2887), .Y(n2361) );
  NAND2X1 U90 ( .A(\mem<31><14> ), .B(n1820), .Y(n2887) );
  OAI21X1 U91 ( .A(n1819), .B(n1826), .C(n2886), .Y(n2360) );
  NAND2X1 U92 ( .A(\mem<31><15> ), .B(n1820), .Y(n2886) );
  OAI21X1 U95 ( .A(n1851), .B(n1816), .C(n2883), .Y(n2359) );
  NAND2X1 U96 ( .A(\mem<30><0> ), .B(n1818), .Y(n2883) );
  OAI21X1 U97 ( .A(n1849), .B(n1816), .C(n2882), .Y(n2358) );
  NAND2X1 U98 ( .A(\mem<30><1> ), .B(n1818), .Y(n2882) );
  OAI21X1 U99 ( .A(n1847), .B(n1816), .C(n2881), .Y(n2357) );
  NAND2X1 U100 ( .A(\mem<30><2> ), .B(n1818), .Y(n2881) );
  OAI21X1 U101 ( .A(n1846), .B(n1816), .C(n2880), .Y(n2356) );
  NAND2X1 U102 ( .A(\mem<30><3> ), .B(n1818), .Y(n2880) );
  OAI21X1 U103 ( .A(n1845), .B(n1816), .C(n2879), .Y(n2355) );
  NAND2X1 U104 ( .A(\mem<30><4> ), .B(n1818), .Y(n2879) );
  OAI21X1 U105 ( .A(n1843), .B(n1816), .C(n2878), .Y(n2354) );
  NAND2X1 U106 ( .A(\mem<30><5> ), .B(n1818), .Y(n2878) );
  OAI21X1 U107 ( .A(n1841), .B(n1816), .C(n2877), .Y(n2353) );
  NAND2X1 U108 ( .A(\mem<30><6> ), .B(n1818), .Y(n2877) );
  OAI21X1 U109 ( .A(n1840), .B(n1816), .C(n2876), .Y(n2352) );
  NAND2X1 U110 ( .A(\mem<30><7> ), .B(n1818), .Y(n2876) );
  OAI21X1 U111 ( .A(n1839), .B(n1816), .C(n2875), .Y(n2351) );
  NAND2X1 U112 ( .A(\mem<30><8> ), .B(n1817), .Y(n2875) );
  OAI21X1 U113 ( .A(n1837), .B(n1816), .C(n2874), .Y(n2350) );
  NAND2X1 U114 ( .A(\mem<30><9> ), .B(n1817), .Y(n2874) );
  OAI21X1 U115 ( .A(n1835), .B(n1816), .C(n2873), .Y(n2349) );
  NAND2X1 U116 ( .A(\mem<30><10> ), .B(n1817), .Y(n2873) );
  OAI21X1 U117 ( .A(n1834), .B(n1816), .C(n2872), .Y(n2348) );
  NAND2X1 U118 ( .A(\mem<30><11> ), .B(n1817), .Y(n2872) );
  OAI21X1 U119 ( .A(n1832), .B(n1816), .C(n2871), .Y(n2347) );
  NAND2X1 U120 ( .A(\mem<30><12> ), .B(n1817), .Y(n2871) );
  OAI21X1 U121 ( .A(n1830), .B(n1816), .C(n2870), .Y(n2346) );
  NAND2X1 U122 ( .A(\mem<30><13> ), .B(n1817), .Y(n2870) );
  OAI21X1 U123 ( .A(n1828), .B(n1816), .C(n2869), .Y(n2345) );
  NAND2X1 U124 ( .A(\mem<30><14> ), .B(n1817), .Y(n2869) );
  OAI21X1 U125 ( .A(n1826), .B(n1816), .C(n2868), .Y(n2344) );
  NAND2X1 U126 ( .A(\mem<30><15> ), .B(n1817), .Y(n2868) );
  OAI21X1 U129 ( .A(n1851), .B(n1813), .C(n2866), .Y(n2343) );
  NAND2X1 U130 ( .A(\mem<29><0> ), .B(n1815), .Y(n2866) );
  OAI21X1 U131 ( .A(n1849), .B(n1813), .C(n2865), .Y(n2342) );
  NAND2X1 U132 ( .A(\mem<29><1> ), .B(n1815), .Y(n2865) );
  OAI21X1 U133 ( .A(n1847), .B(n1813), .C(n2864), .Y(n2341) );
  NAND2X1 U134 ( .A(\mem<29><2> ), .B(n1815), .Y(n2864) );
  OAI21X1 U135 ( .A(n1846), .B(n1813), .C(n2863), .Y(n2340) );
  NAND2X1 U136 ( .A(\mem<29><3> ), .B(n1815), .Y(n2863) );
  OAI21X1 U137 ( .A(n1845), .B(n1813), .C(n2862), .Y(n2339) );
  NAND2X1 U138 ( .A(\mem<29><4> ), .B(n1815), .Y(n2862) );
  OAI21X1 U139 ( .A(n1843), .B(n1813), .C(n2861), .Y(n2338) );
  NAND2X1 U140 ( .A(\mem<29><5> ), .B(n1815), .Y(n2861) );
  OAI21X1 U141 ( .A(n1841), .B(n1813), .C(n2860), .Y(n2337) );
  NAND2X1 U142 ( .A(\mem<29><6> ), .B(n1815), .Y(n2860) );
  OAI21X1 U143 ( .A(n1840), .B(n1813), .C(n2859), .Y(n2336) );
  NAND2X1 U144 ( .A(\mem<29><7> ), .B(n1815), .Y(n2859) );
  OAI21X1 U145 ( .A(n1839), .B(n1813), .C(n2858), .Y(n2335) );
  NAND2X1 U146 ( .A(\mem<29><8> ), .B(n1814), .Y(n2858) );
  OAI21X1 U147 ( .A(n1837), .B(n1813), .C(n2857), .Y(n2334) );
  NAND2X1 U148 ( .A(\mem<29><9> ), .B(n1814), .Y(n2857) );
  OAI21X1 U149 ( .A(n1835), .B(n1813), .C(n2856), .Y(n2333) );
  NAND2X1 U150 ( .A(\mem<29><10> ), .B(n1814), .Y(n2856) );
  OAI21X1 U151 ( .A(n1834), .B(n1813), .C(n2855), .Y(n2332) );
  NAND2X1 U152 ( .A(\mem<29><11> ), .B(n1814), .Y(n2855) );
  OAI21X1 U153 ( .A(n1832), .B(n1813), .C(n2854), .Y(n2331) );
  NAND2X1 U154 ( .A(\mem<29><12> ), .B(n1814), .Y(n2854) );
  OAI21X1 U155 ( .A(n1830), .B(n1813), .C(n2853), .Y(n2330) );
  NAND2X1 U156 ( .A(\mem<29><13> ), .B(n1814), .Y(n2853) );
  OAI21X1 U157 ( .A(n1828), .B(n1813), .C(n2852), .Y(n2329) );
  NAND2X1 U158 ( .A(\mem<29><14> ), .B(n1814), .Y(n2852) );
  OAI21X1 U159 ( .A(n1826), .B(n1813), .C(n2851), .Y(n2328) );
  NAND2X1 U160 ( .A(\mem<29><15> ), .B(n1814), .Y(n2851) );
  OAI21X1 U163 ( .A(n1851), .B(n1810), .C(n2849), .Y(n2327) );
  NAND2X1 U164 ( .A(\mem<28><0> ), .B(n1812), .Y(n2849) );
  OAI21X1 U165 ( .A(n1849), .B(n1810), .C(n2848), .Y(n2326) );
  NAND2X1 U166 ( .A(\mem<28><1> ), .B(n1812), .Y(n2848) );
  OAI21X1 U167 ( .A(n1847), .B(n1810), .C(n2847), .Y(n2325) );
  NAND2X1 U168 ( .A(\mem<28><2> ), .B(n1812), .Y(n2847) );
  OAI21X1 U169 ( .A(n1846), .B(n1810), .C(n2846), .Y(n2324) );
  NAND2X1 U170 ( .A(\mem<28><3> ), .B(n1812), .Y(n2846) );
  OAI21X1 U171 ( .A(n1845), .B(n1810), .C(n2845), .Y(n2323) );
  NAND2X1 U172 ( .A(\mem<28><4> ), .B(n1812), .Y(n2845) );
  OAI21X1 U173 ( .A(n1843), .B(n1810), .C(n2844), .Y(n2322) );
  NAND2X1 U174 ( .A(\mem<28><5> ), .B(n1812), .Y(n2844) );
  OAI21X1 U175 ( .A(n1841), .B(n1810), .C(n2843), .Y(n2321) );
  NAND2X1 U176 ( .A(\mem<28><6> ), .B(n1812), .Y(n2843) );
  OAI21X1 U177 ( .A(n1840), .B(n1810), .C(n2842), .Y(n2320) );
  NAND2X1 U178 ( .A(\mem<28><7> ), .B(n1812), .Y(n2842) );
  OAI21X1 U179 ( .A(n1839), .B(n1810), .C(n2841), .Y(n2319) );
  NAND2X1 U180 ( .A(\mem<28><8> ), .B(n1811), .Y(n2841) );
  OAI21X1 U181 ( .A(n1837), .B(n1810), .C(n2840), .Y(n2318) );
  NAND2X1 U182 ( .A(\mem<28><9> ), .B(n1811), .Y(n2840) );
  OAI21X1 U183 ( .A(n1835), .B(n1810), .C(n2839), .Y(n2317) );
  NAND2X1 U184 ( .A(\mem<28><10> ), .B(n1811), .Y(n2839) );
  OAI21X1 U185 ( .A(n1834), .B(n1810), .C(n2838), .Y(n2316) );
  NAND2X1 U186 ( .A(\mem<28><11> ), .B(n1811), .Y(n2838) );
  OAI21X1 U187 ( .A(n1832), .B(n1810), .C(n2837), .Y(n2315) );
  NAND2X1 U188 ( .A(\mem<28><12> ), .B(n1811), .Y(n2837) );
  OAI21X1 U189 ( .A(n1830), .B(n1810), .C(n2836), .Y(n2314) );
  NAND2X1 U190 ( .A(\mem<28><13> ), .B(n1811), .Y(n2836) );
  OAI21X1 U191 ( .A(n1828), .B(n1810), .C(n2835), .Y(n2313) );
  NAND2X1 U192 ( .A(\mem<28><14> ), .B(n1811), .Y(n2835) );
  OAI21X1 U193 ( .A(n1826), .B(n1810), .C(n2834), .Y(n2312) );
  NAND2X1 U194 ( .A(\mem<28><15> ), .B(n1811), .Y(n2834) );
  OAI21X1 U197 ( .A(n1851), .B(n1807), .C(n2832), .Y(n2311) );
  NAND2X1 U198 ( .A(\mem<27><0> ), .B(n1809), .Y(n2832) );
  OAI21X1 U199 ( .A(n1849), .B(n1807), .C(n2831), .Y(n2310) );
  NAND2X1 U200 ( .A(\mem<27><1> ), .B(n1809), .Y(n2831) );
  OAI21X1 U201 ( .A(n1847), .B(n1807), .C(n2830), .Y(n2309) );
  NAND2X1 U202 ( .A(\mem<27><2> ), .B(n1809), .Y(n2830) );
  OAI21X1 U203 ( .A(n1846), .B(n1807), .C(n2829), .Y(n2308) );
  NAND2X1 U204 ( .A(\mem<27><3> ), .B(n1809), .Y(n2829) );
  OAI21X1 U205 ( .A(n1845), .B(n1807), .C(n2828), .Y(n2307) );
  NAND2X1 U206 ( .A(\mem<27><4> ), .B(n1809), .Y(n2828) );
  OAI21X1 U207 ( .A(n1843), .B(n1807), .C(n2827), .Y(n2306) );
  NAND2X1 U208 ( .A(\mem<27><5> ), .B(n1809), .Y(n2827) );
  OAI21X1 U209 ( .A(n1841), .B(n1807), .C(n2826), .Y(n2305) );
  NAND2X1 U210 ( .A(\mem<27><6> ), .B(n1809), .Y(n2826) );
  OAI21X1 U211 ( .A(n1840), .B(n1807), .C(n2825), .Y(n2304) );
  NAND2X1 U212 ( .A(\mem<27><7> ), .B(n1809), .Y(n2825) );
  OAI21X1 U213 ( .A(n1839), .B(n1807), .C(n2824), .Y(n2303) );
  NAND2X1 U214 ( .A(\mem<27><8> ), .B(n1808), .Y(n2824) );
  OAI21X1 U215 ( .A(n1837), .B(n1807), .C(n2823), .Y(n2302) );
  NAND2X1 U216 ( .A(\mem<27><9> ), .B(n1808), .Y(n2823) );
  OAI21X1 U217 ( .A(n1835), .B(n1807), .C(n2822), .Y(n2301) );
  NAND2X1 U218 ( .A(\mem<27><10> ), .B(n1808), .Y(n2822) );
  OAI21X1 U219 ( .A(n1834), .B(n1807), .C(n2821), .Y(n2300) );
  NAND2X1 U220 ( .A(\mem<27><11> ), .B(n1808), .Y(n2821) );
  OAI21X1 U221 ( .A(n1832), .B(n1807), .C(n2820), .Y(n2299) );
  NAND2X1 U222 ( .A(\mem<27><12> ), .B(n1808), .Y(n2820) );
  OAI21X1 U223 ( .A(n1830), .B(n1807), .C(n2819), .Y(n2298) );
  NAND2X1 U224 ( .A(\mem<27><13> ), .B(n1808), .Y(n2819) );
  OAI21X1 U225 ( .A(n1828), .B(n1807), .C(n2818), .Y(n2297) );
  NAND2X1 U226 ( .A(\mem<27><14> ), .B(n1808), .Y(n2818) );
  OAI21X1 U227 ( .A(n1826), .B(n1807), .C(n2817), .Y(n2296) );
  NAND2X1 U228 ( .A(\mem<27><15> ), .B(n1808), .Y(n2817) );
  OAI21X1 U231 ( .A(n1851), .B(n1804), .C(n2815), .Y(n2295) );
  NAND2X1 U232 ( .A(\mem<26><0> ), .B(n1806), .Y(n2815) );
  OAI21X1 U233 ( .A(n1849), .B(n1804), .C(n2814), .Y(n2294) );
  NAND2X1 U234 ( .A(\mem<26><1> ), .B(n1806), .Y(n2814) );
  OAI21X1 U235 ( .A(n1847), .B(n1804), .C(n2813), .Y(n2293) );
  NAND2X1 U236 ( .A(\mem<26><2> ), .B(n1806), .Y(n2813) );
  OAI21X1 U237 ( .A(n1846), .B(n1804), .C(n2812), .Y(n2292) );
  NAND2X1 U238 ( .A(\mem<26><3> ), .B(n1806), .Y(n2812) );
  OAI21X1 U239 ( .A(n1845), .B(n1804), .C(n2811), .Y(n2291) );
  NAND2X1 U240 ( .A(\mem<26><4> ), .B(n1806), .Y(n2811) );
  OAI21X1 U241 ( .A(n1843), .B(n1804), .C(n2810), .Y(n2290) );
  NAND2X1 U242 ( .A(\mem<26><5> ), .B(n1806), .Y(n2810) );
  OAI21X1 U243 ( .A(n1841), .B(n1804), .C(n2809), .Y(n2289) );
  NAND2X1 U244 ( .A(\mem<26><6> ), .B(n1806), .Y(n2809) );
  OAI21X1 U245 ( .A(n1840), .B(n1804), .C(n2808), .Y(n2288) );
  NAND2X1 U246 ( .A(\mem<26><7> ), .B(n1806), .Y(n2808) );
  OAI21X1 U247 ( .A(n1839), .B(n1804), .C(n2807), .Y(n2287) );
  NAND2X1 U248 ( .A(\mem<26><8> ), .B(n1805), .Y(n2807) );
  OAI21X1 U249 ( .A(n1837), .B(n1804), .C(n2806), .Y(n2286) );
  NAND2X1 U250 ( .A(\mem<26><9> ), .B(n1805), .Y(n2806) );
  OAI21X1 U251 ( .A(n1835), .B(n1804), .C(n2805), .Y(n2285) );
  NAND2X1 U252 ( .A(\mem<26><10> ), .B(n1805), .Y(n2805) );
  OAI21X1 U253 ( .A(n1834), .B(n1804), .C(n2804), .Y(n2284) );
  NAND2X1 U254 ( .A(\mem<26><11> ), .B(n1805), .Y(n2804) );
  OAI21X1 U255 ( .A(n1832), .B(n1804), .C(n2803), .Y(n2283) );
  NAND2X1 U256 ( .A(\mem<26><12> ), .B(n1805), .Y(n2803) );
  OAI21X1 U257 ( .A(n1830), .B(n1804), .C(n2802), .Y(n2282) );
  NAND2X1 U258 ( .A(\mem<26><13> ), .B(n1805), .Y(n2802) );
  OAI21X1 U259 ( .A(n1828), .B(n1804), .C(n2801), .Y(n2281) );
  NAND2X1 U260 ( .A(\mem<26><14> ), .B(n1805), .Y(n2801) );
  OAI21X1 U261 ( .A(n1826), .B(n1804), .C(n2800), .Y(n2280) );
  NAND2X1 U262 ( .A(\mem<26><15> ), .B(n1805), .Y(n2800) );
  OAI21X1 U265 ( .A(n1851), .B(n1801), .C(n2798), .Y(n2279) );
  NAND2X1 U266 ( .A(\mem<25><0> ), .B(n1803), .Y(n2798) );
  OAI21X1 U267 ( .A(n1849), .B(n1801), .C(n2797), .Y(n2278) );
  NAND2X1 U268 ( .A(\mem<25><1> ), .B(n1803), .Y(n2797) );
  OAI21X1 U269 ( .A(n1847), .B(n1801), .C(n2796), .Y(n2277) );
  NAND2X1 U270 ( .A(\mem<25><2> ), .B(n1803), .Y(n2796) );
  OAI21X1 U271 ( .A(n1846), .B(n1801), .C(n2795), .Y(n2276) );
  NAND2X1 U272 ( .A(\mem<25><3> ), .B(n1803), .Y(n2795) );
  OAI21X1 U273 ( .A(n1845), .B(n1801), .C(n2794), .Y(n2275) );
  NAND2X1 U274 ( .A(\mem<25><4> ), .B(n1803), .Y(n2794) );
  OAI21X1 U275 ( .A(n1843), .B(n1801), .C(n2793), .Y(n2274) );
  NAND2X1 U276 ( .A(\mem<25><5> ), .B(n1803), .Y(n2793) );
  OAI21X1 U277 ( .A(n1841), .B(n1801), .C(n2792), .Y(n2273) );
  NAND2X1 U278 ( .A(\mem<25><6> ), .B(n1803), .Y(n2792) );
  OAI21X1 U279 ( .A(n1840), .B(n1801), .C(n2791), .Y(n2272) );
  NAND2X1 U280 ( .A(\mem<25><7> ), .B(n1803), .Y(n2791) );
  OAI21X1 U281 ( .A(n1839), .B(n1801), .C(n2790), .Y(n2271) );
  NAND2X1 U282 ( .A(\mem<25><8> ), .B(n1802), .Y(n2790) );
  OAI21X1 U283 ( .A(n1837), .B(n1801), .C(n2789), .Y(n2270) );
  NAND2X1 U284 ( .A(\mem<25><9> ), .B(n1802), .Y(n2789) );
  OAI21X1 U285 ( .A(n1835), .B(n1801), .C(n2788), .Y(n2269) );
  NAND2X1 U286 ( .A(\mem<25><10> ), .B(n1802), .Y(n2788) );
  OAI21X1 U287 ( .A(n1834), .B(n1801), .C(n2787), .Y(n2268) );
  NAND2X1 U288 ( .A(\mem<25><11> ), .B(n1802), .Y(n2787) );
  OAI21X1 U289 ( .A(n1832), .B(n1801), .C(n2786), .Y(n2267) );
  NAND2X1 U290 ( .A(\mem<25><12> ), .B(n1802), .Y(n2786) );
  OAI21X1 U291 ( .A(n1830), .B(n1801), .C(n2785), .Y(n2266) );
  NAND2X1 U292 ( .A(\mem<25><13> ), .B(n1802), .Y(n2785) );
  OAI21X1 U293 ( .A(n1828), .B(n1801), .C(n2784), .Y(n2265) );
  NAND2X1 U294 ( .A(\mem<25><14> ), .B(n1802), .Y(n2784) );
  OAI21X1 U295 ( .A(n1826), .B(n1801), .C(n2783), .Y(n2264) );
  NAND2X1 U296 ( .A(\mem<25><15> ), .B(n1802), .Y(n2783) );
  OAI21X1 U299 ( .A(n1851), .B(n1798), .C(n2781), .Y(n2263) );
  NAND2X1 U300 ( .A(\mem<24><0> ), .B(n1800), .Y(n2781) );
  OAI21X1 U301 ( .A(n1849), .B(n1798), .C(n2780), .Y(n2262) );
  NAND2X1 U302 ( .A(\mem<24><1> ), .B(n1800), .Y(n2780) );
  OAI21X1 U303 ( .A(n1847), .B(n1798), .C(n2779), .Y(n2261) );
  NAND2X1 U304 ( .A(\mem<24><2> ), .B(n1800), .Y(n2779) );
  OAI21X1 U305 ( .A(n1846), .B(n1798), .C(n2778), .Y(n2260) );
  NAND2X1 U306 ( .A(\mem<24><3> ), .B(n1800), .Y(n2778) );
  OAI21X1 U307 ( .A(n1845), .B(n1798), .C(n2777), .Y(n2259) );
  NAND2X1 U308 ( .A(\mem<24><4> ), .B(n1800), .Y(n2777) );
  OAI21X1 U309 ( .A(n1843), .B(n1798), .C(n2776), .Y(n2258) );
  NAND2X1 U310 ( .A(\mem<24><5> ), .B(n1800), .Y(n2776) );
  OAI21X1 U311 ( .A(n1841), .B(n1798), .C(n2775), .Y(n2257) );
  NAND2X1 U312 ( .A(\mem<24><6> ), .B(n1800), .Y(n2775) );
  OAI21X1 U313 ( .A(n1840), .B(n1798), .C(n2774), .Y(n2256) );
  NAND2X1 U314 ( .A(\mem<24><7> ), .B(n1800), .Y(n2774) );
  OAI21X1 U315 ( .A(n1839), .B(n1798), .C(n2773), .Y(n2255) );
  NAND2X1 U316 ( .A(\mem<24><8> ), .B(n1799), .Y(n2773) );
  OAI21X1 U317 ( .A(n1837), .B(n1798), .C(n2772), .Y(n2254) );
  NAND2X1 U318 ( .A(\mem<24><9> ), .B(n1799), .Y(n2772) );
  OAI21X1 U319 ( .A(n1835), .B(n1798), .C(n2771), .Y(n2253) );
  NAND2X1 U320 ( .A(\mem<24><10> ), .B(n1799), .Y(n2771) );
  OAI21X1 U321 ( .A(n1834), .B(n1798), .C(n2770), .Y(n2252) );
  NAND2X1 U322 ( .A(\mem<24><11> ), .B(n1799), .Y(n2770) );
  OAI21X1 U323 ( .A(n1832), .B(n1798), .C(n2769), .Y(n2251) );
  NAND2X1 U324 ( .A(\mem<24><12> ), .B(n1799), .Y(n2769) );
  OAI21X1 U325 ( .A(n1830), .B(n1798), .C(n2768), .Y(n2250) );
  NAND2X1 U326 ( .A(\mem<24><13> ), .B(n1799), .Y(n2768) );
  OAI21X1 U327 ( .A(n1828), .B(n1798), .C(n2767), .Y(n2249) );
  NAND2X1 U328 ( .A(\mem<24><14> ), .B(n1799), .Y(n2767) );
  OAI21X1 U329 ( .A(n1826), .B(n1798), .C(n2766), .Y(n2248) );
  NAND2X1 U330 ( .A(\mem<24><15> ), .B(n1799), .Y(n2766) );
  NAND3X1 U333 ( .A(n1855), .B(n2763), .C(n1857), .Y(n2764) );
  OAI21X1 U334 ( .A(n1851), .B(n1795), .C(n2762), .Y(n2247) );
  NAND2X1 U335 ( .A(\mem<23><0> ), .B(n1797), .Y(n2762) );
  OAI21X1 U336 ( .A(n1849), .B(n1795), .C(n2761), .Y(n2246) );
  NAND2X1 U337 ( .A(\mem<23><1> ), .B(n1797), .Y(n2761) );
  OAI21X1 U338 ( .A(n1847), .B(n1795), .C(n2760), .Y(n2245) );
  NAND2X1 U339 ( .A(\mem<23><2> ), .B(n1797), .Y(n2760) );
  OAI21X1 U340 ( .A(n1846), .B(n1795), .C(n2759), .Y(n2244) );
  NAND2X1 U341 ( .A(\mem<23><3> ), .B(n1797), .Y(n2759) );
  OAI21X1 U342 ( .A(n1845), .B(n1795), .C(n2758), .Y(n2243) );
  NAND2X1 U343 ( .A(\mem<23><4> ), .B(n1797), .Y(n2758) );
  OAI21X1 U344 ( .A(n1843), .B(n1795), .C(n2757), .Y(n2242) );
  NAND2X1 U345 ( .A(\mem<23><5> ), .B(n1797), .Y(n2757) );
  OAI21X1 U346 ( .A(n1841), .B(n1795), .C(n2756), .Y(n2241) );
  NAND2X1 U347 ( .A(\mem<23><6> ), .B(n1797), .Y(n2756) );
  OAI21X1 U348 ( .A(n1840), .B(n1795), .C(n2755), .Y(n2240) );
  NAND2X1 U349 ( .A(\mem<23><7> ), .B(n1797), .Y(n2755) );
  OAI21X1 U350 ( .A(n1839), .B(n1795), .C(n2754), .Y(n2239) );
  NAND2X1 U351 ( .A(\mem<23><8> ), .B(n1796), .Y(n2754) );
  OAI21X1 U352 ( .A(n1837), .B(n1795), .C(n2753), .Y(n2238) );
  NAND2X1 U353 ( .A(\mem<23><9> ), .B(n1796), .Y(n2753) );
  OAI21X1 U354 ( .A(n1835), .B(n1795), .C(n2752), .Y(n2237) );
  NAND2X1 U355 ( .A(\mem<23><10> ), .B(n1796), .Y(n2752) );
  OAI21X1 U356 ( .A(n1834), .B(n1795), .C(n2751), .Y(n2236) );
  NAND2X1 U357 ( .A(\mem<23><11> ), .B(n1796), .Y(n2751) );
  OAI21X1 U358 ( .A(n1832), .B(n1795), .C(n2750), .Y(n2235) );
  NAND2X1 U359 ( .A(\mem<23><12> ), .B(n1796), .Y(n2750) );
  OAI21X1 U360 ( .A(n1830), .B(n1795), .C(n2749), .Y(n2234) );
  NAND2X1 U361 ( .A(\mem<23><13> ), .B(n1796), .Y(n2749) );
  OAI21X1 U362 ( .A(n1828), .B(n1795), .C(n2748), .Y(n2233) );
  NAND2X1 U363 ( .A(\mem<23><14> ), .B(n1796), .Y(n2748) );
  OAI21X1 U364 ( .A(n1826), .B(n1795), .C(n2747), .Y(n2232) );
  NAND2X1 U365 ( .A(\mem<23><15> ), .B(n1796), .Y(n2747) );
  OAI21X1 U368 ( .A(n1851), .B(n1792), .C(n2746), .Y(n2231) );
  NAND2X1 U369 ( .A(\mem<22><0> ), .B(n1794), .Y(n2746) );
  OAI21X1 U370 ( .A(n1849), .B(n1792), .C(n2745), .Y(n2230) );
  NAND2X1 U371 ( .A(\mem<22><1> ), .B(n1794), .Y(n2745) );
  OAI21X1 U372 ( .A(n1847), .B(n1792), .C(n2744), .Y(n2229) );
  NAND2X1 U373 ( .A(\mem<22><2> ), .B(n1794), .Y(n2744) );
  OAI21X1 U374 ( .A(n1846), .B(n1792), .C(n2743), .Y(n2228) );
  NAND2X1 U375 ( .A(\mem<22><3> ), .B(n1794), .Y(n2743) );
  OAI21X1 U376 ( .A(n1845), .B(n1792), .C(n2742), .Y(n2227) );
  NAND2X1 U377 ( .A(\mem<22><4> ), .B(n1794), .Y(n2742) );
  OAI21X1 U378 ( .A(n1843), .B(n1792), .C(n2741), .Y(n2226) );
  NAND2X1 U379 ( .A(\mem<22><5> ), .B(n1794), .Y(n2741) );
  OAI21X1 U380 ( .A(n1841), .B(n1792), .C(n2740), .Y(n2225) );
  NAND2X1 U381 ( .A(\mem<22><6> ), .B(n1794), .Y(n2740) );
  OAI21X1 U382 ( .A(n1840), .B(n1792), .C(n2739), .Y(n2224) );
  NAND2X1 U383 ( .A(\mem<22><7> ), .B(n1794), .Y(n2739) );
  OAI21X1 U384 ( .A(n1839), .B(n1792), .C(n2738), .Y(n2223) );
  NAND2X1 U385 ( .A(\mem<22><8> ), .B(n1793), .Y(n2738) );
  OAI21X1 U386 ( .A(n1837), .B(n1792), .C(n2737), .Y(n2222) );
  NAND2X1 U387 ( .A(\mem<22><9> ), .B(n1793), .Y(n2737) );
  OAI21X1 U388 ( .A(n1835), .B(n1792), .C(n2736), .Y(n2221) );
  NAND2X1 U389 ( .A(\mem<22><10> ), .B(n1793), .Y(n2736) );
  OAI21X1 U390 ( .A(n1834), .B(n1792), .C(n2735), .Y(n2220) );
  NAND2X1 U391 ( .A(\mem<22><11> ), .B(n1793), .Y(n2735) );
  OAI21X1 U392 ( .A(n1832), .B(n1792), .C(n2734), .Y(n2219) );
  NAND2X1 U393 ( .A(\mem<22><12> ), .B(n1793), .Y(n2734) );
  OAI21X1 U394 ( .A(n1830), .B(n1792), .C(n2733), .Y(n2218) );
  NAND2X1 U395 ( .A(\mem<22><13> ), .B(n1793), .Y(n2733) );
  OAI21X1 U396 ( .A(n1828), .B(n1792), .C(n2732), .Y(n2217) );
  NAND2X1 U397 ( .A(\mem<22><14> ), .B(n1793), .Y(n2732) );
  OAI21X1 U398 ( .A(n1826), .B(n1792), .C(n2731), .Y(n2216) );
  NAND2X1 U399 ( .A(\mem<22><15> ), .B(n1793), .Y(n2731) );
  OAI21X1 U402 ( .A(n1851), .B(n1789), .C(n2730), .Y(n2215) );
  NAND2X1 U403 ( .A(\mem<21><0> ), .B(n1791), .Y(n2730) );
  OAI21X1 U404 ( .A(n1849), .B(n1789), .C(n2729), .Y(n2214) );
  NAND2X1 U405 ( .A(\mem<21><1> ), .B(n1791), .Y(n2729) );
  OAI21X1 U406 ( .A(n1847), .B(n1789), .C(n2728), .Y(n2213) );
  NAND2X1 U407 ( .A(\mem<21><2> ), .B(n1791), .Y(n2728) );
  OAI21X1 U408 ( .A(n1846), .B(n1789), .C(n2727), .Y(n2212) );
  NAND2X1 U409 ( .A(\mem<21><3> ), .B(n1791), .Y(n2727) );
  OAI21X1 U410 ( .A(n1845), .B(n1789), .C(n2726), .Y(n2211) );
  NAND2X1 U411 ( .A(\mem<21><4> ), .B(n1791), .Y(n2726) );
  OAI21X1 U412 ( .A(n1843), .B(n1789), .C(n2725), .Y(n2210) );
  NAND2X1 U413 ( .A(\mem<21><5> ), .B(n1791), .Y(n2725) );
  OAI21X1 U414 ( .A(n1841), .B(n1789), .C(n2724), .Y(n2209) );
  NAND2X1 U415 ( .A(\mem<21><6> ), .B(n1791), .Y(n2724) );
  OAI21X1 U416 ( .A(n1840), .B(n1789), .C(n2723), .Y(n2208) );
  NAND2X1 U417 ( .A(\mem<21><7> ), .B(n1791), .Y(n2723) );
  OAI21X1 U418 ( .A(n1839), .B(n1789), .C(n2722), .Y(n2207) );
  NAND2X1 U419 ( .A(\mem<21><8> ), .B(n1790), .Y(n2722) );
  OAI21X1 U420 ( .A(n1837), .B(n1789), .C(n2721), .Y(n2206) );
  NAND2X1 U421 ( .A(\mem<21><9> ), .B(n1790), .Y(n2721) );
  OAI21X1 U422 ( .A(n1835), .B(n1789), .C(n2720), .Y(n2205) );
  NAND2X1 U423 ( .A(\mem<21><10> ), .B(n1790), .Y(n2720) );
  OAI21X1 U424 ( .A(n1834), .B(n1789), .C(n2719), .Y(n2204) );
  NAND2X1 U425 ( .A(\mem<21><11> ), .B(n1790), .Y(n2719) );
  OAI21X1 U426 ( .A(n1832), .B(n1789), .C(n2718), .Y(n2203) );
  NAND2X1 U427 ( .A(\mem<21><12> ), .B(n1790), .Y(n2718) );
  OAI21X1 U428 ( .A(n1830), .B(n1789), .C(n2717), .Y(n2202) );
  NAND2X1 U429 ( .A(\mem<21><13> ), .B(n1790), .Y(n2717) );
  OAI21X1 U430 ( .A(n1828), .B(n1789), .C(n2716), .Y(n2201) );
  NAND2X1 U431 ( .A(\mem<21><14> ), .B(n1790), .Y(n2716) );
  OAI21X1 U432 ( .A(n1826), .B(n1789), .C(n2715), .Y(n2200) );
  NAND2X1 U433 ( .A(\mem<21><15> ), .B(n1790), .Y(n2715) );
  OAI21X1 U436 ( .A(n1851), .B(n1786), .C(n2714), .Y(n2199) );
  NAND2X1 U437 ( .A(\mem<20><0> ), .B(n1788), .Y(n2714) );
  OAI21X1 U438 ( .A(n1849), .B(n1786), .C(n2713), .Y(n2198) );
  NAND2X1 U439 ( .A(\mem<20><1> ), .B(n1788), .Y(n2713) );
  OAI21X1 U440 ( .A(n1847), .B(n1786), .C(n2712), .Y(n2197) );
  NAND2X1 U441 ( .A(\mem<20><2> ), .B(n1788), .Y(n2712) );
  OAI21X1 U442 ( .A(n1846), .B(n1786), .C(n2711), .Y(n2196) );
  NAND2X1 U443 ( .A(\mem<20><3> ), .B(n1788), .Y(n2711) );
  OAI21X1 U444 ( .A(n1845), .B(n1786), .C(n2710), .Y(n2195) );
  NAND2X1 U445 ( .A(\mem<20><4> ), .B(n1788), .Y(n2710) );
  OAI21X1 U446 ( .A(n1843), .B(n1786), .C(n2709), .Y(n2194) );
  NAND2X1 U447 ( .A(\mem<20><5> ), .B(n1788), .Y(n2709) );
  OAI21X1 U448 ( .A(n1841), .B(n1786), .C(n2708), .Y(n2193) );
  NAND2X1 U449 ( .A(\mem<20><6> ), .B(n1788), .Y(n2708) );
  OAI21X1 U450 ( .A(n1840), .B(n1786), .C(n2707), .Y(n2192) );
  NAND2X1 U451 ( .A(\mem<20><7> ), .B(n1788), .Y(n2707) );
  OAI21X1 U452 ( .A(n1839), .B(n1786), .C(n2706), .Y(n2191) );
  NAND2X1 U453 ( .A(\mem<20><8> ), .B(n1787), .Y(n2706) );
  OAI21X1 U454 ( .A(n1837), .B(n1786), .C(n2705), .Y(n2190) );
  NAND2X1 U455 ( .A(\mem<20><9> ), .B(n1787), .Y(n2705) );
  OAI21X1 U456 ( .A(n1835), .B(n1786), .C(n2704), .Y(n2189) );
  NAND2X1 U457 ( .A(\mem<20><10> ), .B(n1787), .Y(n2704) );
  OAI21X1 U458 ( .A(n1834), .B(n1786), .C(n2703), .Y(n2188) );
  NAND2X1 U459 ( .A(\mem<20><11> ), .B(n1787), .Y(n2703) );
  OAI21X1 U460 ( .A(n1832), .B(n1786), .C(n2702), .Y(n2187) );
  NAND2X1 U461 ( .A(\mem<20><12> ), .B(n1787), .Y(n2702) );
  OAI21X1 U462 ( .A(n1830), .B(n1786), .C(n2701), .Y(n2186) );
  NAND2X1 U463 ( .A(\mem<20><13> ), .B(n1787), .Y(n2701) );
  OAI21X1 U464 ( .A(n1828), .B(n1786), .C(n2700), .Y(n2185) );
  NAND2X1 U465 ( .A(\mem<20><14> ), .B(n1787), .Y(n2700) );
  OAI21X1 U466 ( .A(n1826), .B(n1786), .C(n2699), .Y(n2184) );
  NAND2X1 U467 ( .A(\mem<20><15> ), .B(n1787), .Y(n2699) );
  OAI21X1 U470 ( .A(n1851), .B(n1783), .C(n2698), .Y(n2183) );
  NAND2X1 U471 ( .A(\mem<19><0> ), .B(n1785), .Y(n2698) );
  OAI21X1 U472 ( .A(n1849), .B(n1783), .C(n2697), .Y(n2182) );
  NAND2X1 U473 ( .A(\mem<19><1> ), .B(n1785), .Y(n2697) );
  OAI21X1 U474 ( .A(n1847), .B(n1783), .C(n2696), .Y(n2181) );
  NAND2X1 U475 ( .A(\mem<19><2> ), .B(n1785), .Y(n2696) );
  OAI21X1 U476 ( .A(n1846), .B(n1783), .C(n2695), .Y(n2180) );
  NAND2X1 U477 ( .A(\mem<19><3> ), .B(n1785), .Y(n2695) );
  OAI21X1 U478 ( .A(n1845), .B(n1783), .C(n2694), .Y(n2179) );
  NAND2X1 U479 ( .A(\mem<19><4> ), .B(n1785), .Y(n2694) );
  OAI21X1 U480 ( .A(n1843), .B(n1783), .C(n2693), .Y(n2178) );
  NAND2X1 U481 ( .A(\mem<19><5> ), .B(n1785), .Y(n2693) );
  OAI21X1 U482 ( .A(n1841), .B(n1783), .C(n2692), .Y(n2177) );
  NAND2X1 U483 ( .A(\mem<19><6> ), .B(n1785), .Y(n2692) );
  OAI21X1 U484 ( .A(n1840), .B(n1783), .C(n2691), .Y(n2176) );
  NAND2X1 U485 ( .A(\mem<19><7> ), .B(n1785), .Y(n2691) );
  OAI21X1 U486 ( .A(n1839), .B(n1783), .C(n2690), .Y(n2175) );
  NAND2X1 U487 ( .A(\mem<19><8> ), .B(n1784), .Y(n2690) );
  OAI21X1 U488 ( .A(n1837), .B(n1783), .C(n2689), .Y(n2174) );
  NAND2X1 U489 ( .A(\mem<19><9> ), .B(n1784), .Y(n2689) );
  OAI21X1 U490 ( .A(n1835), .B(n1783), .C(n2688), .Y(n2173) );
  NAND2X1 U491 ( .A(\mem<19><10> ), .B(n1784), .Y(n2688) );
  OAI21X1 U492 ( .A(n1834), .B(n1783), .C(n2687), .Y(n2172) );
  NAND2X1 U493 ( .A(\mem<19><11> ), .B(n1784), .Y(n2687) );
  OAI21X1 U494 ( .A(n1832), .B(n1783), .C(n2686), .Y(n2171) );
  NAND2X1 U495 ( .A(\mem<19><12> ), .B(n1784), .Y(n2686) );
  OAI21X1 U496 ( .A(n1830), .B(n1783), .C(n2685), .Y(n2170) );
  NAND2X1 U497 ( .A(\mem<19><13> ), .B(n1784), .Y(n2685) );
  OAI21X1 U498 ( .A(n1828), .B(n1783), .C(n2684), .Y(n2169) );
  NAND2X1 U499 ( .A(\mem<19><14> ), .B(n1784), .Y(n2684) );
  OAI21X1 U500 ( .A(n1826), .B(n1783), .C(n2683), .Y(n2168) );
  NAND2X1 U501 ( .A(\mem<19><15> ), .B(n1784), .Y(n2683) );
  OAI21X1 U504 ( .A(n1851), .B(n1780), .C(n2682), .Y(n2167) );
  NAND2X1 U505 ( .A(\mem<18><0> ), .B(n1782), .Y(n2682) );
  OAI21X1 U506 ( .A(n1850), .B(n1780), .C(n2681), .Y(n2166) );
  NAND2X1 U507 ( .A(\mem<18><1> ), .B(n1782), .Y(n2681) );
  OAI21X1 U508 ( .A(n1848), .B(n1780), .C(n2680), .Y(n2165) );
  NAND2X1 U509 ( .A(\mem<18><2> ), .B(n1782), .Y(n2680) );
  OAI21X1 U510 ( .A(n1846), .B(n1780), .C(n2679), .Y(n2164) );
  NAND2X1 U511 ( .A(\mem<18><3> ), .B(n1782), .Y(n2679) );
  OAI21X1 U512 ( .A(n1845), .B(n1780), .C(n2678), .Y(n2163) );
  NAND2X1 U513 ( .A(\mem<18><4> ), .B(n1782), .Y(n2678) );
  OAI21X1 U514 ( .A(n1844), .B(n1780), .C(n2677), .Y(n2162) );
  NAND2X1 U515 ( .A(\mem<18><5> ), .B(n1782), .Y(n2677) );
  OAI21X1 U516 ( .A(n1842), .B(n1780), .C(n2676), .Y(n2161) );
  NAND2X1 U517 ( .A(\mem<18><6> ), .B(n1782), .Y(n2676) );
  OAI21X1 U518 ( .A(n1840), .B(n1780), .C(n2675), .Y(n2160) );
  NAND2X1 U519 ( .A(\mem<18><7> ), .B(n1782), .Y(n2675) );
  OAI21X1 U520 ( .A(n1839), .B(n1780), .C(n2674), .Y(n2159) );
  NAND2X1 U521 ( .A(\mem<18><8> ), .B(n1781), .Y(n2674) );
  OAI21X1 U522 ( .A(n1838), .B(n1780), .C(n2673), .Y(n2158) );
  NAND2X1 U523 ( .A(\mem<18><9> ), .B(n1781), .Y(n2673) );
  OAI21X1 U524 ( .A(n1836), .B(n1780), .C(n2672), .Y(n2157) );
  NAND2X1 U525 ( .A(\mem<18><10> ), .B(n1781), .Y(n2672) );
  OAI21X1 U526 ( .A(n1834), .B(n1780), .C(n2671), .Y(n2156) );
  NAND2X1 U527 ( .A(\mem<18><11> ), .B(n1781), .Y(n2671) );
  OAI21X1 U528 ( .A(n1833), .B(n1780), .C(n2670), .Y(n2155) );
  NAND2X1 U529 ( .A(\mem<18><12> ), .B(n1781), .Y(n2670) );
  OAI21X1 U530 ( .A(n1831), .B(n1780), .C(n2669), .Y(n2154) );
  NAND2X1 U531 ( .A(\mem<18><13> ), .B(n1781), .Y(n2669) );
  OAI21X1 U532 ( .A(n1829), .B(n1780), .C(n2668), .Y(n2153) );
  NAND2X1 U533 ( .A(\mem<18><14> ), .B(n1781), .Y(n2668) );
  OAI21X1 U534 ( .A(n1827), .B(n1780), .C(n2667), .Y(n2152) );
  NAND2X1 U535 ( .A(\mem<18><15> ), .B(n1781), .Y(n2667) );
  OAI21X1 U538 ( .A(n1851), .B(n1777), .C(n2666), .Y(n2151) );
  NAND2X1 U539 ( .A(\mem<17><0> ), .B(n1779), .Y(n2666) );
  OAI21X1 U540 ( .A(n1850), .B(n1777), .C(n2665), .Y(n2150) );
  NAND2X1 U541 ( .A(\mem<17><1> ), .B(n1779), .Y(n2665) );
  OAI21X1 U542 ( .A(n1848), .B(n1777), .C(n2664), .Y(n2149) );
  NAND2X1 U543 ( .A(\mem<17><2> ), .B(n1779), .Y(n2664) );
  OAI21X1 U544 ( .A(n1846), .B(n1777), .C(n2663), .Y(n2148) );
  NAND2X1 U545 ( .A(\mem<17><3> ), .B(n1779), .Y(n2663) );
  OAI21X1 U546 ( .A(n1845), .B(n1777), .C(n2662), .Y(n2147) );
  NAND2X1 U547 ( .A(\mem<17><4> ), .B(n1779), .Y(n2662) );
  OAI21X1 U548 ( .A(n1844), .B(n1777), .C(n2661), .Y(n2146) );
  NAND2X1 U549 ( .A(\mem<17><5> ), .B(n1779), .Y(n2661) );
  OAI21X1 U550 ( .A(n1842), .B(n1777), .C(n2660), .Y(n2145) );
  NAND2X1 U551 ( .A(\mem<17><6> ), .B(n1779), .Y(n2660) );
  OAI21X1 U552 ( .A(n1840), .B(n1777), .C(n2659), .Y(n2144) );
  NAND2X1 U553 ( .A(\mem<17><7> ), .B(n1779), .Y(n2659) );
  OAI21X1 U554 ( .A(n1839), .B(n1777), .C(n2658), .Y(n2143) );
  NAND2X1 U555 ( .A(\mem<17><8> ), .B(n1778), .Y(n2658) );
  OAI21X1 U556 ( .A(n1838), .B(n1777), .C(n2657), .Y(n2142) );
  NAND2X1 U557 ( .A(\mem<17><9> ), .B(n1778), .Y(n2657) );
  OAI21X1 U558 ( .A(n1836), .B(n1777), .C(n2656), .Y(n2141) );
  NAND2X1 U559 ( .A(\mem<17><10> ), .B(n1778), .Y(n2656) );
  OAI21X1 U560 ( .A(n1834), .B(n1777), .C(n2655), .Y(n2140) );
  NAND2X1 U561 ( .A(\mem<17><11> ), .B(n1778), .Y(n2655) );
  OAI21X1 U562 ( .A(n1833), .B(n1777), .C(n2654), .Y(n2139) );
  NAND2X1 U563 ( .A(\mem<17><12> ), .B(n1778), .Y(n2654) );
  OAI21X1 U564 ( .A(n1831), .B(n1777), .C(n2653), .Y(n2138) );
  NAND2X1 U565 ( .A(\mem<17><13> ), .B(n1778), .Y(n2653) );
  OAI21X1 U566 ( .A(n1829), .B(n1777), .C(n2652), .Y(n2137) );
  NAND2X1 U567 ( .A(\mem<17><14> ), .B(n1778), .Y(n2652) );
  OAI21X1 U568 ( .A(n1827), .B(n1777), .C(n2651), .Y(n2136) );
  NAND2X1 U569 ( .A(\mem<17><15> ), .B(n1778), .Y(n2651) );
  OAI21X1 U572 ( .A(n1851), .B(n1774), .C(n2650), .Y(n2135) );
  NAND2X1 U573 ( .A(\mem<16><0> ), .B(n1776), .Y(n2650) );
  OAI21X1 U574 ( .A(n1850), .B(n1774), .C(n2649), .Y(n2134) );
  NAND2X1 U575 ( .A(\mem<16><1> ), .B(n1776), .Y(n2649) );
  OAI21X1 U576 ( .A(n1848), .B(n1774), .C(n2648), .Y(n2133) );
  NAND2X1 U577 ( .A(\mem<16><2> ), .B(n1776), .Y(n2648) );
  OAI21X1 U578 ( .A(n1846), .B(n1774), .C(n2647), .Y(n2132) );
  NAND2X1 U579 ( .A(\mem<16><3> ), .B(n1776), .Y(n2647) );
  OAI21X1 U580 ( .A(n1845), .B(n1774), .C(n2646), .Y(n2131) );
  NAND2X1 U581 ( .A(\mem<16><4> ), .B(n1776), .Y(n2646) );
  OAI21X1 U582 ( .A(n1844), .B(n1774), .C(n2645), .Y(n2130) );
  NAND2X1 U583 ( .A(\mem<16><5> ), .B(n1776), .Y(n2645) );
  OAI21X1 U584 ( .A(n1842), .B(n1774), .C(n2644), .Y(n2129) );
  NAND2X1 U585 ( .A(\mem<16><6> ), .B(n1776), .Y(n2644) );
  OAI21X1 U586 ( .A(n1840), .B(n1774), .C(n2643), .Y(n2128) );
  NAND2X1 U587 ( .A(\mem<16><7> ), .B(n1776), .Y(n2643) );
  OAI21X1 U588 ( .A(n1839), .B(n1774), .C(n2642), .Y(n2127) );
  NAND2X1 U589 ( .A(\mem<16><8> ), .B(n1775), .Y(n2642) );
  OAI21X1 U590 ( .A(n1838), .B(n1774), .C(n2641), .Y(n2126) );
  NAND2X1 U591 ( .A(\mem<16><9> ), .B(n1775), .Y(n2641) );
  OAI21X1 U592 ( .A(n1836), .B(n1774), .C(n2640), .Y(n2125) );
  NAND2X1 U593 ( .A(\mem<16><10> ), .B(n1775), .Y(n2640) );
  OAI21X1 U594 ( .A(n1834), .B(n1774), .C(n2639), .Y(n2124) );
  NAND2X1 U595 ( .A(\mem<16><11> ), .B(n1775), .Y(n2639) );
  OAI21X1 U596 ( .A(n1833), .B(n1774), .C(n2638), .Y(n2123) );
  NAND2X1 U597 ( .A(\mem<16><12> ), .B(n1775), .Y(n2638) );
  OAI21X1 U598 ( .A(n1831), .B(n1774), .C(n2637), .Y(n2122) );
  NAND2X1 U599 ( .A(\mem<16><13> ), .B(n1775), .Y(n2637) );
  OAI21X1 U600 ( .A(n1829), .B(n1774), .C(n2636), .Y(n2121) );
  NAND2X1 U601 ( .A(\mem<16><14> ), .B(n1775), .Y(n2636) );
  OAI21X1 U602 ( .A(n1827), .B(n1774), .C(n2635), .Y(n2120) );
  NAND2X1 U603 ( .A(\mem<16><15> ), .B(n1775), .Y(n2635) );
  NAND3X1 U606 ( .A(n2763), .B(n1856), .C(n1857), .Y(n2634) );
  OAI21X1 U607 ( .A(n1851), .B(n1771), .C(n2633), .Y(n2119) );
  NAND2X1 U608 ( .A(\mem<15><0> ), .B(n1773), .Y(n2633) );
  OAI21X1 U609 ( .A(n1850), .B(n1771), .C(n2632), .Y(n2118) );
  NAND2X1 U610 ( .A(\mem<15><1> ), .B(n1773), .Y(n2632) );
  OAI21X1 U611 ( .A(n1848), .B(n1771), .C(n2631), .Y(n2117) );
  NAND2X1 U612 ( .A(\mem<15><2> ), .B(n1773), .Y(n2631) );
  OAI21X1 U613 ( .A(n1846), .B(n1771), .C(n2630), .Y(n2116) );
  NAND2X1 U614 ( .A(\mem<15><3> ), .B(n1773), .Y(n2630) );
  OAI21X1 U615 ( .A(n1845), .B(n1771), .C(n2629), .Y(n2115) );
  NAND2X1 U616 ( .A(\mem<15><4> ), .B(n1773), .Y(n2629) );
  OAI21X1 U617 ( .A(n1844), .B(n1771), .C(n2628), .Y(n2114) );
  NAND2X1 U618 ( .A(\mem<15><5> ), .B(n1773), .Y(n2628) );
  OAI21X1 U619 ( .A(n1842), .B(n1771), .C(n2627), .Y(n2113) );
  NAND2X1 U620 ( .A(\mem<15><6> ), .B(n1773), .Y(n2627) );
  OAI21X1 U621 ( .A(n1840), .B(n1771), .C(n2626), .Y(n2112) );
  NAND2X1 U622 ( .A(\mem<15><7> ), .B(n1773), .Y(n2626) );
  OAI21X1 U623 ( .A(n1839), .B(n1771), .C(n2625), .Y(n2111) );
  NAND2X1 U624 ( .A(\mem<15><8> ), .B(n1772), .Y(n2625) );
  OAI21X1 U625 ( .A(n1838), .B(n1771), .C(n2624), .Y(n2110) );
  NAND2X1 U626 ( .A(\mem<15><9> ), .B(n1772), .Y(n2624) );
  OAI21X1 U627 ( .A(n1836), .B(n1771), .C(n2623), .Y(n2109) );
  NAND2X1 U628 ( .A(\mem<15><10> ), .B(n1772), .Y(n2623) );
  OAI21X1 U629 ( .A(n1834), .B(n1771), .C(n2622), .Y(n2108) );
  NAND2X1 U630 ( .A(\mem<15><11> ), .B(n1772), .Y(n2622) );
  OAI21X1 U631 ( .A(n1833), .B(n1771), .C(n2621), .Y(n2107) );
  NAND2X1 U632 ( .A(\mem<15><12> ), .B(n1772), .Y(n2621) );
  OAI21X1 U633 ( .A(n1831), .B(n1771), .C(n2620), .Y(n2106) );
  NAND2X1 U634 ( .A(\mem<15><13> ), .B(n1772), .Y(n2620) );
  OAI21X1 U635 ( .A(n1829), .B(n1771), .C(n2619), .Y(n2105) );
  NAND2X1 U636 ( .A(\mem<15><14> ), .B(n1772), .Y(n2619) );
  OAI21X1 U637 ( .A(n1827), .B(n1771), .C(n2618), .Y(n2104) );
  NAND2X1 U638 ( .A(\mem<15><15> ), .B(n1772), .Y(n2618) );
  OAI21X1 U641 ( .A(n1851), .B(n1768), .C(n2617), .Y(n2103) );
  NAND2X1 U642 ( .A(\mem<14><0> ), .B(n1770), .Y(n2617) );
  OAI21X1 U643 ( .A(n1850), .B(n1768), .C(n2616), .Y(n2102) );
  NAND2X1 U644 ( .A(\mem<14><1> ), .B(n1770), .Y(n2616) );
  OAI21X1 U645 ( .A(n1848), .B(n1768), .C(n2615), .Y(n2101) );
  NAND2X1 U646 ( .A(\mem<14><2> ), .B(n1770), .Y(n2615) );
  OAI21X1 U647 ( .A(n1846), .B(n1768), .C(n2614), .Y(n2100) );
  NAND2X1 U648 ( .A(\mem<14><3> ), .B(n1770), .Y(n2614) );
  OAI21X1 U649 ( .A(n1845), .B(n1768), .C(n2613), .Y(n2099) );
  NAND2X1 U650 ( .A(\mem<14><4> ), .B(n1770), .Y(n2613) );
  OAI21X1 U651 ( .A(n1844), .B(n1768), .C(n2612), .Y(n2098) );
  NAND2X1 U652 ( .A(\mem<14><5> ), .B(n1770), .Y(n2612) );
  OAI21X1 U653 ( .A(n1842), .B(n1768), .C(n2611), .Y(n2097) );
  NAND2X1 U654 ( .A(\mem<14><6> ), .B(n1770), .Y(n2611) );
  OAI21X1 U655 ( .A(n1840), .B(n1768), .C(n2610), .Y(n2096) );
  NAND2X1 U656 ( .A(\mem<14><7> ), .B(n1770), .Y(n2610) );
  OAI21X1 U657 ( .A(n1839), .B(n1768), .C(n2609), .Y(n2095) );
  NAND2X1 U658 ( .A(\mem<14><8> ), .B(n1769), .Y(n2609) );
  OAI21X1 U659 ( .A(n1838), .B(n1768), .C(n2608), .Y(n2094) );
  NAND2X1 U660 ( .A(\mem<14><9> ), .B(n1769), .Y(n2608) );
  OAI21X1 U661 ( .A(n1836), .B(n1768), .C(n2607), .Y(n2093) );
  NAND2X1 U662 ( .A(\mem<14><10> ), .B(n1769), .Y(n2607) );
  OAI21X1 U663 ( .A(n1834), .B(n1768), .C(n2606), .Y(n2092) );
  NAND2X1 U664 ( .A(\mem<14><11> ), .B(n1769), .Y(n2606) );
  OAI21X1 U665 ( .A(n1833), .B(n1768), .C(n2605), .Y(n2091) );
  NAND2X1 U666 ( .A(\mem<14><12> ), .B(n1769), .Y(n2605) );
  OAI21X1 U667 ( .A(n1831), .B(n1768), .C(n2604), .Y(n2090) );
  NAND2X1 U668 ( .A(\mem<14><13> ), .B(n1769), .Y(n2604) );
  OAI21X1 U669 ( .A(n1829), .B(n1768), .C(n2603), .Y(n2089) );
  NAND2X1 U670 ( .A(\mem<14><14> ), .B(n1769), .Y(n2603) );
  OAI21X1 U671 ( .A(n1827), .B(n1768), .C(n2602), .Y(n2088) );
  NAND2X1 U672 ( .A(\mem<14><15> ), .B(n1769), .Y(n2602) );
  OAI21X1 U675 ( .A(n1851), .B(n1765), .C(n2601), .Y(n2087) );
  NAND2X1 U676 ( .A(\mem<13><0> ), .B(n1767), .Y(n2601) );
  OAI21X1 U677 ( .A(n1850), .B(n1765), .C(n2600), .Y(n2086) );
  NAND2X1 U678 ( .A(\mem<13><1> ), .B(n1767), .Y(n2600) );
  OAI21X1 U679 ( .A(n1848), .B(n1765), .C(n2599), .Y(n2085) );
  NAND2X1 U680 ( .A(\mem<13><2> ), .B(n1767), .Y(n2599) );
  OAI21X1 U681 ( .A(n1846), .B(n1765), .C(n2598), .Y(n2084) );
  NAND2X1 U682 ( .A(\mem<13><3> ), .B(n1767), .Y(n2598) );
  OAI21X1 U683 ( .A(n1845), .B(n1765), .C(n2597), .Y(n2083) );
  NAND2X1 U684 ( .A(\mem<13><4> ), .B(n1767), .Y(n2597) );
  OAI21X1 U685 ( .A(n1844), .B(n1765), .C(n2596), .Y(n2082) );
  NAND2X1 U686 ( .A(\mem<13><5> ), .B(n1767), .Y(n2596) );
  OAI21X1 U687 ( .A(n1842), .B(n1765), .C(n2595), .Y(n2081) );
  NAND2X1 U688 ( .A(\mem<13><6> ), .B(n1767), .Y(n2595) );
  OAI21X1 U689 ( .A(n1840), .B(n1765), .C(n2594), .Y(n2080) );
  NAND2X1 U690 ( .A(\mem<13><7> ), .B(n1767), .Y(n2594) );
  OAI21X1 U691 ( .A(n1839), .B(n1765), .C(n2593), .Y(n2079) );
  NAND2X1 U692 ( .A(\mem<13><8> ), .B(n1766), .Y(n2593) );
  OAI21X1 U693 ( .A(n1838), .B(n1765), .C(n2592), .Y(n2078) );
  NAND2X1 U694 ( .A(\mem<13><9> ), .B(n1766), .Y(n2592) );
  OAI21X1 U695 ( .A(n1836), .B(n1765), .C(n2591), .Y(n2077) );
  NAND2X1 U696 ( .A(\mem<13><10> ), .B(n1766), .Y(n2591) );
  OAI21X1 U697 ( .A(n1834), .B(n1765), .C(n2590), .Y(n2076) );
  NAND2X1 U698 ( .A(\mem<13><11> ), .B(n1766), .Y(n2590) );
  OAI21X1 U699 ( .A(n1833), .B(n1765), .C(n2589), .Y(n2075) );
  NAND2X1 U700 ( .A(\mem<13><12> ), .B(n1766), .Y(n2589) );
  OAI21X1 U701 ( .A(n1831), .B(n1765), .C(n2588), .Y(n2074) );
  NAND2X1 U702 ( .A(\mem<13><13> ), .B(n1766), .Y(n2588) );
  OAI21X1 U703 ( .A(n1829), .B(n1765), .C(n2587), .Y(n2073) );
  NAND2X1 U704 ( .A(\mem<13><14> ), .B(n1766), .Y(n2587) );
  OAI21X1 U705 ( .A(n1827), .B(n1765), .C(n2586), .Y(n2072) );
  NAND2X1 U706 ( .A(\mem<13><15> ), .B(n1766), .Y(n2586) );
  OAI21X1 U709 ( .A(n1851), .B(n1762), .C(n2585), .Y(n2071) );
  NAND2X1 U710 ( .A(\mem<12><0> ), .B(n1764), .Y(n2585) );
  OAI21X1 U711 ( .A(n1850), .B(n1762), .C(n2584), .Y(n2070) );
  NAND2X1 U712 ( .A(\mem<12><1> ), .B(n1764), .Y(n2584) );
  OAI21X1 U713 ( .A(n1848), .B(n1762), .C(n2583), .Y(n2069) );
  NAND2X1 U714 ( .A(\mem<12><2> ), .B(n1764), .Y(n2583) );
  OAI21X1 U715 ( .A(n1846), .B(n1762), .C(n2582), .Y(n2068) );
  NAND2X1 U716 ( .A(\mem<12><3> ), .B(n1764), .Y(n2582) );
  OAI21X1 U717 ( .A(n1845), .B(n1762), .C(n2581), .Y(n2067) );
  NAND2X1 U718 ( .A(\mem<12><4> ), .B(n1764), .Y(n2581) );
  OAI21X1 U719 ( .A(n1844), .B(n1762), .C(n2580), .Y(n2066) );
  NAND2X1 U720 ( .A(\mem<12><5> ), .B(n1764), .Y(n2580) );
  OAI21X1 U721 ( .A(n1842), .B(n1762), .C(n2579), .Y(n2065) );
  NAND2X1 U722 ( .A(\mem<12><6> ), .B(n1764), .Y(n2579) );
  OAI21X1 U723 ( .A(n1840), .B(n1762), .C(n2578), .Y(n2064) );
  NAND2X1 U724 ( .A(\mem<12><7> ), .B(n1764), .Y(n2578) );
  OAI21X1 U725 ( .A(n1839), .B(n1762), .C(n2577), .Y(n2063) );
  NAND2X1 U726 ( .A(\mem<12><8> ), .B(n1763), .Y(n2577) );
  OAI21X1 U727 ( .A(n1838), .B(n1762), .C(n2576), .Y(n2062) );
  NAND2X1 U728 ( .A(\mem<12><9> ), .B(n1763), .Y(n2576) );
  OAI21X1 U729 ( .A(n1836), .B(n1762), .C(n2575), .Y(n2061) );
  NAND2X1 U730 ( .A(\mem<12><10> ), .B(n1763), .Y(n2575) );
  OAI21X1 U731 ( .A(n1834), .B(n1762), .C(n2574), .Y(n2060) );
  NAND2X1 U732 ( .A(\mem<12><11> ), .B(n1763), .Y(n2574) );
  OAI21X1 U733 ( .A(n1833), .B(n1762), .C(n2573), .Y(n2059) );
  NAND2X1 U734 ( .A(\mem<12><12> ), .B(n1763), .Y(n2573) );
  OAI21X1 U735 ( .A(n1831), .B(n1762), .C(n2572), .Y(n2058) );
  NAND2X1 U736 ( .A(\mem<12><13> ), .B(n1763), .Y(n2572) );
  OAI21X1 U737 ( .A(n1829), .B(n1762), .C(n2571), .Y(n2057) );
  NAND2X1 U738 ( .A(\mem<12><14> ), .B(n1763), .Y(n2571) );
  OAI21X1 U739 ( .A(n1827), .B(n1762), .C(n2570), .Y(n2056) );
  NAND2X1 U740 ( .A(\mem<12><15> ), .B(n1763), .Y(n2570) );
  OAI21X1 U743 ( .A(n1851), .B(n1759), .C(n2569), .Y(n2055) );
  NAND2X1 U744 ( .A(\mem<11><0> ), .B(n1761), .Y(n2569) );
  OAI21X1 U745 ( .A(n1850), .B(n1759), .C(n2568), .Y(n2054) );
  NAND2X1 U746 ( .A(\mem<11><1> ), .B(n1761), .Y(n2568) );
  OAI21X1 U747 ( .A(n1848), .B(n1759), .C(n2567), .Y(n2053) );
  NAND2X1 U748 ( .A(\mem<11><2> ), .B(n1761), .Y(n2567) );
  OAI21X1 U749 ( .A(n1846), .B(n1759), .C(n2566), .Y(n2052) );
  NAND2X1 U750 ( .A(\mem<11><3> ), .B(n1761), .Y(n2566) );
  OAI21X1 U751 ( .A(n1845), .B(n1759), .C(n2565), .Y(n2051) );
  NAND2X1 U752 ( .A(\mem<11><4> ), .B(n1761), .Y(n2565) );
  OAI21X1 U753 ( .A(n1844), .B(n1759), .C(n2564), .Y(n2050) );
  NAND2X1 U754 ( .A(\mem<11><5> ), .B(n1761), .Y(n2564) );
  OAI21X1 U755 ( .A(n1842), .B(n1759), .C(n2563), .Y(n2049) );
  NAND2X1 U756 ( .A(\mem<11><6> ), .B(n1761), .Y(n2563) );
  OAI21X1 U757 ( .A(n1840), .B(n1759), .C(n2562), .Y(n2048) );
  NAND2X1 U758 ( .A(\mem<11><7> ), .B(n1761), .Y(n2562) );
  OAI21X1 U759 ( .A(n1839), .B(n1759), .C(n2561), .Y(n2047) );
  NAND2X1 U760 ( .A(\mem<11><8> ), .B(n1760), .Y(n2561) );
  OAI21X1 U761 ( .A(n1838), .B(n1759), .C(n2560), .Y(n2046) );
  NAND2X1 U762 ( .A(\mem<11><9> ), .B(n1760), .Y(n2560) );
  OAI21X1 U763 ( .A(n1836), .B(n1759), .C(n2559), .Y(n2045) );
  NAND2X1 U764 ( .A(\mem<11><10> ), .B(n1760), .Y(n2559) );
  OAI21X1 U765 ( .A(n1834), .B(n1759), .C(n2558), .Y(n2044) );
  NAND2X1 U766 ( .A(\mem<11><11> ), .B(n1760), .Y(n2558) );
  OAI21X1 U767 ( .A(n1833), .B(n1759), .C(n2557), .Y(n2043) );
  NAND2X1 U768 ( .A(\mem<11><12> ), .B(n1760), .Y(n2557) );
  OAI21X1 U769 ( .A(n1831), .B(n1759), .C(n2556), .Y(n2042) );
  NAND2X1 U770 ( .A(\mem<11><13> ), .B(n1760), .Y(n2556) );
  OAI21X1 U771 ( .A(n1829), .B(n1759), .C(n2555), .Y(n2041) );
  NAND2X1 U772 ( .A(\mem<11><14> ), .B(n1760), .Y(n2555) );
  OAI21X1 U773 ( .A(n1827), .B(n1759), .C(n2554), .Y(n2040) );
  NAND2X1 U774 ( .A(\mem<11><15> ), .B(n1760), .Y(n2554) );
  OAI21X1 U777 ( .A(n1851), .B(n1756), .C(n2553), .Y(n2039) );
  NAND2X1 U778 ( .A(\mem<10><0> ), .B(n1758), .Y(n2553) );
  OAI21X1 U779 ( .A(n1850), .B(n1756), .C(n2552), .Y(n2038) );
  NAND2X1 U780 ( .A(\mem<10><1> ), .B(n1758), .Y(n2552) );
  OAI21X1 U781 ( .A(n1848), .B(n1756), .C(n2551), .Y(n2037) );
  NAND2X1 U782 ( .A(\mem<10><2> ), .B(n1758), .Y(n2551) );
  OAI21X1 U783 ( .A(n1846), .B(n1756), .C(n2550), .Y(n2036) );
  NAND2X1 U784 ( .A(\mem<10><3> ), .B(n1758), .Y(n2550) );
  OAI21X1 U785 ( .A(n1845), .B(n1756), .C(n2549), .Y(n2035) );
  NAND2X1 U786 ( .A(\mem<10><4> ), .B(n1758), .Y(n2549) );
  OAI21X1 U787 ( .A(n1844), .B(n1756), .C(n2548), .Y(n2034) );
  NAND2X1 U788 ( .A(\mem<10><5> ), .B(n1758), .Y(n2548) );
  OAI21X1 U789 ( .A(n1842), .B(n1756), .C(n2547), .Y(n2033) );
  NAND2X1 U790 ( .A(\mem<10><6> ), .B(n1758), .Y(n2547) );
  OAI21X1 U791 ( .A(n1840), .B(n1756), .C(n2546), .Y(n2032) );
  NAND2X1 U792 ( .A(\mem<10><7> ), .B(n1758), .Y(n2546) );
  OAI21X1 U793 ( .A(n1839), .B(n1756), .C(n2545), .Y(n2031) );
  NAND2X1 U794 ( .A(\mem<10><8> ), .B(n1757), .Y(n2545) );
  OAI21X1 U795 ( .A(n1838), .B(n1756), .C(n2544), .Y(n2030) );
  NAND2X1 U796 ( .A(\mem<10><9> ), .B(n1757), .Y(n2544) );
  OAI21X1 U797 ( .A(n1836), .B(n1756), .C(n2543), .Y(n2029) );
  NAND2X1 U798 ( .A(\mem<10><10> ), .B(n1757), .Y(n2543) );
  OAI21X1 U799 ( .A(n1834), .B(n1756), .C(n2542), .Y(n2028) );
  NAND2X1 U800 ( .A(\mem<10><11> ), .B(n1757), .Y(n2542) );
  OAI21X1 U801 ( .A(n1833), .B(n1756), .C(n2541), .Y(n2027) );
  NAND2X1 U802 ( .A(\mem<10><12> ), .B(n1757), .Y(n2541) );
  OAI21X1 U803 ( .A(n1831), .B(n1756), .C(n2540), .Y(n2026) );
  NAND2X1 U804 ( .A(\mem<10><13> ), .B(n1757), .Y(n2540) );
  OAI21X1 U805 ( .A(n1829), .B(n1756), .C(n2539), .Y(n2025) );
  NAND2X1 U806 ( .A(\mem<10><14> ), .B(n1757), .Y(n2539) );
  OAI21X1 U807 ( .A(n1827), .B(n1756), .C(n2538), .Y(n2024) );
  NAND2X1 U808 ( .A(\mem<10><15> ), .B(n1757), .Y(n2538) );
  OAI21X1 U811 ( .A(n1851), .B(n1753), .C(n2537), .Y(n2023) );
  NAND2X1 U812 ( .A(\mem<9><0> ), .B(n1755), .Y(n2537) );
  OAI21X1 U813 ( .A(n1850), .B(n1753), .C(n2536), .Y(n2022) );
  NAND2X1 U814 ( .A(\mem<9><1> ), .B(n1755), .Y(n2536) );
  OAI21X1 U815 ( .A(n1848), .B(n1753), .C(n2535), .Y(n2021) );
  NAND2X1 U816 ( .A(\mem<9><2> ), .B(n1755), .Y(n2535) );
  OAI21X1 U817 ( .A(n1846), .B(n1753), .C(n2534), .Y(n2020) );
  NAND2X1 U818 ( .A(\mem<9><3> ), .B(n1755), .Y(n2534) );
  OAI21X1 U819 ( .A(n1845), .B(n1753), .C(n2533), .Y(n2019) );
  NAND2X1 U820 ( .A(\mem<9><4> ), .B(n1755), .Y(n2533) );
  OAI21X1 U821 ( .A(n1844), .B(n1753), .C(n2532), .Y(n2018) );
  NAND2X1 U822 ( .A(\mem<9><5> ), .B(n1755), .Y(n2532) );
  OAI21X1 U823 ( .A(n1842), .B(n1753), .C(n2531), .Y(n2017) );
  NAND2X1 U824 ( .A(\mem<9><6> ), .B(n1755), .Y(n2531) );
  OAI21X1 U825 ( .A(n1840), .B(n1753), .C(n2530), .Y(n2016) );
  NAND2X1 U826 ( .A(\mem<9><7> ), .B(n1755), .Y(n2530) );
  OAI21X1 U827 ( .A(n1839), .B(n1753), .C(n2529), .Y(n2015) );
  NAND2X1 U828 ( .A(\mem<9><8> ), .B(n1754), .Y(n2529) );
  OAI21X1 U829 ( .A(n1838), .B(n1753), .C(n2528), .Y(n2014) );
  NAND2X1 U830 ( .A(\mem<9><9> ), .B(n1754), .Y(n2528) );
  OAI21X1 U831 ( .A(n1836), .B(n1753), .C(n2527), .Y(n2013) );
  NAND2X1 U832 ( .A(\mem<9><10> ), .B(n1754), .Y(n2527) );
  OAI21X1 U833 ( .A(n1834), .B(n1753), .C(n2526), .Y(n2012) );
  NAND2X1 U834 ( .A(\mem<9><11> ), .B(n1754), .Y(n2526) );
  OAI21X1 U835 ( .A(n1833), .B(n1753), .C(n2525), .Y(n2011) );
  NAND2X1 U836 ( .A(\mem<9><12> ), .B(n1754), .Y(n2525) );
  OAI21X1 U837 ( .A(n1831), .B(n1753), .C(n2524), .Y(n2010) );
  NAND2X1 U838 ( .A(\mem<9><13> ), .B(n1754), .Y(n2524) );
  OAI21X1 U839 ( .A(n1829), .B(n1753), .C(n2523), .Y(n2009) );
  NAND2X1 U840 ( .A(\mem<9><14> ), .B(n1754), .Y(n2523) );
  OAI21X1 U841 ( .A(n1827), .B(n1753), .C(n2522), .Y(n2008) );
  NAND2X1 U842 ( .A(\mem<9><15> ), .B(n1754), .Y(n2522) );
  OAI21X1 U845 ( .A(n1851), .B(n1750), .C(n2521), .Y(n2007) );
  NAND2X1 U846 ( .A(\mem<8><0> ), .B(n1752), .Y(n2521) );
  OAI21X1 U847 ( .A(n1850), .B(n1750), .C(n2520), .Y(n2006) );
  NAND2X1 U848 ( .A(\mem<8><1> ), .B(n1752), .Y(n2520) );
  OAI21X1 U849 ( .A(n1848), .B(n1750), .C(n2519), .Y(n2005) );
  NAND2X1 U850 ( .A(\mem<8><2> ), .B(n1752), .Y(n2519) );
  OAI21X1 U851 ( .A(n1846), .B(n1750), .C(n2518), .Y(n2004) );
  NAND2X1 U852 ( .A(\mem<8><3> ), .B(n1752), .Y(n2518) );
  OAI21X1 U853 ( .A(n1845), .B(n1750), .C(n2517), .Y(n2003) );
  NAND2X1 U854 ( .A(\mem<8><4> ), .B(n1752), .Y(n2517) );
  OAI21X1 U855 ( .A(n1844), .B(n1750), .C(n2516), .Y(n2002) );
  NAND2X1 U856 ( .A(\mem<8><5> ), .B(n1752), .Y(n2516) );
  OAI21X1 U857 ( .A(n1842), .B(n1750), .C(n2515), .Y(n2001) );
  NAND2X1 U858 ( .A(\mem<8><6> ), .B(n1752), .Y(n2515) );
  OAI21X1 U859 ( .A(n1840), .B(n1750), .C(n2514), .Y(n2000) );
  NAND2X1 U860 ( .A(\mem<8><7> ), .B(n1752), .Y(n2514) );
  OAI21X1 U861 ( .A(n1839), .B(n1750), .C(n2513), .Y(n1999) );
  NAND2X1 U862 ( .A(\mem<8><8> ), .B(n1751), .Y(n2513) );
  OAI21X1 U863 ( .A(n1838), .B(n1750), .C(n2512), .Y(n1998) );
  NAND2X1 U864 ( .A(\mem<8><9> ), .B(n1751), .Y(n2512) );
  OAI21X1 U865 ( .A(n1836), .B(n1750), .C(n2511), .Y(n1997) );
  NAND2X1 U866 ( .A(\mem<8><10> ), .B(n1751), .Y(n2511) );
  OAI21X1 U867 ( .A(n1834), .B(n1750), .C(n2510), .Y(n1996) );
  NAND2X1 U868 ( .A(\mem<8><11> ), .B(n1751), .Y(n2510) );
  OAI21X1 U869 ( .A(n1833), .B(n1750), .C(n2509), .Y(n1995) );
  NAND2X1 U870 ( .A(\mem<8><12> ), .B(n1751), .Y(n2509) );
  OAI21X1 U871 ( .A(n1831), .B(n1750), .C(n2508), .Y(n1994) );
  NAND2X1 U872 ( .A(\mem<8><13> ), .B(n1751), .Y(n2508) );
  OAI21X1 U873 ( .A(n1829), .B(n1750), .C(n2507), .Y(n1993) );
  NAND2X1 U874 ( .A(\mem<8><14> ), .B(n1751), .Y(n2507) );
  OAI21X1 U875 ( .A(n1827), .B(n1750), .C(n2506), .Y(n1992) );
  NAND2X1 U876 ( .A(\mem<8><15> ), .B(n1751), .Y(n2506) );
  NAND3X1 U879 ( .A(n2763), .B(n1858), .C(n1855), .Y(n2505) );
  OAI21X1 U880 ( .A(n1851), .B(n1747), .C(n2504), .Y(n1991) );
  NAND2X1 U881 ( .A(\mem<7><0> ), .B(n1749), .Y(n2504) );
  OAI21X1 U882 ( .A(n1850), .B(n1747), .C(n2503), .Y(n1990) );
  NAND2X1 U883 ( .A(\mem<7><1> ), .B(n1749), .Y(n2503) );
  OAI21X1 U884 ( .A(n1848), .B(n1747), .C(n2502), .Y(n1989) );
  NAND2X1 U885 ( .A(\mem<7><2> ), .B(n1749), .Y(n2502) );
  OAI21X1 U886 ( .A(n1846), .B(n1747), .C(n2501), .Y(n1988) );
  NAND2X1 U887 ( .A(\mem<7><3> ), .B(n1749), .Y(n2501) );
  OAI21X1 U888 ( .A(n1845), .B(n1747), .C(n2500), .Y(n1987) );
  NAND2X1 U889 ( .A(\mem<7><4> ), .B(n1749), .Y(n2500) );
  OAI21X1 U890 ( .A(n1844), .B(n1747), .C(n2499), .Y(n1986) );
  NAND2X1 U891 ( .A(\mem<7><5> ), .B(n1749), .Y(n2499) );
  OAI21X1 U892 ( .A(n1842), .B(n1747), .C(n2498), .Y(n1985) );
  NAND2X1 U893 ( .A(\mem<7><6> ), .B(n1749), .Y(n2498) );
  OAI21X1 U894 ( .A(n1840), .B(n1747), .C(n2497), .Y(n1984) );
  NAND2X1 U895 ( .A(\mem<7><7> ), .B(n1749), .Y(n2497) );
  OAI21X1 U896 ( .A(n1839), .B(n1747), .C(n2496), .Y(n1983) );
  NAND2X1 U897 ( .A(\mem<7><8> ), .B(n1748), .Y(n2496) );
  OAI21X1 U898 ( .A(n1838), .B(n1747), .C(n2495), .Y(n1982) );
  NAND2X1 U899 ( .A(\mem<7><9> ), .B(n1748), .Y(n2495) );
  OAI21X1 U900 ( .A(n1836), .B(n1747), .C(n2494), .Y(n1981) );
  NAND2X1 U901 ( .A(\mem<7><10> ), .B(n1748), .Y(n2494) );
  OAI21X1 U902 ( .A(n1834), .B(n1747), .C(n2493), .Y(n1980) );
  NAND2X1 U903 ( .A(\mem<7><11> ), .B(n1748), .Y(n2493) );
  OAI21X1 U904 ( .A(n1833), .B(n1747), .C(n2492), .Y(n1979) );
  NAND2X1 U905 ( .A(\mem<7><12> ), .B(n1748), .Y(n2492) );
  OAI21X1 U906 ( .A(n1831), .B(n1747), .C(n2491), .Y(n1978) );
  NAND2X1 U907 ( .A(\mem<7><13> ), .B(n1748), .Y(n2491) );
  OAI21X1 U908 ( .A(n1829), .B(n1747), .C(n2490), .Y(n1977) );
  NAND2X1 U909 ( .A(\mem<7><14> ), .B(n1748), .Y(n2490) );
  OAI21X1 U910 ( .A(n1827), .B(n1747), .C(n2489), .Y(n1976) );
  NAND2X1 U911 ( .A(\mem<7><15> ), .B(n1748), .Y(n2489) );
  NOR3X1 U914 ( .A(n1853), .B(n1710), .C(n1854), .Y(n2884) );
  OAI21X1 U915 ( .A(n1851), .B(n1744), .C(n2488), .Y(n1975) );
  NAND2X1 U916 ( .A(\mem<6><0> ), .B(n1746), .Y(n2488) );
  OAI21X1 U917 ( .A(n1850), .B(n1744), .C(n2487), .Y(n1974) );
  NAND2X1 U918 ( .A(\mem<6><1> ), .B(n1746), .Y(n2487) );
  OAI21X1 U919 ( .A(n1848), .B(n1744), .C(n2486), .Y(n1973) );
  NAND2X1 U920 ( .A(\mem<6><2> ), .B(n1746), .Y(n2486) );
  OAI21X1 U921 ( .A(n1846), .B(n1744), .C(n2485), .Y(n1972) );
  NAND2X1 U922 ( .A(\mem<6><3> ), .B(n1746), .Y(n2485) );
  OAI21X1 U923 ( .A(n1845), .B(n1744), .C(n2484), .Y(n1971) );
  NAND2X1 U924 ( .A(\mem<6><4> ), .B(n1746), .Y(n2484) );
  OAI21X1 U925 ( .A(n1844), .B(n1744), .C(n2483), .Y(n1970) );
  NAND2X1 U926 ( .A(\mem<6><5> ), .B(n1746), .Y(n2483) );
  OAI21X1 U927 ( .A(n1842), .B(n1744), .C(n2482), .Y(n1969) );
  NAND2X1 U928 ( .A(\mem<6><6> ), .B(n1746), .Y(n2482) );
  OAI21X1 U929 ( .A(n1840), .B(n1744), .C(n2481), .Y(n1968) );
  NAND2X1 U930 ( .A(\mem<6><7> ), .B(n1746), .Y(n2481) );
  OAI21X1 U931 ( .A(n1839), .B(n1744), .C(n2480), .Y(n1967) );
  NAND2X1 U932 ( .A(\mem<6><8> ), .B(n1745), .Y(n2480) );
  OAI21X1 U933 ( .A(n1838), .B(n1744), .C(n2479), .Y(n1966) );
  NAND2X1 U934 ( .A(\mem<6><9> ), .B(n1745), .Y(n2479) );
  OAI21X1 U935 ( .A(n1836), .B(n1744), .C(n2478), .Y(n1965) );
  NAND2X1 U936 ( .A(\mem<6><10> ), .B(n1745), .Y(n2478) );
  OAI21X1 U937 ( .A(n1834), .B(n1744), .C(n2477), .Y(n1964) );
  NAND2X1 U938 ( .A(\mem<6><11> ), .B(n1745), .Y(n2477) );
  OAI21X1 U939 ( .A(n1833), .B(n1744), .C(n2476), .Y(n1963) );
  NAND2X1 U940 ( .A(\mem<6><12> ), .B(n1745), .Y(n2476) );
  OAI21X1 U941 ( .A(n1831), .B(n1744), .C(n2475), .Y(n1962) );
  NAND2X1 U942 ( .A(\mem<6><13> ), .B(n1745), .Y(n2475) );
  OAI21X1 U943 ( .A(n1829), .B(n1744), .C(n2474), .Y(n1961) );
  NAND2X1 U944 ( .A(\mem<6><14> ), .B(n1745), .Y(n2474) );
  OAI21X1 U945 ( .A(n1827), .B(n1744), .C(n2473), .Y(n1960) );
  NAND2X1 U946 ( .A(\mem<6><15> ), .B(n1745), .Y(n2473) );
  NOR3X1 U949 ( .A(n1853), .B(n1723), .C(n1854), .Y(n2867) );
  OAI21X1 U950 ( .A(n1851), .B(n1741), .C(n2472), .Y(n1959) );
  NAND2X1 U951 ( .A(\mem<5><0> ), .B(n1743), .Y(n2472) );
  OAI21X1 U952 ( .A(n1849), .B(n1741), .C(n2471), .Y(n1958) );
  NAND2X1 U953 ( .A(\mem<5><1> ), .B(n1743), .Y(n2471) );
  OAI21X1 U954 ( .A(n1847), .B(n1741), .C(n2470), .Y(n1957) );
  NAND2X1 U955 ( .A(\mem<5><2> ), .B(n1743), .Y(n2470) );
  OAI21X1 U956 ( .A(n1846), .B(n1741), .C(n2469), .Y(n1956) );
  NAND2X1 U957 ( .A(\mem<5><3> ), .B(n1743), .Y(n2469) );
  OAI21X1 U958 ( .A(n1845), .B(n1741), .C(n2468), .Y(n1955) );
  NAND2X1 U959 ( .A(\mem<5><4> ), .B(n1743), .Y(n2468) );
  OAI21X1 U960 ( .A(n1843), .B(n1741), .C(n2467), .Y(n1954) );
  NAND2X1 U961 ( .A(\mem<5><5> ), .B(n1743), .Y(n2467) );
  OAI21X1 U962 ( .A(n1841), .B(n1741), .C(n2466), .Y(n1953) );
  NAND2X1 U963 ( .A(\mem<5><6> ), .B(n1743), .Y(n2466) );
  OAI21X1 U964 ( .A(n1840), .B(n1741), .C(n2465), .Y(n1952) );
  NAND2X1 U965 ( .A(\mem<5><7> ), .B(n1743), .Y(n2465) );
  OAI21X1 U966 ( .A(n1839), .B(n1741), .C(n2464), .Y(n1951) );
  NAND2X1 U967 ( .A(\mem<5><8> ), .B(n1742), .Y(n2464) );
  OAI21X1 U968 ( .A(n1837), .B(n1741), .C(n2463), .Y(n1950) );
  NAND2X1 U969 ( .A(\mem<5><9> ), .B(n1742), .Y(n2463) );
  OAI21X1 U970 ( .A(n1835), .B(n1741), .C(n2462), .Y(n1949) );
  NAND2X1 U971 ( .A(\mem<5><10> ), .B(n1742), .Y(n2462) );
  OAI21X1 U972 ( .A(n1834), .B(n1741), .C(n2461), .Y(n1948) );
  NAND2X1 U973 ( .A(\mem<5><11> ), .B(n1742), .Y(n2461) );
  OAI21X1 U974 ( .A(n1832), .B(n1741), .C(n2460), .Y(n1947) );
  NAND2X1 U975 ( .A(\mem<5><12> ), .B(n1742), .Y(n2460) );
  OAI21X1 U976 ( .A(n1830), .B(n1741), .C(n2459), .Y(n1946) );
  NAND2X1 U977 ( .A(\mem<5><13> ), .B(n1742), .Y(n2459) );
  OAI21X1 U978 ( .A(n1828), .B(n1741), .C(n2458), .Y(n1945) );
  NAND2X1 U979 ( .A(\mem<5><14> ), .B(n1742), .Y(n2458) );
  OAI21X1 U980 ( .A(n1826), .B(n1741), .C(n2457), .Y(n1944) );
  NAND2X1 U981 ( .A(\mem<5><15> ), .B(n1742), .Y(n2457) );
  NOR3X1 U984 ( .A(n1711), .B(n1852), .C(n1854), .Y(n2850) );
  OAI21X1 U985 ( .A(n1851), .B(n1738), .C(n2456), .Y(n1943) );
  NAND2X1 U986 ( .A(\mem<4><0> ), .B(n1740), .Y(n2456) );
  OAI21X1 U987 ( .A(n1850), .B(n1738), .C(n2455), .Y(n1942) );
  NAND2X1 U988 ( .A(\mem<4><1> ), .B(n1740), .Y(n2455) );
  OAI21X1 U989 ( .A(n1848), .B(n1738), .C(n2454), .Y(n1941) );
  NAND2X1 U990 ( .A(\mem<4><2> ), .B(n1740), .Y(n2454) );
  OAI21X1 U991 ( .A(n1846), .B(n1738), .C(n2453), .Y(n1940) );
  NAND2X1 U992 ( .A(\mem<4><3> ), .B(n1740), .Y(n2453) );
  OAI21X1 U993 ( .A(n1845), .B(n1738), .C(n2452), .Y(n1939) );
  NAND2X1 U994 ( .A(\mem<4><4> ), .B(n1740), .Y(n2452) );
  OAI21X1 U995 ( .A(n1844), .B(n1738), .C(n2451), .Y(n1938) );
  NAND2X1 U996 ( .A(\mem<4><5> ), .B(n1740), .Y(n2451) );
  OAI21X1 U997 ( .A(n1842), .B(n1738), .C(n2450), .Y(n1937) );
  NAND2X1 U998 ( .A(\mem<4><6> ), .B(n1740), .Y(n2450) );
  OAI21X1 U999 ( .A(n1840), .B(n1738), .C(n2449), .Y(n1936) );
  NAND2X1 U1000 ( .A(\mem<4><7> ), .B(n1740), .Y(n2449) );
  OAI21X1 U1001 ( .A(n1839), .B(n1738), .C(n2448), .Y(n1935) );
  NAND2X1 U1002 ( .A(\mem<4><8> ), .B(n1739), .Y(n2448) );
  OAI21X1 U1003 ( .A(n1838), .B(n1738), .C(n2447), .Y(n1934) );
  NAND2X1 U1004 ( .A(\mem<4><9> ), .B(n1739), .Y(n2447) );
  OAI21X1 U1005 ( .A(n1836), .B(n1738), .C(n2446), .Y(n1933) );
  NAND2X1 U1006 ( .A(\mem<4><10> ), .B(n1739), .Y(n2446) );
  OAI21X1 U1007 ( .A(n1834), .B(n1738), .C(n2445), .Y(n1932) );
  NAND2X1 U1008 ( .A(\mem<4><11> ), .B(n1739), .Y(n2445) );
  OAI21X1 U1009 ( .A(n1833), .B(n1738), .C(n2444), .Y(n1931) );
  NAND2X1 U1010 ( .A(\mem<4><12> ), .B(n1739), .Y(n2444) );
  OAI21X1 U1011 ( .A(n1831), .B(n1738), .C(n2443), .Y(n1930) );
  NAND2X1 U1012 ( .A(\mem<4><13> ), .B(n1739), .Y(n2443) );
  OAI21X1 U1013 ( .A(n1829), .B(n1738), .C(n2442), .Y(n1929) );
  NAND2X1 U1014 ( .A(\mem<4><14> ), .B(n1739), .Y(n2442) );
  OAI21X1 U1015 ( .A(n1827), .B(n1738), .C(n2441), .Y(n1928) );
  NAND2X1 U1016 ( .A(\mem<4><15> ), .B(n1739), .Y(n2441) );
  NOR3X1 U1019 ( .A(n1723), .B(n1852), .C(n1854), .Y(n2833) );
  OAI21X1 U1020 ( .A(n1851), .B(n1735), .C(n2440), .Y(n1927) );
  NAND2X1 U1021 ( .A(\mem<3><0> ), .B(n1737), .Y(n2440) );
  OAI21X1 U1022 ( .A(n1849), .B(n1735), .C(n2439), .Y(n1926) );
  NAND2X1 U1023 ( .A(\mem<3><1> ), .B(n1737), .Y(n2439) );
  OAI21X1 U1024 ( .A(n1847), .B(n1735), .C(n2438), .Y(n1925) );
  NAND2X1 U1025 ( .A(\mem<3><2> ), .B(n1737), .Y(n2438) );
  OAI21X1 U1026 ( .A(n1846), .B(n1735), .C(n2437), .Y(n1924) );
  NAND2X1 U1027 ( .A(\mem<3><3> ), .B(n1737), .Y(n2437) );
  OAI21X1 U1028 ( .A(n1845), .B(n1735), .C(n2436), .Y(n1923) );
  NAND2X1 U1029 ( .A(\mem<3><4> ), .B(n1737), .Y(n2436) );
  OAI21X1 U1030 ( .A(n1843), .B(n1735), .C(n2435), .Y(n1922) );
  NAND2X1 U1031 ( .A(\mem<3><5> ), .B(n1737), .Y(n2435) );
  OAI21X1 U1032 ( .A(n1841), .B(n1735), .C(n2434), .Y(n1921) );
  NAND2X1 U1033 ( .A(\mem<3><6> ), .B(n1737), .Y(n2434) );
  OAI21X1 U1034 ( .A(n1840), .B(n1735), .C(n2433), .Y(n1920) );
  NAND2X1 U1035 ( .A(\mem<3><7> ), .B(n1737), .Y(n2433) );
  OAI21X1 U1036 ( .A(n1839), .B(n1735), .C(n2432), .Y(n1919) );
  NAND2X1 U1037 ( .A(\mem<3><8> ), .B(n1736), .Y(n2432) );
  OAI21X1 U1038 ( .A(n1837), .B(n1735), .C(n2431), .Y(n1918) );
  NAND2X1 U1039 ( .A(\mem<3><9> ), .B(n1736), .Y(n2431) );
  OAI21X1 U1040 ( .A(n1835), .B(n1735), .C(n2430), .Y(n1917) );
  NAND2X1 U1041 ( .A(\mem<3><10> ), .B(n1736), .Y(n2430) );
  OAI21X1 U1042 ( .A(n1834), .B(n1735), .C(n2429), .Y(n1916) );
  NAND2X1 U1043 ( .A(\mem<3><11> ), .B(n1736), .Y(n2429) );
  OAI21X1 U1044 ( .A(n1832), .B(n1735), .C(n2428), .Y(n1915) );
  NAND2X1 U1045 ( .A(\mem<3><12> ), .B(n1736), .Y(n2428) );
  OAI21X1 U1046 ( .A(n1830), .B(n1735), .C(n2427), .Y(n1914) );
  NAND2X1 U1047 ( .A(\mem<3><13> ), .B(n1736), .Y(n2427) );
  OAI21X1 U1048 ( .A(n1828), .B(n1735), .C(n2426), .Y(n1913) );
  NAND2X1 U1049 ( .A(\mem<3><14> ), .B(n1736), .Y(n2426) );
  OAI21X1 U1050 ( .A(n1826), .B(n1735), .C(n2425), .Y(n1912) );
  NAND2X1 U1051 ( .A(\mem<3><15> ), .B(n1736), .Y(n2425) );
  NOR3X1 U1054 ( .A(n1711), .B(n1691), .C(n1853), .Y(n2816) );
  OAI21X1 U1055 ( .A(n1851), .B(n1732), .C(n2424), .Y(n1911) );
  NAND2X1 U1056 ( .A(\mem<2><0> ), .B(n1734), .Y(n2424) );
  OAI21X1 U1057 ( .A(n1850), .B(n1732), .C(n2423), .Y(n1910) );
  NAND2X1 U1058 ( .A(\mem<2><1> ), .B(n1734), .Y(n2423) );
  OAI21X1 U1059 ( .A(n1848), .B(n1732), .C(n2422), .Y(n1909) );
  NAND2X1 U1060 ( .A(\mem<2><2> ), .B(n1734), .Y(n2422) );
  OAI21X1 U1061 ( .A(n1846), .B(n1732), .C(n2421), .Y(n1908) );
  NAND2X1 U1062 ( .A(\mem<2><3> ), .B(n1734), .Y(n2421) );
  OAI21X1 U1063 ( .A(n1845), .B(n1732), .C(n2420), .Y(n1907) );
  NAND2X1 U1064 ( .A(\mem<2><4> ), .B(n1734), .Y(n2420) );
  OAI21X1 U1065 ( .A(n1844), .B(n1732), .C(n2419), .Y(n1906) );
  NAND2X1 U1066 ( .A(\mem<2><5> ), .B(n1734), .Y(n2419) );
  OAI21X1 U1067 ( .A(n1842), .B(n1732), .C(n2418), .Y(n1905) );
  NAND2X1 U1068 ( .A(\mem<2><6> ), .B(n1734), .Y(n2418) );
  OAI21X1 U1069 ( .A(n1840), .B(n1732), .C(n2417), .Y(n1904) );
  NAND2X1 U1070 ( .A(\mem<2><7> ), .B(n1734), .Y(n2417) );
  OAI21X1 U1071 ( .A(n1839), .B(n1732), .C(n2416), .Y(n1903) );
  NAND2X1 U1072 ( .A(\mem<2><8> ), .B(n1733), .Y(n2416) );
  OAI21X1 U1073 ( .A(n1838), .B(n1732), .C(n2415), .Y(n1902) );
  NAND2X1 U1074 ( .A(\mem<2><9> ), .B(n1733), .Y(n2415) );
  OAI21X1 U1075 ( .A(n1836), .B(n1732), .C(n2414), .Y(n1901) );
  NAND2X1 U1076 ( .A(\mem<2><10> ), .B(n1733), .Y(n2414) );
  OAI21X1 U1077 ( .A(n1834), .B(n1732), .C(n2413), .Y(n1900) );
  NAND2X1 U1078 ( .A(\mem<2><11> ), .B(n1733), .Y(n2413) );
  OAI21X1 U1079 ( .A(n1833), .B(n1732), .C(n2412), .Y(n1899) );
  NAND2X1 U1080 ( .A(\mem<2><12> ), .B(n1733), .Y(n2412) );
  OAI21X1 U1081 ( .A(n1831), .B(n1732), .C(n2411), .Y(n1898) );
  NAND2X1 U1082 ( .A(\mem<2><13> ), .B(n1733), .Y(n2411) );
  OAI21X1 U1083 ( .A(n1829), .B(n1732), .C(n2410), .Y(n1897) );
  NAND2X1 U1084 ( .A(\mem<2><14> ), .B(n1733), .Y(n2410) );
  OAI21X1 U1085 ( .A(n1827), .B(n1732), .C(n2409), .Y(n1896) );
  NAND2X1 U1086 ( .A(\mem<2><15> ), .B(n1733), .Y(n2409) );
  NOR3X1 U1089 ( .A(n1722), .B(n1691), .C(n1853), .Y(n2799) );
  OAI21X1 U1090 ( .A(n1851), .B(n1729), .C(n2408), .Y(n1895) );
  NAND2X1 U1091 ( .A(\mem<1><0> ), .B(n1731), .Y(n2408) );
  OAI21X1 U1092 ( .A(n1849), .B(n1729), .C(n2407), .Y(n1894) );
  NAND2X1 U1093 ( .A(\mem<1><1> ), .B(n1731), .Y(n2407) );
  OAI21X1 U1094 ( .A(n1847), .B(n1729), .C(n2406), .Y(n1893) );
  NAND2X1 U1095 ( .A(\mem<1><2> ), .B(n1731), .Y(n2406) );
  OAI21X1 U1096 ( .A(n1846), .B(n1729), .C(n2405), .Y(n1892) );
  NAND2X1 U1097 ( .A(\mem<1><3> ), .B(n1731), .Y(n2405) );
  OAI21X1 U1098 ( .A(n1845), .B(n1729), .C(n2404), .Y(n1891) );
  NAND2X1 U1099 ( .A(\mem<1><4> ), .B(n1731), .Y(n2404) );
  OAI21X1 U1100 ( .A(n1843), .B(n1729), .C(n2403), .Y(n1890) );
  NAND2X1 U1101 ( .A(\mem<1><5> ), .B(n1731), .Y(n2403) );
  OAI21X1 U1102 ( .A(n1841), .B(n1729), .C(n2402), .Y(n1889) );
  NAND2X1 U1103 ( .A(\mem<1><6> ), .B(n1731), .Y(n2402) );
  OAI21X1 U1104 ( .A(n1840), .B(n1729), .C(n2401), .Y(n1888) );
  NAND2X1 U1105 ( .A(\mem<1><7> ), .B(n1731), .Y(n2401) );
  OAI21X1 U1106 ( .A(n1839), .B(n1729), .C(n2400), .Y(n1887) );
  NAND2X1 U1107 ( .A(\mem<1><8> ), .B(n1730), .Y(n2400) );
  OAI21X1 U1108 ( .A(n1837), .B(n1729), .C(n2399), .Y(n1886) );
  NAND2X1 U1109 ( .A(\mem<1><9> ), .B(n1730), .Y(n2399) );
  OAI21X1 U1110 ( .A(n1835), .B(n1729), .C(n2398), .Y(n1885) );
  NAND2X1 U1111 ( .A(\mem<1><10> ), .B(n1730), .Y(n2398) );
  OAI21X1 U1112 ( .A(n1834), .B(n1729), .C(n2397), .Y(n1884) );
  NAND2X1 U1113 ( .A(\mem<1><11> ), .B(n1730), .Y(n2397) );
  OAI21X1 U1114 ( .A(n1832), .B(n1729), .C(n2396), .Y(n1883) );
  NAND2X1 U1115 ( .A(\mem<1><12> ), .B(n1730), .Y(n2396) );
  OAI21X1 U1116 ( .A(n1830), .B(n1729), .C(n2395), .Y(n1882) );
  NAND2X1 U1117 ( .A(\mem<1><13> ), .B(n1730), .Y(n2395) );
  OAI21X1 U1118 ( .A(n1828), .B(n1729), .C(n2394), .Y(n1881) );
  NAND2X1 U1119 ( .A(\mem<1><14> ), .B(n1730), .Y(n2394) );
  OAI21X1 U1120 ( .A(n1826), .B(n1729), .C(n2393), .Y(n1880) );
  NAND2X1 U1121 ( .A(\mem<1><15> ), .B(n1730), .Y(n2393) );
  NOR3X1 U1124 ( .A(n1852), .B(n1691), .C(n1709), .Y(n2782) );
  OAI21X1 U1125 ( .A(n1851), .B(n1726), .C(n2392), .Y(n1879) );
  NAND2X1 U1126 ( .A(\mem<0><0> ), .B(n1728), .Y(n2392) );
  OAI21X1 U1128 ( .A(n1850), .B(n1726), .C(n2391), .Y(n1878) );
  NAND2X1 U1129 ( .A(\mem<0><1> ), .B(n1728), .Y(n2391) );
  OAI21X1 U1131 ( .A(n1848), .B(n1726), .C(n2390), .Y(n1877) );
  NAND2X1 U1132 ( .A(\mem<0><2> ), .B(n1728), .Y(n2390) );
  OAI21X1 U1134 ( .A(n1846), .B(n1726), .C(n2389), .Y(n1876) );
  NAND2X1 U1135 ( .A(\mem<0><3> ), .B(n1728), .Y(n2389) );
  OAI21X1 U1137 ( .A(n1845), .B(n1726), .C(n2388), .Y(n1875) );
  NAND2X1 U1138 ( .A(\mem<0><4> ), .B(n1728), .Y(n2388) );
  OAI21X1 U1140 ( .A(n1844), .B(n1726), .C(n2387), .Y(n1874) );
  NAND2X1 U1141 ( .A(\mem<0><5> ), .B(n1728), .Y(n2387) );
  OAI21X1 U1143 ( .A(n1842), .B(n1726), .C(n2386), .Y(n1873) );
  NAND2X1 U1144 ( .A(\mem<0><6> ), .B(n1728), .Y(n2386) );
  OAI21X1 U1146 ( .A(n1840), .B(n1726), .C(n2385), .Y(n1872) );
  NAND2X1 U1147 ( .A(\mem<0><7> ), .B(n1728), .Y(n2385) );
  OAI21X1 U1149 ( .A(n1839), .B(n1726), .C(n2384), .Y(n1871) );
  NAND2X1 U1150 ( .A(\mem<0><8> ), .B(n1727), .Y(n2384) );
  OAI21X1 U1152 ( .A(n1838), .B(n1726), .C(n2383), .Y(n1870) );
  NAND2X1 U1153 ( .A(\mem<0><9> ), .B(n1727), .Y(n2383) );
  OAI21X1 U1155 ( .A(n1836), .B(n1726), .C(n2382), .Y(n1869) );
  NAND2X1 U1156 ( .A(\mem<0><10> ), .B(n1727), .Y(n2382) );
  OAI21X1 U1158 ( .A(n1834), .B(n1726), .C(n2381), .Y(n1868) );
  NAND2X1 U1159 ( .A(\mem<0><11> ), .B(n1727), .Y(n2381) );
  OAI21X1 U1161 ( .A(n1833), .B(n1726), .C(n2380), .Y(n1867) );
  NAND2X1 U1162 ( .A(\mem<0><12> ), .B(n1727), .Y(n2380) );
  OAI21X1 U1164 ( .A(n1831), .B(n1726), .C(n2379), .Y(n1866) );
  NAND2X1 U1165 ( .A(\mem<0><13> ), .B(n1727), .Y(n2379) );
  OAI21X1 U1167 ( .A(n1829), .B(n1726), .C(n2378), .Y(n1865) );
  NAND2X1 U1168 ( .A(\mem<0><14> ), .B(n1727), .Y(n2378) );
  OAI21X1 U1170 ( .A(n1827), .B(n1726), .C(n2377), .Y(n1864) );
  NAND2X1 U1171 ( .A(\mem<0><15> ), .B(n1727), .Y(n2377) );
  NOR3X1 U1174 ( .A(n1852), .B(n1691), .C(n1724), .Y(n2765) );
  NAND3X1 U1175 ( .A(n1856), .B(n1858), .C(n2763), .Y(n2376) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2763) );
  INVX4 U3 ( .A(n5), .Y(n4) );
  AND2X2 U4 ( .A(\data_in<9> ), .B(n1822), .Y(n43) );
  AND2X2 U5 ( .A(\data_in<10> ), .B(n1822), .Y(n42) );
  AND2X2 U6 ( .A(\data_in<0> ), .B(n1824), .Y(n58) );
  AND2X2 U7 ( .A(\data_in<1> ), .B(n1824), .Y(n56) );
  AND2X2 U8 ( .A(\data_in<2> ), .B(n1824), .Y(n54) );
  AND2X2 U9 ( .A(\data_in<3> ), .B(n1824), .Y(n52) );
  AND2X2 U10 ( .A(\data_in<4> ), .B(n1824), .Y(n50) );
  AND2X2 U11 ( .A(\data_in<5> ), .B(n1824), .Y(n48) );
  AND2X2 U12 ( .A(\data_in<6> ), .B(n1824), .Y(n47) );
  AND2X2 U13 ( .A(\data_in<7> ), .B(n1824), .Y(n45) );
  AND2X2 U14 ( .A(\data_in<11> ), .B(n1824), .Y(n41) );
  AND2X2 U15 ( .A(\data_in<12> ), .B(n1824), .Y(n40) );
  AND2X2 U16 ( .A(\data_in<15> ), .B(n1824), .Y(n37) );
  AND2X2 U17 ( .A(\data_in<8> ), .B(n1823), .Y(n44) );
  AND2X2 U18 ( .A(\data_in<13> ), .B(n1823), .Y(n39) );
  AND2X2 U19 ( .A(\data_in<14> ), .B(n1823), .Y(n38) );
  INVX1 U20 ( .A(N10), .Y(n1710) );
  INVX2 U21 ( .A(n1711), .Y(n1712) );
  INVX2 U22 ( .A(n1709), .Y(n1718) );
  INVX2 U23 ( .A(n1709), .Y(n1717) );
  INVX2 U24 ( .A(n1709), .Y(n1716) );
  INVX2 U25 ( .A(n1710), .Y(n1715) );
  INVX2 U26 ( .A(n1710), .Y(n1714) );
  INVX1 U27 ( .A(n1709), .Y(n1721) );
  INVX1 U28 ( .A(n1710), .Y(n1713) );
  INVX1 U29 ( .A(n1725), .Y(n1720) );
  INVX1 U30 ( .A(n1725), .Y(n1723) );
  INVX1 U31 ( .A(n1725), .Y(n1722) );
  INVX1 U32 ( .A(n1725), .Y(n1724) );
  INVX1 U33 ( .A(N10), .Y(n1709) );
  INVX1 U34 ( .A(n1719), .Y(n1711) );
  INVX1 U35 ( .A(n1698), .Y(n1703) );
  INVX1 U36 ( .A(n1697), .Y(n1705) );
  INVX1 U37 ( .A(n1697), .Y(n1706) );
  INVX1 U38 ( .A(n1698), .Y(n1707) );
  INVX2 U39 ( .A(n1697), .Y(n1708) );
  INVX1 U40 ( .A(n1853), .Y(n1700) );
  INVX2 U41 ( .A(n1698), .Y(n1701) );
  INVX2 U42 ( .A(n1698), .Y(n1702) );
  INVX2 U43 ( .A(n1697), .Y(n1704) );
  INVX1 U44 ( .A(n1856), .Y(n1688) );
  INVX1 U45 ( .A(n1856), .Y(n1690) );
  INVX1 U46 ( .A(n1856), .Y(n1689) );
  INVX2 U47 ( .A(n1854), .Y(n1691) );
  INVX1 U48 ( .A(n1853), .Y(n1699) );
  INVX1 U49 ( .A(n1858), .Y(n1687) );
  INVX1 U50 ( .A(N14), .Y(n1858) );
  INVX1 U51 ( .A(N13), .Y(n1856) );
  INVX1 U52 ( .A(N10), .Y(n1725) );
  INVX1 U53 ( .A(n1853), .Y(n1852) );
  INVX1 U54 ( .A(rst), .Y(n1859) );
  INVX1 U55 ( .A(n68), .Y(n1726) );
  INVX1 U56 ( .A(N12), .Y(n1854) );
  INVX1 U57 ( .A(n70), .Y(n1729) );
  INVX1 U58 ( .A(n101), .Y(n1750) );
  INVX1 U59 ( .A(n118), .Y(n1753) );
  INVX1 U60 ( .A(n177), .Y(n1774) );
  INVX1 U93 ( .A(n194), .Y(n1777) );
  INVX4 U94 ( .A(n2885), .Y(n1825) );
  INVX1 U127 ( .A(n1852), .Y(n1697) );
  INVX1 U128 ( .A(n1852), .Y(n1698) );
  INVX1 U161 ( .A(n72), .Y(n1732) );
  INVX1 U162 ( .A(n74), .Y(n1735) );
  INVX1 U195 ( .A(n76), .Y(n1738) );
  INVX1 U196 ( .A(n80), .Y(n1741) );
  INVX1 U229 ( .A(n82), .Y(n1744) );
  INVX1 U230 ( .A(n99), .Y(n1747) );
  INVX1 U263 ( .A(n120), .Y(n1756) );
  INVX1 U264 ( .A(n137), .Y(n1759) );
  INVX1 U297 ( .A(n139), .Y(n1762) );
  INVX1 U298 ( .A(n156), .Y(n1765) );
  INVX1 U331 ( .A(n158), .Y(n1768) );
  INVX1 U332 ( .A(n175), .Y(n1771) );
  INVX1 U366 ( .A(n196), .Y(n1780) );
  INVX1 U367 ( .A(n215), .Y(n1783) );
  INVX1 U400 ( .A(n217), .Y(n1786) );
  INVX1 U401 ( .A(n233), .Y(n1789) );
  INVX1 U434 ( .A(n235), .Y(n1792) );
  INVX1 U435 ( .A(n251), .Y(n1795) );
  INVX1 U468 ( .A(n253), .Y(n1798) );
  INVX1 U469 ( .A(n269), .Y(n1801) );
  INVX1 U502 ( .A(n271), .Y(n1804) );
  INVX1 U503 ( .A(n287), .Y(n1807) );
  INVX1 U536 ( .A(n289), .Y(n1810) );
  INVX1 U537 ( .A(n305), .Y(n1813) );
  INVX1 U570 ( .A(n307), .Y(n1816) );
  INVX1 U571 ( .A(n323), .Y(n1819) );
  AND2X2 U604 ( .A(n3), .B(N31), .Y(\data_out<1> ) );
  INVX1 U605 ( .A(n1672), .Y(N31) );
  INVX1 U639 ( .A(n5), .Y(n2) );
  INVX1 U640 ( .A(n4), .Y(n3) );
  AND2X2 U673 ( .A(n6), .B(n1859), .Y(n5) );
  INVX1 U674 ( .A(write), .Y(n6) );
  OR2X2 U707 ( .A(n4), .B(n1671), .Y(n7) );
  INVX1 U708 ( .A(n7), .Y(\data_out<0> ) );
  OR2X2 U741 ( .A(n4), .B(n1673), .Y(n9) );
  INVX1 U742 ( .A(n9), .Y(\data_out<2> ) );
  OR2X2 U775 ( .A(n2), .B(n1674), .Y(n11) );
  INVX1 U776 ( .A(n11), .Y(\data_out<3> ) );
  OR2X2 U809 ( .A(n4), .B(n1675), .Y(n13) );
  INVX1 U810 ( .A(n13), .Y(\data_out<4> ) );
  OR2X2 U843 ( .A(n4), .B(n1676), .Y(n15) );
  INVX1 U844 ( .A(n15), .Y(\data_out<5> ) );
  OR2X2 U877 ( .A(n4), .B(n1677), .Y(n17) );
  INVX1 U878 ( .A(n17), .Y(\data_out<6> ) );
  OR2X2 U912 ( .A(n2), .B(n1678), .Y(n19) );
  INVX1 U913 ( .A(n19), .Y(\data_out<7> ) );
  OR2X2 U947 ( .A(n4), .B(n1679), .Y(n21) );
  INVX1 U948 ( .A(n21), .Y(\data_out<8> ) );
  OR2X2 U982 ( .A(n4), .B(n1680), .Y(n23) );
  INVX1 U983 ( .A(n23), .Y(\data_out<9> ) );
  OR2X2 U1017 ( .A(n4), .B(n1681), .Y(n25) );
  INVX1 U1018 ( .A(n25), .Y(\data_out<10> ) );
  OR2X2 U1052 ( .A(n2), .B(n1682), .Y(n27) );
  INVX1 U1053 ( .A(n27), .Y(\data_out<11> ) );
  OR2X2 U1087 ( .A(n2), .B(n1683), .Y(n29) );
  INVX1 U1088 ( .A(n29), .Y(\data_out<12> ) );
  OR2X2 U1122 ( .A(n4), .B(n1684), .Y(n31) );
  INVX1 U1123 ( .A(n31), .Y(\data_out<13> ) );
  OR2X2 U1127 ( .A(n4), .B(n1686), .Y(n33) );
  INVX1 U1130 ( .A(n33), .Y(\data_out<15> ) );
  OR2X2 U1133 ( .A(n4), .B(n1685), .Y(n35) );
  INVX1 U1136 ( .A(n35), .Y(\data_out<14> ) );
  BUFX2 U1139 ( .A(n341), .Y(n1727) );
  BUFX2 U1142 ( .A(n341), .Y(n1728) );
  BUFX2 U1145 ( .A(n360), .Y(n1730) );
  BUFX2 U1148 ( .A(n360), .Y(n1731) );
  BUFX2 U1151 ( .A(n378), .Y(n1733) );
  BUFX2 U1154 ( .A(n378), .Y(n1734) );
  BUFX2 U1157 ( .A(n396), .Y(n1736) );
  BUFX2 U1160 ( .A(n396), .Y(n1737) );
  BUFX2 U1163 ( .A(n414), .Y(n1739) );
  BUFX2 U1166 ( .A(n414), .Y(n1740) );
  BUFX2 U1169 ( .A(n432), .Y(n1742) );
  BUFX2 U1172 ( .A(n432), .Y(n1743) );
  BUFX2 U1173 ( .A(n450), .Y(n1745) );
  BUFX2 U1177 ( .A(n450), .Y(n1746) );
  BUFX2 U1178 ( .A(n468), .Y(n1748) );
  BUFX2 U1179 ( .A(n468), .Y(n1749) );
  BUFX2 U1180 ( .A(n486), .Y(n1751) );
  BUFX2 U1181 ( .A(n486), .Y(n1752) );
  BUFX2 U1182 ( .A(n505), .Y(n1754) );
  BUFX2 U1183 ( .A(n505), .Y(n1755) );
  BUFX2 U1184 ( .A(n523), .Y(n1757) );
  BUFX2 U1185 ( .A(n523), .Y(n1758) );
  BUFX2 U1186 ( .A(n541), .Y(n1760) );
  BUFX2 U1187 ( .A(n541), .Y(n1761) );
  BUFX2 U1188 ( .A(n559), .Y(n1763) );
  BUFX2 U1189 ( .A(n559), .Y(n1764) );
  BUFX2 U1190 ( .A(n577), .Y(n1766) );
  BUFX2 U1191 ( .A(n577), .Y(n1767) );
  BUFX2 U1192 ( .A(n595), .Y(n1769) );
  BUFX2 U1193 ( .A(n595), .Y(n1770) );
  BUFX2 U1194 ( .A(n613), .Y(n1772) );
  BUFX2 U1195 ( .A(n613), .Y(n1773) );
  BUFX2 U1196 ( .A(n631), .Y(n1775) );
  BUFX2 U1197 ( .A(n631), .Y(n1776) );
  BUFX2 U1198 ( .A(n650), .Y(n1778) );
  BUFX2 U1199 ( .A(n650), .Y(n1779) );
  BUFX2 U1200 ( .A(n1164), .Y(n1781) );
  BUFX2 U1201 ( .A(n1164), .Y(n1782) );
  BUFX2 U1202 ( .A(n1166), .Y(n1784) );
  BUFX2 U1203 ( .A(n1166), .Y(n1785) );
  BUFX2 U1204 ( .A(n1168), .Y(n1787) );
  BUFX2 U1205 ( .A(n1168), .Y(n1788) );
  BUFX2 U1206 ( .A(n1170), .Y(n1790) );
  BUFX2 U1207 ( .A(n1170), .Y(n1791) );
  BUFX2 U1208 ( .A(n1172), .Y(n1793) );
  BUFX2 U1209 ( .A(n1172), .Y(n1794) );
  BUFX2 U1210 ( .A(n1174), .Y(n1796) );
  BUFX2 U1211 ( .A(n1174), .Y(n1797) );
  BUFX2 U1212 ( .A(n1176), .Y(n1799) );
  BUFX2 U1213 ( .A(n1176), .Y(n1800) );
  BUFX2 U1214 ( .A(n1178), .Y(n1802) );
  BUFX2 U1215 ( .A(n1178), .Y(n1803) );
  BUFX2 U1216 ( .A(n1180), .Y(n1805) );
  BUFX2 U1217 ( .A(n1180), .Y(n1806) );
  BUFX2 U1218 ( .A(n1182), .Y(n1808) );
  BUFX2 U1219 ( .A(n1182), .Y(n1809) );
  BUFX2 U1220 ( .A(n1184), .Y(n1811) );
  BUFX2 U1221 ( .A(n1184), .Y(n1812) );
  BUFX2 U1222 ( .A(n1186), .Y(n1814) );
  BUFX2 U1223 ( .A(n1186), .Y(n1815) );
  BUFX2 U1224 ( .A(n1188), .Y(n1817) );
  BUFX2 U1225 ( .A(n1188), .Y(n1818) );
  BUFX2 U1226 ( .A(n1190), .Y(n1820) );
  BUFX2 U1227 ( .A(n1190), .Y(n1821) );
  INVX1 U1228 ( .A(n1858), .Y(n1857) );
  INVX1 U1229 ( .A(n1856), .Y(n1855) );
  BUFX2 U1230 ( .A(n2376), .Y(n60) );
  INVX1 U1231 ( .A(n60), .Y(n1860) );
  BUFX2 U1232 ( .A(n2505), .Y(n62) );
  INVX1 U1233 ( .A(n62), .Y(n1863) );
  BUFX2 U1234 ( .A(n2634), .Y(n64) );
  INVX1 U1235 ( .A(n64), .Y(n1861) );
  BUFX2 U1236 ( .A(n2764), .Y(n66) );
  INVX1 U1237 ( .A(n66), .Y(n1862) );
  AND2X1 U1238 ( .A(n1860), .B(n2765), .Y(n68) );
  AND2X1 U1239 ( .A(n1860), .B(n2782), .Y(n70) );
  AND2X1 U1240 ( .A(n1860), .B(n2799), .Y(n72) );
  AND2X1 U1241 ( .A(n1860), .B(n2816), .Y(n74) );
  AND2X1 U1242 ( .A(n1860), .B(n2833), .Y(n76) );
  AND2X1 U1243 ( .A(n1860), .B(n2850), .Y(n80) );
  AND2X1 U1244 ( .A(n1860), .B(n2867), .Y(n82) );
  AND2X1 U1245 ( .A(n1860), .B(n2884), .Y(n99) );
  AND2X1 U1246 ( .A(n1863), .B(n2765), .Y(n101) );
  AND2X1 U1247 ( .A(n1863), .B(n2782), .Y(n118) );
  AND2X1 U1248 ( .A(n1863), .B(n2799), .Y(n120) );
  AND2X1 U1249 ( .A(n1863), .B(n2816), .Y(n137) );
  AND2X1 U1250 ( .A(n1863), .B(n2833), .Y(n139) );
  AND2X1 U1251 ( .A(n1863), .B(n2850), .Y(n156) );
  AND2X1 U1252 ( .A(n1863), .B(n2867), .Y(n158) );
  AND2X1 U1253 ( .A(n1863), .B(n2884), .Y(n175) );
  AND2X1 U1254 ( .A(n1861), .B(n2765), .Y(n177) );
  AND2X1 U1255 ( .A(n1861), .B(n2782), .Y(n194) );
  AND2X1 U1256 ( .A(n1861), .B(n2799), .Y(n196) );
  AND2X1 U1257 ( .A(n1861), .B(n2816), .Y(n215) );
  AND2X1 U1258 ( .A(n1861), .B(n2833), .Y(n217) );
  AND2X1 U1259 ( .A(n1861), .B(n2850), .Y(n233) );
  AND2X1 U1260 ( .A(n1861), .B(n2867), .Y(n235) );
  AND2X1 U1261 ( .A(n1861), .B(n2884), .Y(n251) );
  AND2X1 U1262 ( .A(n2765), .B(n1862), .Y(n253) );
  AND2X1 U1263 ( .A(n2782), .B(n1862), .Y(n269) );
  AND2X1 U1264 ( .A(n2799), .B(n1862), .Y(n271) );
  AND2X1 U1265 ( .A(n2816), .B(n1862), .Y(n287) );
  AND2X1 U1266 ( .A(n2833), .B(n1862), .Y(n289) );
  AND2X1 U1267 ( .A(n2850), .B(n1862), .Y(n305) );
  AND2X1 U1268 ( .A(n2867), .B(n1862), .Y(n307) );
  AND2X1 U1269 ( .A(n2884), .B(n1862), .Y(n323) );
  AND2X1 U1270 ( .A(n68), .B(n1823), .Y(n325) );
  INVX1 U1271 ( .A(n325), .Y(n341) );
  AND2X1 U1272 ( .A(n70), .B(n1824), .Y(n343) );
  INVX1 U1273 ( .A(n343), .Y(n360) );
  AND2X1 U1274 ( .A(n72), .B(n1824), .Y(n362) );
  INVX1 U1275 ( .A(n362), .Y(n378) );
  AND2X1 U1276 ( .A(n74), .B(n1824), .Y(n380) );
  INVX1 U1277 ( .A(n380), .Y(n396) );
  AND2X1 U1278 ( .A(n76), .B(n1824), .Y(n398) );
  INVX1 U1279 ( .A(n398), .Y(n414) );
  AND2X1 U1280 ( .A(n80), .B(n1824), .Y(n416) );
  INVX1 U1281 ( .A(n416), .Y(n432) );
  AND2X1 U1282 ( .A(n82), .B(n1823), .Y(n434) );
  INVX1 U1283 ( .A(n434), .Y(n450) );
  AND2X1 U1284 ( .A(n99), .B(n1823), .Y(n452) );
  INVX1 U1285 ( .A(n452), .Y(n468) );
  AND2X1 U1286 ( .A(n101), .B(n1823), .Y(n470) );
  INVX1 U1287 ( .A(n470), .Y(n486) );
  AND2X1 U1288 ( .A(n118), .B(n1823), .Y(n488) );
  INVX1 U1289 ( .A(n488), .Y(n505) );
  AND2X1 U1290 ( .A(n120), .B(n1823), .Y(n507) );
  INVX1 U1291 ( .A(n507), .Y(n523) );
  AND2X1 U1292 ( .A(n137), .B(n1823), .Y(n525) );
  INVX1 U1293 ( .A(n525), .Y(n541) );
  AND2X1 U1294 ( .A(n139), .B(n1823), .Y(n543) );
  INVX1 U1295 ( .A(n543), .Y(n559) );
  AND2X1 U1296 ( .A(n156), .B(n1823), .Y(n561) );
  INVX1 U1297 ( .A(n561), .Y(n577) );
  AND2X1 U1298 ( .A(n158), .B(n1823), .Y(n579) );
  INVX1 U1299 ( .A(n579), .Y(n595) );
  AND2X1 U1300 ( .A(n175), .B(n1823), .Y(n597) );
  INVX1 U1301 ( .A(n597), .Y(n613) );
  AND2X1 U1302 ( .A(n177), .B(n1823), .Y(n615) );
  INVX1 U1303 ( .A(n615), .Y(n631) );
  AND2X1 U1304 ( .A(n194), .B(n1823), .Y(n633) );
  INVX1 U1305 ( .A(n633), .Y(n650) );
  AND2X1 U1306 ( .A(n196), .B(n1823), .Y(n1163) );
  INVX1 U1307 ( .A(n1163), .Y(n1164) );
  AND2X1 U1308 ( .A(n215), .B(n1822), .Y(n1165) );
  INVX1 U1309 ( .A(n1165), .Y(n1166) );
  AND2X1 U1310 ( .A(n217), .B(n1822), .Y(n1167) );
  INVX1 U1311 ( .A(n1167), .Y(n1168) );
  AND2X1 U1312 ( .A(n233), .B(n1822), .Y(n1169) );
  INVX1 U1313 ( .A(n1169), .Y(n1170) );
  AND2X1 U1314 ( .A(n235), .B(n1822), .Y(n1171) );
  INVX1 U1315 ( .A(n1171), .Y(n1172) );
  AND2X1 U1316 ( .A(n251), .B(n1822), .Y(n1173) );
  INVX1 U1317 ( .A(n1173), .Y(n1174) );
  AND2X1 U1318 ( .A(n253), .B(n1822), .Y(n1175) );
  INVX1 U1319 ( .A(n1175), .Y(n1176) );
  AND2X1 U1320 ( .A(n269), .B(n1822), .Y(n1177) );
  INVX1 U1321 ( .A(n1177), .Y(n1178) );
  AND2X1 U1322 ( .A(n271), .B(n1822), .Y(n1179) );
  INVX1 U1323 ( .A(n1179), .Y(n1180) );
  AND2X1 U1324 ( .A(n287), .B(n1822), .Y(n1181) );
  INVX1 U1325 ( .A(n1181), .Y(n1182) );
  AND2X1 U1326 ( .A(n289), .B(n1822), .Y(n1183) );
  INVX1 U1327 ( .A(n1183), .Y(n1184) );
  AND2X1 U1328 ( .A(n305), .B(n1822), .Y(n1185) );
  INVX1 U1329 ( .A(n1185), .Y(n1186) );
  AND2X1 U1330 ( .A(n307), .B(n1822), .Y(n1187) );
  INVX1 U1331 ( .A(n1187), .Y(n1188) );
  AND2X1 U1332 ( .A(n323), .B(n1822), .Y(n1189) );
  INVX1 U1333 ( .A(n1189), .Y(n1190) );
  MUX2X1 U1334 ( .B(n1192), .A(n1193), .S(n1699), .Y(n1191) );
  MUX2X1 U1335 ( .B(n1195), .A(n1196), .S(n1699), .Y(n1194) );
  MUX2X1 U1336 ( .B(n1198), .A(n1199), .S(n1699), .Y(n1197) );
  MUX2X1 U1337 ( .B(n1201), .A(n1202), .S(n1699), .Y(n1200) );
  MUX2X1 U1338 ( .B(n1204), .A(n1205), .S(n1690), .Y(n1203) );
  MUX2X1 U1339 ( .B(n1207), .A(n1208), .S(n1699), .Y(n1206) );
  MUX2X1 U1340 ( .B(n1210), .A(n1211), .S(n1699), .Y(n1209) );
  MUX2X1 U1341 ( .B(n1213), .A(n1214), .S(n1699), .Y(n1212) );
  MUX2X1 U1342 ( .B(n1216), .A(n1217), .S(n1699), .Y(n1215) );
  MUX2X1 U1343 ( .B(n1219), .A(n1220), .S(n1690), .Y(n1218) );
  MUX2X1 U1344 ( .B(n1222), .A(n1223), .S(n1700), .Y(n1221) );
  MUX2X1 U1345 ( .B(n1225), .A(n1226), .S(n1700), .Y(n1224) );
  MUX2X1 U1346 ( .B(n1228), .A(n1229), .S(n1700), .Y(n1227) );
  MUX2X1 U1347 ( .B(n1231), .A(n1232), .S(n1700), .Y(n1230) );
  MUX2X1 U1348 ( .B(n1234), .A(n1235), .S(n1690), .Y(n1233) );
  MUX2X1 U1349 ( .B(n1237), .A(n1238), .S(n1700), .Y(n1236) );
  MUX2X1 U1350 ( .B(n1240), .A(n1241), .S(n1700), .Y(n1239) );
  MUX2X1 U1351 ( .B(n1243), .A(n1244), .S(n1700), .Y(n1242) );
  MUX2X1 U1352 ( .B(n1246), .A(n1247), .S(n1700), .Y(n1245) );
  MUX2X1 U1353 ( .B(n1249), .A(n1250), .S(n1690), .Y(n1248) );
  MUX2X1 U1354 ( .B(n1252), .A(n1253), .S(n1700), .Y(n1251) );
  MUX2X1 U1355 ( .B(n1255), .A(n1256), .S(n1700), .Y(n1254) );
  MUX2X1 U1356 ( .B(n1258), .A(n1259), .S(n1700), .Y(n1257) );
  MUX2X1 U1357 ( .B(n1261), .A(n1262), .S(n1700), .Y(n1260) );
  MUX2X1 U1358 ( .B(n1264), .A(n1265), .S(n1690), .Y(n1263) );
  MUX2X1 U1359 ( .B(n1267), .A(n1268), .S(n1700), .Y(n1266) );
  MUX2X1 U1360 ( .B(n1270), .A(n1271), .S(n1699), .Y(n1269) );
  MUX2X1 U1361 ( .B(n1273), .A(n1274), .S(n1700), .Y(n1272) );
  MUX2X1 U1362 ( .B(n1276), .A(n1277), .S(n1699), .Y(n1275) );
  MUX2X1 U1363 ( .B(n1279), .A(n1280), .S(n1690), .Y(n1278) );
  MUX2X1 U1364 ( .B(n1282), .A(n1283), .S(n1700), .Y(n1281) );
  MUX2X1 U1365 ( .B(n1285), .A(n1286), .S(n1700), .Y(n1284) );
  MUX2X1 U1366 ( .B(n1288), .A(n1289), .S(n1699), .Y(n1287) );
  MUX2X1 U1367 ( .B(n1291), .A(n1292), .S(n1700), .Y(n1290) );
  MUX2X1 U1368 ( .B(n1294), .A(n1295), .S(n1690), .Y(n1293) );
  MUX2X1 U1369 ( .B(n1297), .A(n1298), .S(n1699), .Y(n1296) );
  MUX2X1 U1370 ( .B(n1300), .A(n1301), .S(n1700), .Y(n1299) );
  MUX2X1 U1371 ( .B(n1303), .A(n1304), .S(n1699), .Y(n1302) );
  MUX2X1 U1372 ( .B(n1306), .A(n1307), .S(n1700), .Y(n1305) );
  MUX2X1 U1373 ( .B(n1309), .A(n1310), .S(n1690), .Y(n1308) );
  MUX2X1 U1374 ( .B(n1312), .A(n1313), .S(n1701), .Y(n1311) );
  MUX2X1 U1375 ( .B(n1315), .A(n1316), .S(n1701), .Y(n1314) );
  MUX2X1 U1376 ( .B(n1318), .A(n1319), .S(n1701), .Y(n1317) );
  MUX2X1 U1377 ( .B(n1321), .A(n1322), .S(n1701), .Y(n1320) );
  MUX2X1 U1378 ( .B(n1324), .A(n1325), .S(n1690), .Y(n1323) );
  MUX2X1 U1379 ( .B(n1327), .A(n1328), .S(n1701), .Y(n1326) );
  MUX2X1 U1380 ( .B(n1330), .A(n1331), .S(n1701), .Y(n1329) );
  MUX2X1 U1381 ( .B(n1333), .A(n1334), .S(n1701), .Y(n1332) );
  MUX2X1 U1382 ( .B(n1336), .A(n1337), .S(n1701), .Y(n1335) );
  MUX2X1 U1383 ( .B(n1339), .A(n1340), .S(n1690), .Y(n1338) );
  MUX2X1 U1384 ( .B(n1342), .A(n1343), .S(n1701), .Y(n1341) );
  MUX2X1 U1385 ( .B(n1345), .A(n1346), .S(n1701), .Y(n1344) );
  MUX2X1 U1386 ( .B(n1348), .A(n1349), .S(n1701), .Y(n1347) );
  MUX2X1 U1387 ( .B(n1351), .A(n1352), .S(n1701), .Y(n1350) );
  MUX2X1 U1388 ( .B(n1354), .A(n1355), .S(n1690), .Y(n1353) );
  MUX2X1 U1389 ( .B(n1357), .A(n1358), .S(n1702), .Y(n1356) );
  MUX2X1 U1390 ( .B(n1360), .A(n1361), .S(n1702), .Y(n1359) );
  MUX2X1 U1391 ( .B(n1363), .A(n1364), .S(n1702), .Y(n1362) );
  MUX2X1 U1392 ( .B(n1366), .A(n1367), .S(n1702), .Y(n1365) );
  MUX2X1 U1393 ( .B(n1369), .A(n1370), .S(n1690), .Y(n1368) );
  MUX2X1 U1394 ( .B(n1372), .A(n1373), .S(n1702), .Y(n1371) );
  MUX2X1 U1395 ( .B(n1375), .A(n1376), .S(n1702), .Y(n1374) );
  MUX2X1 U1396 ( .B(n1378), .A(n1379), .S(n1702), .Y(n1377) );
  MUX2X1 U1397 ( .B(n1381), .A(n1382), .S(n1702), .Y(n1380) );
  MUX2X1 U1398 ( .B(n1384), .A(n1385), .S(n1689), .Y(n1383) );
  MUX2X1 U1399 ( .B(n1387), .A(n1388), .S(n1702), .Y(n1386) );
  MUX2X1 U1400 ( .B(n1390), .A(n1391), .S(n1702), .Y(n1389) );
  MUX2X1 U1401 ( .B(n1393), .A(n1394), .S(n1702), .Y(n1392) );
  MUX2X1 U1402 ( .B(n1396), .A(n1397), .S(n1702), .Y(n1395) );
  MUX2X1 U1403 ( .B(n1399), .A(n1400), .S(n1689), .Y(n1398) );
  MUX2X1 U1404 ( .B(n1402), .A(n1403), .S(n1703), .Y(n1401) );
  MUX2X1 U1405 ( .B(n1405), .A(n1406), .S(n1703), .Y(n1404) );
  MUX2X1 U1406 ( .B(n1408), .A(n1409), .S(n1703), .Y(n1407) );
  MUX2X1 U1407 ( .B(n1411), .A(n1412), .S(n1703), .Y(n1410) );
  MUX2X1 U1408 ( .B(n1414), .A(n1415), .S(n1689), .Y(n1413) );
  MUX2X1 U1409 ( .B(n1417), .A(n1418), .S(n1703), .Y(n1416) );
  MUX2X1 U1410 ( .B(n1420), .A(n1421), .S(n1703), .Y(n1419) );
  MUX2X1 U1411 ( .B(n1423), .A(n1424), .S(n1703), .Y(n1422) );
  MUX2X1 U1412 ( .B(n1426), .A(n1427), .S(n1703), .Y(n1425) );
  MUX2X1 U1413 ( .B(n1429), .A(n1430), .S(n1689), .Y(n1428) );
  MUX2X1 U1414 ( .B(n1432), .A(n1433), .S(n1703), .Y(n1431) );
  MUX2X1 U1415 ( .B(n1435), .A(n1436), .S(n1703), .Y(n1434) );
  MUX2X1 U1416 ( .B(n1438), .A(n1439), .S(n1703), .Y(n1437) );
  MUX2X1 U1417 ( .B(n1441), .A(n1442), .S(n1703), .Y(n1440) );
  MUX2X1 U1418 ( .B(n1444), .A(n1445), .S(n1689), .Y(n1443) );
  MUX2X1 U1419 ( .B(n1447), .A(n1448), .S(n1704), .Y(n1446) );
  MUX2X1 U1420 ( .B(n1450), .A(n1451), .S(n1704), .Y(n1449) );
  MUX2X1 U1421 ( .B(n1453), .A(n1454), .S(n1704), .Y(n1452) );
  MUX2X1 U1422 ( .B(n1456), .A(n1457), .S(n1704), .Y(n1455) );
  MUX2X1 U1423 ( .B(n1459), .A(n1460), .S(n1689), .Y(n1458) );
  MUX2X1 U1424 ( .B(n1462), .A(n1463), .S(n1704), .Y(n1461) );
  MUX2X1 U1425 ( .B(n1465), .A(n1466), .S(n1704), .Y(n1464) );
  MUX2X1 U1426 ( .B(n1468), .A(n1469), .S(n1704), .Y(n1467) );
  MUX2X1 U1427 ( .B(n1471), .A(n1472), .S(n1704), .Y(n1470) );
  MUX2X1 U1428 ( .B(n1474), .A(n1475), .S(n1689), .Y(n1473) );
  MUX2X1 U1429 ( .B(n1477), .A(n1478), .S(n1704), .Y(n1476) );
  MUX2X1 U1430 ( .B(n1480), .A(n1481), .S(n1704), .Y(n1479) );
  MUX2X1 U1431 ( .B(n1483), .A(n1484), .S(n1704), .Y(n1482) );
  MUX2X1 U1432 ( .B(n1486), .A(n1487), .S(n1704), .Y(n1485) );
  MUX2X1 U1433 ( .B(n1489), .A(n1490), .S(n1689), .Y(n1488) );
  MUX2X1 U1434 ( .B(n1492), .A(n1493), .S(n1705), .Y(n1491) );
  MUX2X1 U1435 ( .B(n1495), .A(n1496), .S(n1705), .Y(n1494) );
  MUX2X1 U1436 ( .B(n1498), .A(n1499), .S(n1705), .Y(n1497) );
  MUX2X1 U1437 ( .B(n1501), .A(n1502), .S(n1705), .Y(n1500) );
  MUX2X1 U1438 ( .B(n1504), .A(n1505), .S(n1689), .Y(n1503) );
  MUX2X1 U1439 ( .B(n1507), .A(n1508), .S(n1705), .Y(n1506) );
  MUX2X1 U1440 ( .B(n1510), .A(n1511), .S(n1705), .Y(n1509) );
  MUX2X1 U1441 ( .B(n1513), .A(n1514), .S(n1705), .Y(n1512) );
  MUX2X1 U1442 ( .B(n1516), .A(n1517), .S(n1705), .Y(n1515) );
  MUX2X1 U1443 ( .B(n1519), .A(n1520), .S(n1689), .Y(n1518) );
  MUX2X1 U1444 ( .B(n1522), .A(n1523), .S(n1705), .Y(n1521) );
  MUX2X1 U1445 ( .B(n1525), .A(n1526), .S(n1705), .Y(n1524) );
  MUX2X1 U1446 ( .B(n1528), .A(n1529), .S(n1705), .Y(n1527) );
  MUX2X1 U1447 ( .B(n1531), .A(n1532), .S(n1705), .Y(n1530) );
  MUX2X1 U1448 ( .B(n1534), .A(n1535), .S(n1689), .Y(n1533) );
  MUX2X1 U1449 ( .B(n1537), .A(n1538), .S(n1706), .Y(n1536) );
  MUX2X1 U1450 ( .B(n1540), .A(n1541), .S(n1706), .Y(n1539) );
  MUX2X1 U1451 ( .B(n1543), .A(n1544), .S(n1706), .Y(n1542) );
  MUX2X1 U1452 ( .B(n1546), .A(n1547), .S(n1706), .Y(n1545) );
  MUX2X1 U1453 ( .B(n1549), .A(n1550), .S(n1689), .Y(n1548) );
  MUX2X1 U1454 ( .B(n1552), .A(n1553), .S(n1706), .Y(n1551) );
  MUX2X1 U1455 ( .B(n1555), .A(n1556), .S(n1706), .Y(n1554) );
  MUX2X1 U1456 ( .B(n1558), .A(n1559), .S(n1706), .Y(n1557) );
  MUX2X1 U1457 ( .B(n1561), .A(n1562), .S(n1706), .Y(n1560) );
  MUX2X1 U1458 ( .B(n1564), .A(n1565), .S(n1688), .Y(n1563) );
  MUX2X1 U1459 ( .B(n1567), .A(n1568), .S(n1706), .Y(n1566) );
  MUX2X1 U1460 ( .B(n1570), .A(n1571), .S(n1706), .Y(n1569) );
  MUX2X1 U1461 ( .B(n1573), .A(n1574), .S(n1706), .Y(n1572) );
  MUX2X1 U1462 ( .B(n1576), .A(n1577), .S(n1706), .Y(n1575) );
  MUX2X1 U1463 ( .B(n1579), .A(n1580), .S(n1688), .Y(n1578) );
  MUX2X1 U1464 ( .B(n1582), .A(n1583), .S(n1707), .Y(n1581) );
  MUX2X1 U1465 ( .B(n1585), .A(n1586), .S(n1707), .Y(n1584) );
  MUX2X1 U1466 ( .B(n1588), .A(n1589), .S(n1707), .Y(n1587) );
  MUX2X1 U1467 ( .B(n1591), .A(n1592), .S(n1707), .Y(n1590) );
  MUX2X1 U1468 ( .B(n1594), .A(n1595), .S(n1688), .Y(n1593) );
  MUX2X1 U1469 ( .B(n1597), .A(n1598), .S(n1707), .Y(n1596) );
  MUX2X1 U1470 ( .B(n1600), .A(n1601), .S(n1707), .Y(n1599) );
  MUX2X1 U1471 ( .B(n1603), .A(n1604), .S(n1707), .Y(n1602) );
  MUX2X1 U1472 ( .B(n1606), .A(n1607), .S(n1707), .Y(n1605) );
  MUX2X1 U1473 ( .B(n1609), .A(n1610), .S(n1688), .Y(n1608) );
  MUX2X1 U1474 ( .B(n1612), .A(n1613), .S(n1707), .Y(n1611) );
  MUX2X1 U1475 ( .B(n1615), .A(n1616), .S(n1707), .Y(n1614) );
  MUX2X1 U1476 ( .B(n1618), .A(n1619), .S(n1707), .Y(n1617) );
  MUX2X1 U1477 ( .B(n1621), .A(n1622), .S(n1707), .Y(n1620) );
  MUX2X1 U1478 ( .B(n1624), .A(n1625), .S(n1688), .Y(n1623) );
  MUX2X1 U1479 ( .B(n1627), .A(n1628), .S(n1708), .Y(n1626) );
  MUX2X1 U1480 ( .B(n1630), .A(n1631), .S(n1708), .Y(n1629) );
  MUX2X1 U1481 ( .B(n1633), .A(n1634), .S(n1708), .Y(n1632) );
  MUX2X1 U1482 ( .B(n1636), .A(n1637), .S(n1708), .Y(n1635) );
  MUX2X1 U1483 ( .B(n1639), .A(n1640), .S(n1688), .Y(n1638) );
  MUX2X1 U1484 ( .B(n1642), .A(n1643), .S(n1708), .Y(n1641) );
  MUX2X1 U1485 ( .B(n1645), .A(n1646), .S(n1708), .Y(n1644) );
  MUX2X1 U1486 ( .B(n1648), .A(n1649), .S(n1708), .Y(n1647) );
  MUX2X1 U1487 ( .B(n1651), .A(n1652), .S(n1708), .Y(n1650) );
  MUX2X1 U1488 ( .B(n1654), .A(n1655), .S(n1688), .Y(n1653) );
  MUX2X1 U1489 ( .B(n1657), .A(n1658), .S(n1708), .Y(n1656) );
  MUX2X1 U1490 ( .B(n1660), .A(n1661), .S(n1708), .Y(n1659) );
  MUX2X1 U1491 ( .B(n1663), .A(n1664), .S(n1708), .Y(n1662) );
  MUX2X1 U1492 ( .B(n1666), .A(n1667), .S(n1708), .Y(n1665) );
  MUX2X1 U1493 ( .B(n1669), .A(n1670), .S(n1688), .Y(n1668) );
  MUX2X1 U1494 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1722), .Y(n1193) );
  MUX2X1 U1495 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1712), .Y(n1192) );
  MUX2X1 U1496 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1716), .Y(n1196) );
  MUX2X1 U1497 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1718), .Y(n1195) );
  MUX2X1 U1498 ( .B(n1194), .A(n1191), .S(n1696), .Y(n1205) );
  MUX2X1 U1499 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1717), .Y(n1199) );
  MUX2X1 U1500 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1714), .Y(n1198) );
  MUX2X1 U1501 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1714), .Y(n1202) );
  MUX2X1 U1502 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1714), .Y(n1201) );
  MUX2X1 U1503 ( .B(n1200), .A(n1197), .S(n1696), .Y(n1204) );
  MUX2X1 U1504 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1714), .Y(n1208) );
  MUX2X1 U1505 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1714), .Y(n1207) );
  MUX2X1 U1506 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1714), .Y(n1211) );
  MUX2X1 U1507 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1714), .Y(n1210) );
  MUX2X1 U1508 ( .B(n1209), .A(n1206), .S(n1696), .Y(n1220) );
  MUX2X1 U1509 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1714), .Y(n1214) );
  MUX2X1 U1510 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1714), .Y(n1213) );
  MUX2X1 U1511 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1714), .Y(n1217) );
  MUX2X1 U1512 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1714), .Y(n1216) );
  MUX2X1 U1513 ( .B(n1215), .A(n1212), .S(n1696), .Y(n1219) );
  MUX2X1 U1514 ( .B(n1218), .A(n1203), .S(n1687), .Y(n1671) );
  MUX2X1 U1515 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1714), .Y(n1223) );
  MUX2X1 U1516 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1714), .Y(n1222) );
  MUX2X1 U1517 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1716), .Y(n1226) );
  MUX2X1 U1518 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1718), .Y(n1225) );
  MUX2X1 U1519 ( .B(n1224), .A(n1221), .S(n1696), .Y(n1235) );
  MUX2X1 U1520 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1716), .Y(n1229) );
  MUX2X1 U1521 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1714), .Y(n1228) );
  MUX2X1 U1522 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1714), .Y(n1232) );
  MUX2X1 U1523 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1722), .Y(n1231) );
  MUX2X1 U1524 ( .B(n1230), .A(n1227), .S(n1696), .Y(n1234) );
  MUX2X1 U1525 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1723), .Y(n1238) );
  MUX2X1 U1526 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1717), .Y(n1237) );
  MUX2X1 U1527 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1716), .Y(n1241) );
  MUX2X1 U1528 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1718), .Y(n1240) );
  MUX2X1 U1529 ( .B(n1239), .A(n1236), .S(n1696), .Y(n1250) );
  MUX2X1 U1530 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1719), .Y(n1244) );
  MUX2X1 U1531 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1719), .Y(n1243) );
  MUX2X1 U1532 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1724), .Y(n1247) );
  MUX2X1 U1533 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1719), .Y(n1246) );
  MUX2X1 U1534 ( .B(n1245), .A(n1242), .S(n1696), .Y(n1249) );
  MUX2X1 U1535 ( .B(n1248), .A(n1233), .S(n1687), .Y(n1672) );
  MUX2X1 U1536 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1719), .Y(n1253) );
  MUX2X1 U1537 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1723), .Y(n1252) );
  MUX2X1 U1538 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1719), .Y(n1256) );
  MUX2X1 U1539 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1719), .Y(n1255) );
  MUX2X1 U1540 ( .B(n1254), .A(n1251), .S(n1696), .Y(n1265) );
  MUX2X1 U1541 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1724), .Y(n1259) );
  MUX2X1 U1542 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1719), .Y(n1258) );
  MUX2X1 U1543 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1719), .Y(n1262) );
  MUX2X1 U1544 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1719), .Y(n1261) );
  MUX2X1 U1545 ( .B(n1260), .A(n1257), .S(n1696), .Y(n1264) );
  MUX2X1 U1546 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1716), .Y(n1268) );
  MUX2X1 U1547 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1716), .Y(n1267) );
  MUX2X1 U1548 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1716), .Y(n1271) );
  MUX2X1 U1549 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1719), .Y(n1270) );
  MUX2X1 U1550 ( .B(n1269), .A(n1266), .S(n1696), .Y(n1280) );
  MUX2X1 U1551 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1719), .Y(n1274) );
  MUX2X1 U1552 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1719), .Y(n1273) );
  MUX2X1 U1553 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1723), .Y(n1277) );
  MUX2X1 U1554 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1719), .Y(n1276) );
  MUX2X1 U1555 ( .B(n1275), .A(n1272), .S(n1696), .Y(n1279) );
  MUX2X1 U1556 ( .B(n1278), .A(n1263), .S(n1687), .Y(n1673) );
  MUX2X1 U1557 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1716), .Y(n1283) );
  MUX2X1 U1558 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1722), .Y(n1282) );
  MUX2X1 U1559 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1722), .Y(n1286) );
  MUX2X1 U1560 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1719), .Y(n1285) );
  MUX2X1 U1561 ( .B(n1284), .A(n1281), .S(n1695), .Y(n1295) );
  MUX2X1 U1562 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1717), .Y(n1289) );
  MUX2X1 U1563 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1717), .Y(n1288) );
  MUX2X1 U1564 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1718), .Y(n1292) );
  MUX2X1 U1565 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1717), .Y(n1291) );
  MUX2X1 U1566 ( .B(n1290), .A(n1287), .S(n1695), .Y(n1294) );
  MUX2X1 U1567 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1718), .Y(n1298) );
  MUX2X1 U1568 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1717), .Y(n1297) );
  MUX2X1 U1569 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1718), .Y(n1301) );
  MUX2X1 U1570 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1717), .Y(n1300) );
  MUX2X1 U1571 ( .B(n1299), .A(n1296), .S(n1695), .Y(n1310) );
  MUX2X1 U1572 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1718), .Y(n1304) );
  MUX2X1 U1573 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1718), .Y(n1303) );
  MUX2X1 U1574 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1717), .Y(n1307) );
  MUX2X1 U1575 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1717), .Y(n1306) );
  MUX2X1 U1576 ( .B(n1305), .A(n1302), .S(n1695), .Y(n1309) );
  MUX2X1 U1577 ( .B(n1308), .A(n1293), .S(n1687), .Y(n1674) );
  MUX2X1 U1578 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1719), .Y(n1313) );
  MUX2X1 U1579 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1719), .Y(n1312) );
  MUX2X1 U1580 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1719), .Y(n1316) );
  MUX2X1 U1581 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1719), .Y(n1315) );
  MUX2X1 U1582 ( .B(n1314), .A(n1311), .S(n1695), .Y(n1325) );
  MUX2X1 U1583 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1724), .Y(n1319) );
  MUX2X1 U1584 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1716), .Y(n1318) );
  MUX2X1 U1585 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1719), .Y(n1322) );
  MUX2X1 U1586 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1719), .Y(n1321) );
  MUX2X1 U1587 ( .B(n1320), .A(n1317), .S(n1695), .Y(n1324) );
  MUX2X1 U1588 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1719), .Y(n1328) );
  MUX2X1 U1589 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1719), .Y(n1327) );
  MUX2X1 U1590 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1719), .Y(n1331) );
  MUX2X1 U1591 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1719), .Y(n1330) );
  MUX2X1 U1592 ( .B(n1329), .A(n1326), .S(n1695), .Y(n1340) );
  MUX2X1 U1593 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1715), .Y(n1334) );
  MUX2X1 U1594 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1715), .Y(n1333) );
  MUX2X1 U1595 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1715), .Y(n1337) );
  MUX2X1 U1596 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1715), .Y(n1336) );
  MUX2X1 U1597 ( .B(n1335), .A(n1332), .S(n1695), .Y(n1339) );
  MUX2X1 U1598 ( .B(n1338), .A(n1323), .S(n1687), .Y(n1675) );
  MUX2X1 U1599 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1715), .Y(n1343) );
  MUX2X1 U1600 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1715), .Y(n1342) );
  MUX2X1 U1601 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1715), .Y(n1346) );
  MUX2X1 U1602 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1715), .Y(n1345) );
  MUX2X1 U1603 ( .B(n1344), .A(n1341), .S(n1695), .Y(n1355) );
  MUX2X1 U1604 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1715), .Y(n1349) );
  MUX2X1 U1605 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1715), .Y(n1348) );
  MUX2X1 U1606 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1715), .Y(n1352) );
  MUX2X1 U1607 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1715), .Y(n1351) );
  MUX2X1 U1608 ( .B(n1350), .A(n1347), .S(n1695), .Y(n1354) );
  MUX2X1 U1609 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1712), .Y(n1358) );
  MUX2X1 U1610 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1712), .Y(n1357) );
  MUX2X1 U1611 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1712), .Y(n1361) );
  MUX2X1 U1612 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1712), .Y(n1360) );
  MUX2X1 U1613 ( .B(n1359), .A(n1356), .S(n1695), .Y(n1370) );
  MUX2X1 U1614 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1712), .Y(n1364) );
  MUX2X1 U1615 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1712), .Y(n1363) );
  MUX2X1 U1616 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1712), .Y(n1367) );
  MUX2X1 U1617 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1712), .Y(n1366) );
  MUX2X1 U1618 ( .B(n1365), .A(n1362), .S(n1695), .Y(n1369) );
  MUX2X1 U1619 ( .B(n1368), .A(n1353), .S(n1687), .Y(n1676) );
  MUX2X1 U1620 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1712), .Y(n1373) );
  MUX2X1 U1621 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1712), .Y(n1372) );
  MUX2X1 U1622 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1712), .Y(n1376) );
  MUX2X1 U1623 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1712), .Y(n1375) );
  MUX2X1 U1624 ( .B(n1374), .A(n1371), .S(n1694), .Y(n1385) );
  MUX2X1 U1625 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1713), .Y(n1379) );
  MUX2X1 U1626 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1713), .Y(n1378) );
  MUX2X1 U1627 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1713), .Y(n1382) );
  MUX2X1 U1628 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1713), .Y(n1381) );
  MUX2X1 U1629 ( .B(n1380), .A(n1377), .S(n1694), .Y(n1384) );
  MUX2X1 U1630 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1713), .Y(n1388) );
  MUX2X1 U1631 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1713), .Y(n1387) );
  MUX2X1 U1632 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1713), .Y(n1391) );
  MUX2X1 U1633 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1713), .Y(n1390) );
  MUX2X1 U1634 ( .B(n1389), .A(n1386), .S(n1694), .Y(n1400) );
  MUX2X1 U1635 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1713), .Y(n1394) );
  MUX2X1 U1636 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1713), .Y(n1393) );
  MUX2X1 U1637 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1713), .Y(n1397) );
  MUX2X1 U1638 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1713), .Y(n1396) );
  MUX2X1 U1639 ( .B(n1395), .A(n1392), .S(n1694), .Y(n1399) );
  MUX2X1 U1640 ( .B(n1398), .A(n1383), .S(n1687), .Y(n1677) );
  MUX2X1 U1641 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1714), .Y(n1403) );
  MUX2X1 U1642 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1714), .Y(n1402) );
  MUX2X1 U1643 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1714), .Y(n1406) );
  MUX2X1 U1644 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1714), .Y(n1405) );
  MUX2X1 U1645 ( .B(n1404), .A(n1401), .S(n1694), .Y(n1415) );
  MUX2X1 U1646 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1714), .Y(n1409) );
  MUX2X1 U1647 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1714), .Y(n1408) );
  MUX2X1 U1648 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1714), .Y(n1412) );
  MUX2X1 U1649 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1714), .Y(n1411) );
  MUX2X1 U1650 ( .B(n1410), .A(n1407), .S(n1694), .Y(n1414) );
  MUX2X1 U1651 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1714), .Y(n1418) );
  MUX2X1 U1652 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1714), .Y(n1417) );
  MUX2X1 U1653 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1714), .Y(n1421) );
  MUX2X1 U1654 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1714), .Y(n1420) );
  MUX2X1 U1655 ( .B(n1419), .A(n1416), .S(n1694), .Y(n1430) );
  MUX2X1 U1656 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1715), .Y(n1424) );
  MUX2X1 U1657 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1715), .Y(n1423) );
  MUX2X1 U1658 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1715), .Y(n1427) );
  MUX2X1 U1659 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1715), .Y(n1426) );
  MUX2X1 U1660 ( .B(n1425), .A(n1422), .S(n1694), .Y(n1429) );
  MUX2X1 U1661 ( .B(n1428), .A(n1413), .S(n1687), .Y(n1678) );
  MUX2X1 U1662 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1715), .Y(n1433) );
  MUX2X1 U1663 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1715), .Y(n1432) );
  MUX2X1 U1664 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1715), .Y(n1436) );
  MUX2X1 U1665 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1715), .Y(n1435) );
  MUX2X1 U1666 ( .B(n1434), .A(n1431), .S(n1694), .Y(n1445) );
  MUX2X1 U1667 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1715), .Y(n1439) );
  MUX2X1 U1668 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1715), .Y(n1438) );
  MUX2X1 U1669 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1715), .Y(n1442) );
  MUX2X1 U1670 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1715), .Y(n1441) );
  MUX2X1 U1671 ( .B(n1440), .A(n1437), .S(n1694), .Y(n1444) );
  MUX2X1 U1672 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1716), .Y(n1448) );
  MUX2X1 U1673 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1716), .Y(n1447) );
  MUX2X1 U1674 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1716), .Y(n1451) );
  MUX2X1 U1675 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1716), .Y(n1450) );
  MUX2X1 U1676 ( .B(n1449), .A(n1446), .S(n1694), .Y(n1460) );
  MUX2X1 U1677 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1716), .Y(n1454) );
  MUX2X1 U1678 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1716), .Y(n1453) );
  MUX2X1 U1679 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1716), .Y(n1457) );
  MUX2X1 U1680 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1716), .Y(n1456) );
  MUX2X1 U1681 ( .B(n1455), .A(n1452), .S(n1694), .Y(n1459) );
  MUX2X1 U1682 ( .B(n1458), .A(n1443), .S(n1687), .Y(n1679) );
  MUX2X1 U1683 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1716), .Y(n1463) );
  MUX2X1 U1684 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1716), .Y(n1462) );
  MUX2X1 U1685 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1716), .Y(n1466) );
  MUX2X1 U1686 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1716), .Y(n1465) );
  MUX2X1 U1687 ( .B(n1464), .A(n1461), .S(n1693), .Y(n1475) );
  MUX2X1 U1688 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1717), .Y(n1469) );
  MUX2X1 U1689 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1717), .Y(n1468) );
  MUX2X1 U1690 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1717), .Y(n1472) );
  MUX2X1 U1691 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1717), .Y(n1471) );
  MUX2X1 U1692 ( .B(n1470), .A(n1467), .S(n1693), .Y(n1474) );
  MUX2X1 U1693 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1717), .Y(n1478) );
  MUX2X1 U1694 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1717), .Y(n1477) );
  MUX2X1 U1695 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1717), .Y(n1481) );
  MUX2X1 U1696 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1717), .Y(n1480) );
  MUX2X1 U1697 ( .B(n1479), .A(n1476), .S(n1693), .Y(n1490) );
  MUX2X1 U1698 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1717), .Y(n1484) );
  MUX2X1 U1699 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1717), .Y(n1483) );
  MUX2X1 U1700 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1717), .Y(n1487) );
  MUX2X1 U1701 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1717), .Y(n1486) );
  MUX2X1 U1702 ( .B(n1485), .A(n1482), .S(n1693), .Y(n1489) );
  MUX2X1 U1703 ( .B(n1488), .A(n1473), .S(n1687), .Y(n1680) );
  MUX2X1 U1704 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1718), .Y(n1493) );
  MUX2X1 U1705 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1718), .Y(n1492) );
  MUX2X1 U1706 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1718), .Y(n1496) );
  MUX2X1 U1707 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1718), .Y(n1495) );
  MUX2X1 U1708 ( .B(n1494), .A(n1491), .S(n1693), .Y(n1505) );
  MUX2X1 U1709 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1718), .Y(n1499) );
  MUX2X1 U1710 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1718), .Y(n1498) );
  MUX2X1 U1711 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1718), .Y(n1502) );
  MUX2X1 U1712 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1718), .Y(n1501) );
  MUX2X1 U1713 ( .B(n1500), .A(n1497), .S(n1693), .Y(n1504) );
  MUX2X1 U1714 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1718), .Y(n1508) );
  MUX2X1 U1715 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1718), .Y(n1507) );
  MUX2X1 U1716 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1718), .Y(n1511) );
  MUX2X1 U1717 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1718), .Y(n1510) );
  MUX2X1 U1718 ( .B(n1509), .A(n1506), .S(n1693), .Y(n1520) );
  MUX2X1 U1719 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1719), .Y(n1514) );
  MUX2X1 U1720 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1719), .Y(n1513) );
  MUX2X1 U1721 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1719), .Y(n1517) );
  MUX2X1 U1722 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1719), .Y(n1516) );
  MUX2X1 U1723 ( .B(n1515), .A(n1512), .S(n1693), .Y(n1519) );
  MUX2X1 U1724 ( .B(n1518), .A(n1503), .S(n1687), .Y(n1681) );
  MUX2X1 U1725 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1719), .Y(n1523) );
  MUX2X1 U1726 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1719), .Y(n1522) );
  MUX2X1 U1727 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1719), .Y(n1526) );
  MUX2X1 U1728 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1719), .Y(n1525) );
  MUX2X1 U1729 ( .B(n1524), .A(n1521), .S(n1693), .Y(n1535) );
  MUX2X1 U1730 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1719), .Y(n1529) );
  MUX2X1 U1731 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1719), .Y(n1528) );
  MUX2X1 U1732 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1719), .Y(n1532) );
  MUX2X1 U1733 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1719), .Y(n1531) );
  MUX2X1 U1734 ( .B(n1530), .A(n1527), .S(n1693), .Y(n1534) );
  MUX2X1 U1735 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1720), .Y(n1538) );
  MUX2X1 U1736 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1720), .Y(n1537) );
  MUX2X1 U1737 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1720), .Y(n1541) );
  MUX2X1 U1738 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1720), .Y(n1540) );
  MUX2X1 U1739 ( .B(n1539), .A(n1536), .S(n1693), .Y(n1550) );
  MUX2X1 U1740 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1720), .Y(n1544) );
  MUX2X1 U1741 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1720), .Y(n1543) );
  MUX2X1 U1742 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1720), .Y(n1547) );
  MUX2X1 U1743 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1720), .Y(n1546) );
  MUX2X1 U1744 ( .B(n1545), .A(n1542), .S(n1693), .Y(n1549) );
  MUX2X1 U1745 ( .B(n1548), .A(n1533), .S(n1687), .Y(n1682) );
  MUX2X1 U1746 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1720), .Y(n1553) );
  MUX2X1 U1747 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1720), .Y(n1552) );
  MUX2X1 U1748 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1720), .Y(n1556) );
  MUX2X1 U1749 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1720), .Y(n1555) );
  MUX2X1 U1750 ( .B(n1554), .A(n1551), .S(n1692), .Y(n1565) );
  MUX2X1 U1751 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1721), .Y(n1559) );
  MUX2X1 U1752 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1721), .Y(n1558) );
  MUX2X1 U1753 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1721), .Y(n1562) );
  MUX2X1 U1754 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1721), .Y(n1561) );
  MUX2X1 U1755 ( .B(n1560), .A(n1557), .S(n1692), .Y(n1564) );
  MUX2X1 U1756 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1721), .Y(n1568) );
  MUX2X1 U1757 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1721), .Y(n1567) );
  MUX2X1 U1758 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1721), .Y(n1571) );
  MUX2X1 U1759 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1721), .Y(n1570) );
  MUX2X1 U1760 ( .B(n1569), .A(n1566), .S(n1692), .Y(n1580) );
  MUX2X1 U1761 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1721), .Y(n1574) );
  MUX2X1 U1762 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1721), .Y(n1573) );
  MUX2X1 U1763 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1721), .Y(n1577) );
  MUX2X1 U1764 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1721), .Y(n1576) );
  MUX2X1 U1765 ( .B(n1575), .A(n1572), .S(n1692), .Y(n1579) );
  MUX2X1 U1766 ( .B(n1578), .A(n1563), .S(n1687), .Y(n1683) );
  MUX2X1 U1767 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1719), .Y(n1583) );
  MUX2X1 U1768 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1719), .Y(n1582) );
  MUX2X1 U1769 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1720), .Y(n1586) );
  MUX2X1 U1770 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1713), .Y(n1585) );
  MUX2X1 U1771 ( .B(n1584), .A(n1581), .S(n1692), .Y(n1595) );
  MUX2X1 U1772 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1720), .Y(n1589) );
  MUX2X1 U1773 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1713), .Y(n1588) );
  MUX2X1 U1774 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1715), .Y(n1592) );
  MUX2X1 U1775 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1715), .Y(n1591) );
  MUX2X1 U1776 ( .B(n1590), .A(n1587), .S(n1692), .Y(n1594) );
  MUX2X1 U1777 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1719), .Y(n1598) );
  MUX2X1 U1778 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1715), .Y(n1597) );
  MUX2X1 U1779 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1714), .Y(n1601) );
  MUX2X1 U1780 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1721), .Y(n1600) );
  MUX2X1 U1781 ( .B(n1599), .A(n1596), .S(n1692), .Y(n1610) );
  MUX2X1 U1782 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1722), .Y(n1604) );
  MUX2X1 U1783 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1722), .Y(n1603) );
  MUX2X1 U1784 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1722), .Y(n1607) );
  MUX2X1 U1785 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1722), .Y(n1606) );
  MUX2X1 U1786 ( .B(n1605), .A(n1602), .S(n1692), .Y(n1609) );
  MUX2X1 U1787 ( .B(n1608), .A(n1593), .S(n1687), .Y(n1684) );
  MUX2X1 U1788 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1722), .Y(n1613) );
  MUX2X1 U1789 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1722), .Y(n1612) );
  MUX2X1 U1790 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1722), .Y(n1616) );
  MUX2X1 U1791 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1722), .Y(n1615) );
  MUX2X1 U1792 ( .B(n1614), .A(n1611), .S(n1692), .Y(n1625) );
  MUX2X1 U1793 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1722), .Y(n1619) );
  MUX2X1 U1794 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1722), .Y(n1618) );
  MUX2X1 U1795 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1722), .Y(n1622) );
  MUX2X1 U1796 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1722), .Y(n1621) );
  MUX2X1 U1797 ( .B(n1620), .A(n1617), .S(n1692), .Y(n1624) );
  MUX2X1 U1798 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1723), .Y(n1628) );
  MUX2X1 U1799 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1723), .Y(n1627) );
  MUX2X1 U1800 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1723), .Y(n1631) );
  MUX2X1 U1801 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1723), .Y(n1630) );
  MUX2X1 U1802 ( .B(n1629), .A(n1626), .S(n1692), .Y(n1640) );
  MUX2X1 U1803 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1723), .Y(n1634) );
  MUX2X1 U1804 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1723), .Y(n1633) );
  MUX2X1 U1805 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1723), .Y(n1637) );
  MUX2X1 U1806 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1723), .Y(n1636) );
  MUX2X1 U1807 ( .B(n1635), .A(n1632), .S(n1692), .Y(n1639) );
  MUX2X1 U1808 ( .B(n1638), .A(n1623), .S(n1687), .Y(n1685) );
  MUX2X1 U1809 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1723), .Y(n1643) );
  MUX2X1 U1810 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1723), .Y(n1642) );
  MUX2X1 U1811 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1723), .Y(n1646) );
  MUX2X1 U1812 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1723), .Y(n1645) );
  MUX2X1 U1813 ( .B(n1644), .A(n1641), .S(n1691), .Y(n1655) );
  MUX2X1 U1814 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1724), .Y(n1649) );
  MUX2X1 U1815 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1724), .Y(n1648) );
  MUX2X1 U1816 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1724), .Y(n1652) );
  MUX2X1 U1817 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1724), .Y(n1651) );
  MUX2X1 U1818 ( .B(n1650), .A(n1647), .S(n1691), .Y(n1654) );
  MUX2X1 U1819 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1724), .Y(n1658) );
  MUX2X1 U1820 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1724), .Y(n1657) );
  MUX2X1 U1821 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1724), .Y(n1661) );
  MUX2X1 U1822 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1724), .Y(n1660) );
  MUX2X1 U1823 ( .B(n1659), .A(n1656), .S(n1691), .Y(n1670) );
  MUX2X1 U1824 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1724), .Y(n1664) );
  MUX2X1 U1825 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1724), .Y(n1663) );
  MUX2X1 U1826 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1724), .Y(n1667) );
  MUX2X1 U1827 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1724), .Y(n1666) );
  MUX2X1 U1828 ( .B(n1665), .A(n1662), .S(n1691), .Y(n1669) );
  MUX2X1 U1829 ( .B(n1668), .A(n1653), .S(n1687), .Y(n1686) );
  INVX8 U1830 ( .A(n1854), .Y(n1692) );
  INVX8 U1831 ( .A(n1854), .Y(n1693) );
  INVX8 U1832 ( .A(n1854), .Y(n1694) );
  INVX8 U1833 ( .A(n1854), .Y(n1695) );
  INVX8 U1834 ( .A(n1854), .Y(n1696) );
  INVX8 U1835 ( .A(n1710), .Y(n1719) );
  INVX1 U1836 ( .A(N11), .Y(n1853) );
  INVX8 U1837 ( .A(n1825), .Y(n1822) );
  INVX8 U1838 ( .A(n1825), .Y(n1823) );
  INVX8 U1839 ( .A(n1825), .Y(n1824) );
  INVX8 U1840 ( .A(n37), .Y(n1826) );
  INVX8 U1841 ( .A(n37), .Y(n1827) );
  INVX8 U1842 ( .A(n38), .Y(n1828) );
  INVX8 U1843 ( .A(n38), .Y(n1829) );
  INVX8 U1844 ( .A(n39), .Y(n1830) );
  INVX8 U1845 ( .A(n39), .Y(n1831) );
  INVX8 U1846 ( .A(n40), .Y(n1832) );
  INVX8 U1847 ( .A(n40), .Y(n1833) );
  INVX8 U1848 ( .A(n41), .Y(n1834) );
  INVX8 U1849 ( .A(n42), .Y(n1835) );
  INVX8 U1850 ( .A(n42), .Y(n1836) );
  INVX8 U1851 ( .A(n43), .Y(n1837) );
  INVX8 U1852 ( .A(n43), .Y(n1838) );
  INVX8 U1853 ( .A(n44), .Y(n1839) );
  INVX8 U1854 ( .A(n45), .Y(n1840) );
  INVX8 U1855 ( .A(n47), .Y(n1841) );
  INVX8 U1856 ( .A(n47), .Y(n1842) );
  INVX8 U1857 ( .A(n48), .Y(n1843) );
  INVX8 U1858 ( .A(n48), .Y(n1844) );
  INVX8 U1859 ( .A(n50), .Y(n1845) );
  INVX8 U1860 ( .A(n52), .Y(n1846) );
  INVX8 U1861 ( .A(n54), .Y(n1847) );
  INVX8 U1862 ( .A(n54), .Y(n1848) );
  INVX8 U1863 ( .A(n56), .Y(n1849) );
  INVX8 U1864 ( .A(n56), .Y(n1850) );
  INVX8 U1865 ( .A(n58), .Y(n1851) );
endmodule


module memc_Size16_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , n1, n2, n3, n5, n7, n9, n11, n13, n15, n17, n19, n21,
         n23, n25, n27, n29, n31, n33, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n47, n48, n50, n52, n54, n56, n58, n60, n62, n64, n66,
         n68, n70, n72, n74, n76, n80, n82, n99, n101, n118, n120, n137, n139,
         n156, n158, n175, n177, n194, n196, n215, n217, n233, n235, n251,
         n253, n269, n271, n287, n289, n305, n307, n323, n325, n341, n343,
         n360, n362, n378, n380, n396, n398, n414, n416, n432, n434, n450,
         n452, n468, n470, n486, n488, n505, n507, n523, n525, n541, n543,
         n559, n561, n577, n579, n595, n597, n613, n615, n631, n633, n650,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1856), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1857), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1858), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1859), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1860), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1861), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1862), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1863), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1864), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1865), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1866), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1867), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1868), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1869), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1870), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1871), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1872), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1873), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1874), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1875), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1876), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1877), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1878), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1879), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1880), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1881), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1882), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1883), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1884), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1885), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1886), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1887), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1888), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1889), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1890), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1891), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1892), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1893), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1894), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1895), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1896), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1897), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1898), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1899), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1900), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1901), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1902), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1903), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1904), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1905), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1906), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1907), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1908), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1909), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1910), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1911), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1912), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1913), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1914), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1915), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1916), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1917), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1918), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1919), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1920), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1921), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1922), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1923), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1924), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1925), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1926), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1927), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1928), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1929), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1930), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1931), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1932), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1933), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1934), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1935), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1936), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1937), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1938), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1939), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1940), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1941), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1942), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1943), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1944), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1945), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1946), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1947), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1948), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1949), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1950), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1951), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1952), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1953), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1954), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1955), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1956), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1957), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1958), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1959), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1960), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1961), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1962), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1963), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1964), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1965), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1966), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1967), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1968), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1969), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1970), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1971), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1972), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1973), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1974), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1975), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1976), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1977), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1978), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1979), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1980), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1981), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1982), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1983), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1984), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1985), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1986), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1987), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1988), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1989), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1990), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1991), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1992), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1993), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1994), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1995), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1996), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1997), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1998), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1999), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2000), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2001), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2002), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2003), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2004), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2005), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2006), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2007), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2008), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2009), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2010), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2011), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2012), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2013), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2014), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2015), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2016), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2017), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2018), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2019), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2020), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2021), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2022), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2023), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2024), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2025), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2026), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2027), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2028), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2029), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2030), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2031), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2032), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2033), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2034), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2035), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2036), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2037), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2038), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2039), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2040), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2041), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2042), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2043), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2044), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2045), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2046), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2047), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2048), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2049), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2050), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2051), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2052), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2053), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2054), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2055), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2056), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2057), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2058), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2059), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2060), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2061), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2062), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2063), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2064), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2065), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2066), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2067), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2068), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2069), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2070), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2071), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2072), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2073), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2074), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2075), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2076), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2077), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2078), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2079), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2080), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2081), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2082), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2083), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2084), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2085), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2086), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2087), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2088), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2089), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2090), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2091), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2092), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2093), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2094), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2095), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2096), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2097), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2098), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2099), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2100), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2101), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2102), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2103), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2104), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2105), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2106), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2107), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2108), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2109), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2110), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2111), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2112), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2113), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2114), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2115), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2116), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2117), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2118), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2119), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2120), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2121), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2122), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2123), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2124), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2125), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2126), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2127), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2128), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2129), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2130), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2131), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2132), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2133), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2134), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2135), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2136), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2137), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2138), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2139), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2140), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2141), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2142), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2143), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2144), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2145), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2146), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2147), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2148), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2149), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2150), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2151), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2152), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2153), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2154), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2155), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2156), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2157), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2158), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2159), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2160), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2161), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2162), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2163), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2164), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2165), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2166), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2167), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2168), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2169), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2170), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2171), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2172), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2173), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2174), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2175), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2176), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2177), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2178), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2179), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2180), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2181), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2182), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2183), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2184), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2185), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2186), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2187), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2188), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2189), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2190), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2191), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2192), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2193), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2194), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2195), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2196), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2197), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2198), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2199), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2200), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2201), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2202), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2203), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2204), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2205), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2206), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2207), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2208), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2209), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2210), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2211), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2212), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2213), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2214), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2215), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2216), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2217), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2218), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2219), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2220), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2221), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2222), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2223), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2224), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2225), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2226), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2227), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2228), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2229), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2230), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2231), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2232), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2233), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2234), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2235), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2236), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2237), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2238), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2239), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2240), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2241), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2242), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2243), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2244), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2245), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2246), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2247), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2248), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2249), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2250), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2251), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2252), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2253), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2254), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2255), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2256), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2257), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2258), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2259), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2260), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2261), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2262), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2263), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2264), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2265), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2266), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2267), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2268), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2269), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2270), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2271), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2272), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2273), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2274), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2275), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2276), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2277), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2278), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2279), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2280), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2281), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2282), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2283), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2284), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2285), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2286), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2287), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2288), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2289), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2290), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2291), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2292), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2293), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2294), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2295), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2296), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2297), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2298), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2299), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2300), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2301), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2302), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2303), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2304), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2305), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2306), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2307), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2308), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2309), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2310), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2311), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2312), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2313), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2314), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2315), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2316), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2317), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2318), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2319), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2320), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2321), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2322), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2323), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2324), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2325), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2326), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2327), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2328), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2329), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2330), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2331), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2332), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2333), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2334), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2335), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2336), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2337), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2338), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2339), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2340), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2341), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2342), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2343), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2344), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2345), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2346), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2347), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2348), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2349), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2350), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2351), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2352), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2353), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2354), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2355), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2356), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2357), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2358), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2359), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2360), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2361), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2362), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2363), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2364), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2365), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2366), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2367), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(write), .B(n1850), .Y(n2877) );
  OAI21X1 U61 ( .A(n1818), .B(n1840), .C(n2893), .Y(n2367) );
  NAND2X1 U62 ( .A(\mem<31><0> ), .B(n1820), .Y(n2893) );
  OAI21X1 U63 ( .A(n1818), .B(n1839), .C(n2892), .Y(n2366) );
  NAND2X1 U64 ( .A(\mem<31><1> ), .B(n1820), .Y(n2892) );
  OAI21X1 U65 ( .A(n1818), .B(n1838), .C(n2891), .Y(n2365) );
  NAND2X1 U66 ( .A(\mem<31><2> ), .B(n1820), .Y(n2891) );
  OAI21X1 U67 ( .A(n1818), .B(n1837), .C(n2890), .Y(n2364) );
  NAND2X1 U68 ( .A(\mem<31><3> ), .B(n1820), .Y(n2890) );
  OAI21X1 U69 ( .A(n1818), .B(n1836), .C(n2889), .Y(n2363) );
  NAND2X1 U70 ( .A(\mem<31><4> ), .B(n1820), .Y(n2889) );
  OAI21X1 U71 ( .A(n1818), .B(n1835), .C(n2888), .Y(n2362) );
  NAND2X1 U72 ( .A(\mem<31><5> ), .B(n1820), .Y(n2888) );
  OAI21X1 U73 ( .A(n1818), .B(n1834), .C(n2887), .Y(n2361) );
  NAND2X1 U74 ( .A(\mem<31><6> ), .B(n1820), .Y(n2887) );
  OAI21X1 U75 ( .A(n1818), .B(n1833), .C(n2886), .Y(n2360) );
  NAND2X1 U76 ( .A(\mem<31><7> ), .B(n1820), .Y(n2886) );
  OAI21X1 U77 ( .A(n1818), .B(n1832), .C(n2885), .Y(n2359) );
  NAND2X1 U78 ( .A(\mem<31><8> ), .B(n1819), .Y(n2885) );
  OAI21X1 U79 ( .A(n1818), .B(n1831), .C(n2884), .Y(n2358) );
  NAND2X1 U80 ( .A(\mem<31><9> ), .B(n1819), .Y(n2884) );
  OAI21X1 U81 ( .A(n1818), .B(n1830), .C(n2883), .Y(n2357) );
  NAND2X1 U82 ( .A(\mem<31><10> ), .B(n1819), .Y(n2883) );
  OAI21X1 U83 ( .A(n1818), .B(n1829), .C(n2882), .Y(n2356) );
  NAND2X1 U84 ( .A(\mem<31><11> ), .B(n1819), .Y(n2882) );
  OAI21X1 U85 ( .A(n1818), .B(n1828), .C(n2881), .Y(n2355) );
  NAND2X1 U86 ( .A(\mem<31><12> ), .B(n1819), .Y(n2881) );
  OAI21X1 U87 ( .A(n1818), .B(n1827), .C(n2880), .Y(n2354) );
  NAND2X1 U88 ( .A(\mem<31><13> ), .B(n1819), .Y(n2880) );
  OAI21X1 U89 ( .A(n1818), .B(n1826), .C(n2879), .Y(n2353) );
  NAND2X1 U90 ( .A(\mem<31><14> ), .B(n1819), .Y(n2879) );
  OAI21X1 U91 ( .A(n1818), .B(n1825), .C(n2878), .Y(n2352) );
  NAND2X1 U92 ( .A(\mem<31><15> ), .B(n1819), .Y(n2878) );
  OAI21X1 U95 ( .A(n1840), .B(n1815), .C(n2875), .Y(n2351) );
  NAND2X1 U96 ( .A(\mem<30><0> ), .B(n1817), .Y(n2875) );
  OAI21X1 U97 ( .A(n1839), .B(n1815), .C(n2874), .Y(n2350) );
  NAND2X1 U98 ( .A(\mem<30><1> ), .B(n1817), .Y(n2874) );
  OAI21X1 U99 ( .A(n1838), .B(n1815), .C(n2873), .Y(n2349) );
  NAND2X1 U100 ( .A(\mem<30><2> ), .B(n1817), .Y(n2873) );
  OAI21X1 U101 ( .A(n1837), .B(n1815), .C(n2872), .Y(n2348) );
  NAND2X1 U102 ( .A(\mem<30><3> ), .B(n1817), .Y(n2872) );
  OAI21X1 U103 ( .A(n1836), .B(n1815), .C(n2871), .Y(n2347) );
  NAND2X1 U104 ( .A(\mem<30><4> ), .B(n1817), .Y(n2871) );
  OAI21X1 U105 ( .A(n1835), .B(n1815), .C(n2870), .Y(n2346) );
  NAND2X1 U106 ( .A(\mem<30><5> ), .B(n1817), .Y(n2870) );
  OAI21X1 U107 ( .A(n1834), .B(n1815), .C(n2869), .Y(n2345) );
  NAND2X1 U108 ( .A(\mem<30><6> ), .B(n1817), .Y(n2869) );
  OAI21X1 U109 ( .A(n1833), .B(n1815), .C(n2868), .Y(n2344) );
  NAND2X1 U110 ( .A(\mem<30><7> ), .B(n1817), .Y(n2868) );
  OAI21X1 U111 ( .A(n1832), .B(n1815), .C(n2867), .Y(n2343) );
  NAND2X1 U112 ( .A(\mem<30><8> ), .B(n1816), .Y(n2867) );
  OAI21X1 U113 ( .A(n1831), .B(n1815), .C(n2866), .Y(n2342) );
  NAND2X1 U114 ( .A(\mem<30><9> ), .B(n1816), .Y(n2866) );
  OAI21X1 U115 ( .A(n1830), .B(n1815), .C(n2865), .Y(n2341) );
  NAND2X1 U116 ( .A(\mem<30><10> ), .B(n1816), .Y(n2865) );
  OAI21X1 U117 ( .A(n1829), .B(n1815), .C(n2864), .Y(n2340) );
  NAND2X1 U118 ( .A(\mem<30><11> ), .B(n1816), .Y(n2864) );
  OAI21X1 U119 ( .A(n1828), .B(n1815), .C(n2863), .Y(n2339) );
  NAND2X1 U120 ( .A(\mem<30><12> ), .B(n1816), .Y(n2863) );
  OAI21X1 U121 ( .A(n1827), .B(n1815), .C(n2862), .Y(n2338) );
  NAND2X1 U122 ( .A(\mem<30><13> ), .B(n1816), .Y(n2862) );
  OAI21X1 U123 ( .A(n1826), .B(n1815), .C(n2861), .Y(n2337) );
  NAND2X1 U124 ( .A(\mem<30><14> ), .B(n1816), .Y(n2861) );
  OAI21X1 U125 ( .A(n1825), .B(n1815), .C(n2860), .Y(n2336) );
  NAND2X1 U126 ( .A(\mem<30><15> ), .B(n1816), .Y(n2860) );
  OAI21X1 U129 ( .A(n1840), .B(n1812), .C(n2858), .Y(n2335) );
  NAND2X1 U130 ( .A(\mem<29><0> ), .B(n1814), .Y(n2858) );
  OAI21X1 U131 ( .A(n1839), .B(n1812), .C(n2857), .Y(n2334) );
  NAND2X1 U132 ( .A(\mem<29><1> ), .B(n1814), .Y(n2857) );
  OAI21X1 U133 ( .A(n1838), .B(n1812), .C(n2856), .Y(n2333) );
  NAND2X1 U134 ( .A(\mem<29><2> ), .B(n1814), .Y(n2856) );
  OAI21X1 U135 ( .A(n1837), .B(n1812), .C(n2855), .Y(n2332) );
  NAND2X1 U136 ( .A(\mem<29><3> ), .B(n1814), .Y(n2855) );
  OAI21X1 U137 ( .A(n1836), .B(n1812), .C(n2854), .Y(n2331) );
  NAND2X1 U138 ( .A(\mem<29><4> ), .B(n1814), .Y(n2854) );
  OAI21X1 U139 ( .A(n1835), .B(n1812), .C(n2853), .Y(n2330) );
  NAND2X1 U140 ( .A(\mem<29><5> ), .B(n1814), .Y(n2853) );
  OAI21X1 U141 ( .A(n1834), .B(n1812), .C(n2852), .Y(n2329) );
  NAND2X1 U142 ( .A(\mem<29><6> ), .B(n1814), .Y(n2852) );
  OAI21X1 U143 ( .A(n1833), .B(n1812), .C(n2851), .Y(n2328) );
  NAND2X1 U144 ( .A(\mem<29><7> ), .B(n1814), .Y(n2851) );
  OAI21X1 U145 ( .A(n1832), .B(n1812), .C(n2850), .Y(n2327) );
  NAND2X1 U146 ( .A(\mem<29><8> ), .B(n1813), .Y(n2850) );
  OAI21X1 U147 ( .A(n1831), .B(n1812), .C(n2849), .Y(n2326) );
  NAND2X1 U148 ( .A(\mem<29><9> ), .B(n1813), .Y(n2849) );
  OAI21X1 U149 ( .A(n1830), .B(n1812), .C(n2848), .Y(n2325) );
  NAND2X1 U150 ( .A(\mem<29><10> ), .B(n1813), .Y(n2848) );
  OAI21X1 U151 ( .A(n1829), .B(n1812), .C(n2847), .Y(n2324) );
  NAND2X1 U152 ( .A(\mem<29><11> ), .B(n1813), .Y(n2847) );
  OAI21X1 U153 ( .A(n1828), .B(n1812), .C(n2846), .Y(n2323) );
  NAND2X1 U154 ( .A(\mem<29><12> ), .B(n1813), .Y(n2846) );
  OAI21X1 U155 ( .A(n1827), .B(n1812), .C(n2845), .Y(n2322) );
  NAND2X1 U156 ( .A(\mem<29><13> ), .B(n1813), .Y(n2845) );
  OAI21X1 U157 ( .A(n1826), .B(n1812), .C(n2844), .Y(n2321) );
  NAND2X1 U158 ( .A(\mem<29><14> ), .B(n1813), .Y(n2844) );
  OAI21X1 U159 ( .A(n1825), .B(n1812), .C(n2843), .Y(n2320) );
  NAND2X1 U160 ( .A(\mem<29><15> ), .B(n1813), .Y(n2843) );
  OAI21X1 U163 ( .A(n1840), .B(n1809), .C(n2841), .Y(n2319) );
  NAND2X1 U164 ( .A(\mem<28><0> ), .B(n1811), .Y(n2841) );
  OAI21X1 U165 ( .A(n1839), .B(n1809), .C(n2840), .Y(n2318) );
  NAND2X1 U166 ( .A(\mem<28><1> ), .B(n1811), .Y(n2840) );
  OAI21X1 U167 ( .A(n1838), .B(n1809), .C(n2839), .Y(n2317) );
  NAND2X1 U168 ( .A(\mem<28><2> ), .B(n1811), .Y(n2839) );
  OAI21X1 U169 ( .A(n1837), .B(n1809), .C(n2838), .Y(n2316) );
  NAND2X1 U170 ( .A(\mem<28><3> ), .B(n1811), .Y(n2838) );
  OAI21X1 U171 ( .A(n1836), .B(n1809), .C(n2837), .Y(n2315) );
  NAND2X1 U172 ( .A(\mem<28><4> ), .B(n1811), .Y(n2837) );
  OAI21X1 U173 ( .A(n1835), .B(n1809), .C(n2836), .Y(n2314) );
  NAND2X1 U174 ( .A(\mem<28><5> ), .B(n1811), .Y(n2836) );
  OAI21X1 U175 ( .A(n1834), .B(n1809), .C(n2835), .Y(n2313) );
  NAND2X1 U176 ( .A(\mem<28><6> ), .B(n1811), .Y(n2835) );
  OAI21X1 U177 ( .A(n1833), .B(n1809), .C(n2834), .Y(n2312) );
  NAND2X1 U178 ( .A(\mem<28><7> ), .B(n1811), .Y(n2834) );
  OAI21X1 U179 ( .A(n1832), .B(n1809), .C(n2833), .Y(n2311) );
  NAND2X1 U180 ( .A(\mem<28><8> ), .B(n1810), .Y(n2833) );
  OAI21X1 U181 ( .A(n1831), .B(n1809), .C(n2832), .Y(n2310) );
  NAND2X1 U182 ( .A(\mem<28><9> ), .B(n1810), .Y(n2832) );
  OAI21X1 U183 ( .A(n1830), .B(n1809), .C(n2831), .Y(n2309) );
  NAND2X1 U184 ( .A(\mem<28><10> ), .B(n1810), .Y(n2831) );
  OAI21X1 U185 ( .A(n1829), .B(n1809), .C(n2830), .Y(n2308) );
  NAND2X1 U186 ( .A(\mem<28><11> ), .B(n1810), .Y(n2830) );
  OAI21X1 U187 ( .A(n1828), .B(n1809), .C(n2829), .Y(n2307) );
  NAND2X1 U188 ( .A(\mem<28><12> ), .B(n1810), .Y(n2829) );
  OAI21X1 U189 ( .A(n1827), .B(n1809), .C(n2828), .Y(n2306) );
  NAND2X1 U190 ( .A(\mem<28><13> ), .B(n1810), .Y(n2828) );
  OAI21X1 U191 ( .A(n1826), .B(n1809), .C(n2827), .Y(n2305) );
  NAND2X1 U192 ( .A(\mem<28><14> ), .B(n1810), .Y(n2827) );
  OAI21X1 U193 ( .A(n1825), .B(n1809), .C(n2826), .Y(n2304) );
  NAND2X1 U194 ( .A(\mem<28><15> ), .B(n1810), .Y(n2826) );
  OAI21X1 U197 ( .A(n1840), .B(n1806), .C(n2824), .Y(n2303) );
  NAND2X1 U198 ( .A(\mem<27><0> ), .B(n1808), .Y(n2824) );
  OAI21X1 U199 ( .A(n1839), .B(n1806), .C(n2823), .Y(n2302) );
  NAND2X1 U200 ( .A(\mem<27><1> ), .B(n1808), .Y(n2823) );
  OAI21X1 U201 ( .A(n1838), .B(n1806), .C(n2822), .Y(n2301) );
  NAND2X1 U202 ( .A(\mem<27><2> ), .B(n1808), .Y(n2822) );
  OAI21X1 U203 ( .A(n1837), .B(n1806), .C(n2821), .Y(n2300) );
  NAND2X1 U204 ( .A(\mem<27><3> ), .B(n1808), .Y(n2821) );
  OAI21X1 U205 ( .A(n1836), .B(n1806), .C(n2820), .Y(n2299) );
  NAND2X1 U206 ( .A(\mem<27><4> ), .B(n1808), .Y(n2820) );
  OAI21X1 U207 ( .A(n1835), .B(n1806), .C(n2819), .Y(n2298) );
  NAND2X1 U208 ( .A(\mem<27><5> ), .B(n1808), .Y(n2819) );
  OAI21X1 U209 ( .A(n1834), .B(n1806), .C(n2818), .Y(n2297) );
  NAND2X1 U210 ( .A(\mem<27><6> ), .B(n1808), .Y(n2818) );
  OAI21X1 U211 ( .A(n1833), .B(n1806), .C(n2817), .Y(n2296) );
  NAND2X1 U212 ( .A(\mem<27><7> ), .B(n1808), .Y(n2817) );
  OAI21X1 U213 ( .A(n1832), .B(n1806), .C(n2816), .Y(n2295) );
  NAND2X1 U214 ( .A(\mem<27><8> ), .B(n1807), .Y(n2816) );
  OAI21X1 U215 ( .A(n1831), .B(n1806), .C(n2815), .Y(n2294) );
  NAND2X1 U216 ( .A(\mem<27><9> ), .B(n1807), .Y(n2815) );
  OAI21X1 U217 ( .A(n1830), .B(n1806), .C(n2814), .Y(n2293) );
  NAND2X1 U218 ( .A(\mem<27><10> ), .B(n1807), .Y(n2814) );
  OAI21X1 U219 ( .A(n1829), .B(n1806), .C(n2813), .Y(n2292) );
  NAND2X1 U220 ( .A(\mem<27><11> ), .B(n1807), .Y(n2813) );
  OAI21X1 U221 ( .A(n1828), .B(n1806), .C(n2812), .Y(n2291) );
  NAND2X1 U222 ( .A(\mem<27><12> ), .B(n1807), .Y(n2812) );
  OAI21X1 U223 ( .A(n1827), .B(n1806), .C(n2811), .Y(n2290) );
  NAND2X1 U224 ( .A(\mem<27><13> ), .B(n1807), .Y(n2811) );
  OAI21X1 U225 ( .A(n1826), .B(n1806), .C(n2810), .Y(n2289) );
  NAND2X1 U226 ( .A(\mem<27><14> ), .B(n1807), .Y(n2810) );
  OAI21X1 U227 ( .A(n1825), .B(n1806), .C(n2809), .Y(n2288) );
  NAND2X1 U228 ( .A(\mem<27><15> ), .B(n1807), .Y(n2809) );
  OAI21X1 U231 ( .A(n1840), .B(n1803), .C(n2807), .Y(n2287) );
  NAND2X1 U232 ( .A(\mem<26><0> ), .B(n1805), .Y(n2807) );
  OAI21X1 U233 ( .A(n1839), .B(n1803), .C(n2806), .Y(n2286) );
  NAND2X1 U234 ( .A(\mem<26><1> ), .B(n1805), .Y(n2806) );
  OAI21X1 U235 ( .A(n1838), .B(n1803), .C(n2805), .Y(n2285) );
  NAND2X1 U236 ( .A(\mem<26><2> ), .B(n1805), .Y(n2805) );
  OAI21X1 U237 ( .A(n1837), .B(n1803), .C(n2804), .Y(n2284) );
  NAND2X1 U238 ( .A(\mem<26><3> ), .B(n1805), .Y(n2804) );
  OAI21X1 U239 ( .A(n1836), .B(n1803), .C(n2803), .Y(n2283) );
  NAND2X1 U240 ( .A(\mem<26><4> ), .B(n1805), .Y(n2803) );
  OAI21X1 U241 ( .A(n1835), .B(n1803), .C(n2802), .Y(n2282) );
  NAND2X1 U242 ( .A(\mem<26><5> ), .B(n1805), .Y(n2802) );
  OAI21X1 U243 ( .A(n1834), .B(n1803), .C(n2801), .Y(n2281) );
  NAND2X1 U244 ( .A(\mem<26><6> ), .B(n1805), .Y(n2801) );
  OAI21X1 U245 ( .A(n1833), .B(n1803), .C(n2800), .Y(n2280) );
  NAND2X1 U246 ( .A(\mem<26><7> ), .B(n1805), .Y(n2800) );
  OAI21X1 U247 ( .A(n1832), .B(n1803), .C(n2799), .Y(n2279) );
  NAND2X1 U248 ( .A(\mem<26><8> ), .B(n1804), .Y(n2799) );
  OAI21X1 U249 ( .A(n1831), .B(n1803), .C(n2798), .Y(n2278) );
  NAND2X1 U250 ( .A(\mem<26><9> ), .B(n1804), .Y(n2798) );
  OAI21X1 U251 ( .A(n1830), .B(n1803), .C(n2797), .Y(n2277) );
  NAND2X1 U252 ( .A(\mem<26><10> ), .B(n1804), .Y(n2797) );
  OAI21X1 U253 ( .A(n1829), .B(n1803), .C(n2796), .Y(n2276) );
  NAND2X1 U254 ( .A(\mem<26><11> ), .B(n1804), .Y(n2796) );
  OAI21X1 U255 ( .A(n1828), .B(n1803), .C(n2795), .Y(n2275) );
  NAND2X1 U256 ( .A(\mem<26><12> ), .B(n1804), .Y(n2795) );
  OAI21X1 U257 ( .A(n1827), .B(n1803), .C(n2794), .Y(n2274) );
  NAND2X1 U258 ( .A(\mem<26><13> ), .B(n1804), .Y(n2794) );
  OAI21X1 U259 ( .A(n1826), .B(n1803), .C(n2793), .Y(n2273) );
  NAND2X1 U260 ( .A(\mem<26><14> ), .B(n1804), .Y(n2793) );
  OAI21X1 U261 ( .A(n1825), .B(n1803), .C(n2792), .Y(n2272) );
  NAND2X1 U262 ( .A(\mem<26><15> ), .B(n1804), .Y(n2792) );
  OAI21X1 U265 ( .A(n1840), .B(n1800), .C(n2790), .Y(n2271) );
  NAND2X1 U266 ( .A(\mem<25><0> ), .B(n1802), .Y(n2790) );
  OAI21X1 U267 ( .A(n1839), .B(n1800), .C(n2789), .Y(n2270) );
  NAND2X1 U268 ( .A(\mem<25><1> ), .B(n1802), .Y(n2789) );
  OAI21X1 U269 ( .A(n1838), .B(n1800), .C(n2788), .Y(n2269) );
  NAND2X1 U270 ( .A(\mem<25><2> ), .B(n1802), .Y(n2788) );
  OAI21X1 U271 ( .A(n1837), .B(n1800), .C(n2787), .Y(n2268) );
  NAND2X1 U272 ( .A(\mem<25><3> ), .B(n1802), .Y(n2787) );
  OAI21X1 U273 ( .A(n1836), .B(n1800), .C(n2786), .Y(n2267) );
  NAND2X1 U274 ( .A(\mem<25><4> ), .B(n1802), .Y(n2786) );
  OAI21X1 U275 ( .A(n1835), .B(n1800), .C(n2785), .Y(n2266) );
  NAND2X1 U276 ( .A(\mem<25><5> ), .B(n1802), .Y(n2785) );
  OAI21X1 U277 ( .A(n1834), .B(n1800), .C(n2784), .Y(n2265) );
  NAND2X1 U278 ( .A(\mem<25><6> ), .B(n1802), .Y(n2784) );
  OAI21X1 U279 ( .A(n1833), .B(n1800), .C(n2783), .Y(n2264) );
  NAND2X1 U280 ( .A(\mem<25><7> ), .B(n1802), .Y(n2783) );
  OAI21X1 U281 ( .A(n1832), .B(n1800), .C(n2782), .Y(n2263) );
  NAND2X1 U282 ( .A(\mem<25><8> ), .B(n1801), .Y(n2782) );
  OAI21X1 U283 ( .A(n1831), .B(n1800), .C(n2781), .Y(n2262) );
  NAND2X1 U284 ( .A(\mem<25><9> ), .B(n1801), .Y(n2781) );
  OAI21X1 U285 ( .A(n1830), .B(n1800), .C(n2780), .Y(n2261) );
  NAND2X1 U286 ( .A(\mem<25><10> ), .B(n1801), .Y(n2780) );
  OAI21X1 U287 ( .A(n1829), .B(n1800), .C(n2779), .Y(n2260) );
  NAND2X1 U288 ( .A(\mem<25><11> ), .B(n1801), .Y(n2779) );
  OAI21X1 U289 ( .A(n1828), .B(n1800), .C(n2778), .Y(n2259) );
  NAND2X1 U290 ( .A(\mem<25><12> ), .B(n1801), .Y(n2778) );
  OAI21X1 U291 ( .A(n1827), .B(n1800), .C(n2777), .Y(n2258) );
  NAND2X1 U292 ( .A(\mem<25><13> ), .B(n1801), .Y(n2777) );
  OAI21X1 U293 ( .A(n1826), .B(n1800), .C(n2776), .Y(n2257) );
  NAND2X1 U294 ( .A(\mem<25><14> ), .B(n1801), .Y(n2776) );
  OAI21X1 U295 ( .A(n1825), .B(n1800), .C(n2775), .Y(n2256) );
  NAND2X1 U296 ( .A(\mem<25><15> ), .B(n1801), .Y(n2775) );
  OAI21X1 U299 ( .A(n1840), .B(n1797), .C(n2773), .Y(n2255) );
  NAND2X1 U300 ( .A(\mem<24><0> ), .B(n1799), .Y(n2773) );
  OAI21X1 U301 ( .A(n1839), .B(n1797), .C(n2772), .Y(n2254) );
  NAND2X1 U302 ( .A(\mem<24><1> ), .B(n1799), .Y(n2772) );
  OAI21X1 U303 ( .A(n1838), .B(n1797), .C(n2771), .Y(n2253) );
  NAND2X1 U304 ( .A(\mem<24><2> ), .B(n1799), .Y(n2771) );
  OAI21X1 U305 ( .A(n1837), .B(n1797), .C(n2770), .Y(n2252) );
  NAND2X1 U306 ( .A(\mem<24><3> ), .B(n1799), .Y(n2770) );
  OAI21X1 U307 ( .A(n1836), .B(n1797), .C(n2769), .Y(n2251) );
  NAND2X1 U308 ( .A(\mem<24><4> ), .B(n1799), .Y(n2769) );
  OAI21X1 U309 ( .A(n1835), .B(n1797), .C(n2768), .Y(n2250) );
  NAND2X1 U310 ( .A(\mem<24><5> ), .B(n1799), .Y(n2768) );
  OAI21X1 U311 ( .A(n1834), .B(n1797), .C(n2767), .Y(n2249) );
  NAND2X1 U312 ( .A(\mem<24><6> ), .B(n1799), .Y(n2767) );
  OAI21X1 U313 ( .A(n1833), .B(n1797), .C(n2766), .Y(n2248) );
  NAND2X1 U314 ( .A(\mem<24><7> ), .B(n1799), .Y(n2766) );
  OAI21X1 U315 ( .A(n1832), .B(n1797), .C(n2765), .Y(n2247) );
  NAND2X1 U316 ( .A(\mem<24><8> ), .B(n1798), .Y(n2765) );
  OAI21X1 U317 ( .A(n1831), .B(n1797), .C(n2764), .Y(n2246) );
  NAND2X1 U318 ( .A(\mem<24><9> ), .B(n1798), .Y(n2764) );
  OAI21X1 U319 ( .A(n1830), .B(n1797), .C(n2763), .Y(n2245) );
  NAND2X1 U320 ( .A(\mem<24><10> ), .B(n1798), .Y(n2763) );
  OAI21X1 U321 ( .A(n1829), .B(n1797), .C(n2762), .Y(n2244) );
  NAND2X1 U322 ( .A(\mem<24><11> ), .B(n1798), .Y(n2762) );
  OAI21X1 U323 ( .A(n1828), .B(n1797), .C(n2761), .Y(n2243) );
  NAND2X1 U324 ( .A(\mem<24><12> ), .B(n1798), .Y(n2761) );
  OAI21X1 U325 ( .A(n1827), .B(n1797), .C(n2760), .Y(n2242) );
  NAND2X1 U326 ( .A(\mem<24><13> ), .B(n1798), .Y(n2760) );
  OAI21X1 U327 ( .A(n1826), .B(n1797), .C(n2759), .Y(n2241) );
  NAND2X1 U328 ( .A(\mem<24><14> ), .B(n1798), .Y(n2759) );
  OAI21X1 U329 ( .A(n1825), .B(n1797), .C(n2758), .Y(n2240) );
  NAND2X1 U330 ( .A(\mem<24><15> ), .B(n1798), .Y(n2758) );
  NAND3X1 U333 ( .A(n1846), .B(n2755), .C(n1848), .Y(n2756) );
  OAI21X1 U334 ( .A(n1840), .B(n1794), .C(n2754), .Y(n2239) );
  NAND2X1 U335 ( .A(\mem<23><0> ), .B(n1796), .Y(n2754) );
  OAI21X1 U336 ( .A(n1839), .B(n1794), .C(n2753), .Y(n2238) );
  NAND2X1 U337 ( .A(\mem<23><1> ), .B(n1796), .Y(n2753) );
  OAI21X1 U338 ( .A(n1838), .B(n1794), .C(n2752), .Y(n2237) );
  NAND2X1 U339 ( .A(\mem<23><2> ), .B(n1796), .Y(n2752) );
  OAI21X1 U340 ( .A(n1837), .B(n1794), .C(n2751), .Y(n2236) );
  NAND2X1 U341 ( .A(\mem<23><3> ), .B(n1796), .Y(n2751) );
  OAI21X1 U342 ( .A(n1836), .B(n1794), .C(n2750), .Y(n2235) );
  NAND2X1 U343 ( .A(\mem<23><4> ), .B(n1796), .Y(n2750) );
  OAI21X1 U344 ( .A(n1835), .B(n1794), .C(n2749), .Y(n2234) );
  NAND2X1 U345 ( .A(\mem<23><5> ), .B(n1796), .Y(n2749) );
  OAI21X1 U346 ( .A(n1834), .B(n1794), .C(n2748), .Y(n2233) );
  NAND2X1 U347 ( .A(\mem<23><6> ), .B(n1796), .Y(n2748) );
  OAI21X1 U348 ( .A(n1833), .B(n1794), .C(n2747), .Y(n2232) );
  NAND2X1 U349 ( .A(\mem<23><7> ), .B(n1796), .Y(n2747) );
  OAI21X1 U350 ( .A(n1832), .B(n1794), .C(n2746), .Y(n2231) );
  NAND2X1 U351 ( .A(\mem<23><8> ), .B(n1795), .Y(n2746) );
  OAI21X1 U352 ( .A(n1831), .B(n1794), .C(n2745), .Y(n2230) );
  NAND2X1 U353 ( .A(\mem<23><9> ), .B(n1795), .Y(n2745) );
  OAI21X1 U354 ( .A(n1830), .B(n1794), .C(n2744), .Y(n2229) );
  NAND2X1 U355 ( .A(\mem<23><10> ), .B(n1795), .Y(n2744) );
  OAI21X1 U356 ( .A(n1829), .B(n1794), .C(n2743), .Y(n2228) );
  NAND2X1 U357 ( .A(\mem<23><11> ), .B(n1795), .Y(n2743) );
  OAI21X1 U358 ( .A(n1828), .B(n1794), .C(n2742), .Y(n2227) );
  NAND2X1 U359 ( .A(\mem<23><12> ), .B(n1795), .Y(n2742) );
  OAI21X1 U360 ( .A(n1827), .B(n1794), .C(n2741), .Y(n2226) );
  NAND2X1 U361 ( .A(\mem<23><13> ), .B(n1795), .Y(n2741) );
  OAI21X1 U362 ( .A(n1826), .B(n1794), .C(n2740), .Y(n2225) );
  NAND2X1 U363 ( .A(\mem<23><14> ), .B(n1795), .Y(n2740) );
  OAI21X1 U364 ( .A(n1825), .B(n1794), .C(n2739), .Y(n2224) );
  NAND2X1 U365 ( .A(\mem<23><15> ), .B(n1795), .Y(n2739) );
  OAI21X1 U368 ( .A(n1840), .B(n1791), .C(n2738), .Y(n2223) );
  NAND2X1 U369 ( .A(\mem<22><0> ), .B(n1793), .Y(n2738) );
  OAI21X1 U370 ( .A(n1839), .B(n1791), .C(n2737), .Y(n2222) );
  NAND2X1 U371 ( .A(\mem<22><1> ), .B(n1793), .Y(n2737) );
  OAI21X1 U372 ( .A(n1838), .B(n1791), .C(n2736), .Y(n2221) );
  NAND2X1 U373 ( .A(\mem<22><2> ), .B(n1793), .Y(n2736) );
  OAI21X1 U374 ( .A(n1837), .B(n1791), .C(n2735), .Y(n2220) );
  NAND2X1 U375 ( .A(\mem<22><3> ), .B(n1793), .Y(n2735) );
  OAI21X1 U376 ( .A(n1836), .B(n1791), .C(n2734), .Y(n2219) );
  NAND2X1 U377 ( .A(\mem<22><4> ), .B(n1793), .Y(n2734) );
  OAI21X1 U378 ( .A(n1835), .B(n1791), .C(n2733), .Y(n2218) );
  NAND2X1 U379 ( .A(\mem<22><5> ), .B(n1793), .Y(n2733) );
  OAI21X1 U380 ( .A(n1834), .B(n1791), .C(n2732), .Y(n2217) );
  NAND2X1 U381 ( .A(\mem<22><6> ), .B(n1793), .Y(n2732) );
  OAI21X1 U382 ( .A(n1833), .B(n1791), .C(n2731), .Y(n2216) );
  NAND2X1 U383 ( .A(\mem<22><7> ), .B(n1793), .Y(n2731) );
  OAI21X1 U384 ( .A(n1832), .B(n1791), .C(n2730), .Y(n2215) );
  NAND2X1 U385 ( .A(\mem<22><8> ), .B(n1792), .Y(n2730) );
  OAI21X1 U386 ( .A(n1831), .B(n1791), .C(n2729), .Y(n2214) );
  NAND2X1 U387 ( .A(\mem<22><9> ), .B(n1792), .Y(n2729) );
  OAI21X1 U388 ( .A(n1830), .B(n1791), .C(n2728), .Y(n2213) );
  NAND2X1 U389 ( .A(\mem<22><10> ), .B(n1792), .Y(n2728) );
  OAI21X1 U390 ( .A(n1829), .B(n1791), .C(n2727), .Y(n2212) );
  NAND2X1 U391 ( .A(\mem<22><11> ), .B(n1792), .Y(n2727) );
  OAI21X1 U392 ( .A(n1828), .B(n1791), .C(n2726), .Y(n2211) );
  NAND2X1 U393 ( .A(\mem<22><12> ), .B(n1792), .Y(n2726) );
  OAI21X1 U394 ( .A(n1827), .B(n1791), .C(n2725), .Y(n2210) );
  NAND2X1 U395 ( .A(\mem<22><13> ), .B(n1792), .Y(n2725) );
  OAI21X1 U396 ( .A(n1826), .B(n1791), .C(n2724), .Y(n2209) );
  NAND2X1 U397 ( .A(\mem<22><14> ), .B(n1792), .Y(n2724) );
  OAI21X1 U398 ( .A(n1825), .B(n1791), .C(n2723), .Y(n2208) );
  NAND2X1 U399 ( .A(\mem<22><15> ), .B(n1792), .Y(n2723) );
  OAI21X1 U402 ( .A(n1840), .B(n1788), .C(n2722), .Y(n2207) );
  NAND2X1 U403 ( .A(\mem<21><0> ), .B(n1790), .Y(n2722) );
  OAI21X1 U404 ( .A(n1839), .B(n1788), .C(n2721), .Y(n2206) );
  NAND2X1 U405 ( .A(\mem<21><1> ), .B(n1790), .Y(n2721) );
  OAI21X1 U406 ( .A(n1838), .B(n1788), .C(n2720), .Y(n2205) );
  NAND2X1 U407 ( .A(\mem<21><2> ), .B(n1790), .Y(n2720) );
  OAI21X1 U408 ( .A(n1837), .B(n1788), .C(n2719), .Y(n2204) );
  NAND2X1 U409 ( .A(\mem<21><3> ), .B(n1790), .Y(n2719) );
  OAI21X1 U410 ( .A(n1836), .B(n1788), .C(n2718), .Y(n2203) );
  NAND2X1 U411 ( .A(\mem<21><4> ), .B(n1790), .Y(n2718) );
  OAI21X1 U412 ( .A(n1835), .B(n1788), .C(n2717), .Y(n2202) );
  NAND2X1 U413 ( .A(\mem<21><5> ), .B(n1790), .Y(n2717) );
  OAI21X1 U414 ( .A(n1834), .B(n1788), .C(n2716), .Y(n2201) );
  NAND2X1 U415 ( .A(\mem<21><6> ), .B(n1790), .Y(n2716) );
  OAI21X1 U416 ( .A(n1833), .B(n1788), .C(n2715), .Y(n2200) );
  NAND2X1 U417 ( .A(\mem<21><7> ), .B(n1790), .Y(n2715) );
  OAI21X1 U418 ( .A(n1832), .B(n1788), .C(n2714), .Y(n2199) );
  NAND2X1 U419 ( .A(\mem<21><8> ), .B(n1789), .Y(n2714) );
  OAI21X1 U420 ( .A(n1831), .B(n1788), .C(n2713), .Y(n2198) );
  NAND2X1 U421 ( .A(\mem<21><9> ), .B(n1789), .Y(n2713) );
  OAI21X1 U422 ( .A(n1830), .B(n1788), .C(n2712), .Y(n2197) );
  NAND2X1 U423 ( .A(\mem<21><10> ), .B(n1789), .Y(n2712) );
  OAI21X1 U424 ( .A(n1829), .B(n1788), .C(n2711), .Y(n2196) );
  NAND2X1 U425 ( .A(\mem<21><11> ), .B(n1789), .Y(n2711) );
  OAI21X1 U426 ( .A(n1828), .B(n1788), .C(n2710), .Y(n2195) );
  NAND2X1 U427 ( .A(\mem<21><12> ), .B(n1789), .Y(n2710) );
  OAI21X1 U428 ( .A(n1827), .B(n1788), .C(n2709), .Y(n2194) );
  NAND2X1 U429 ( .A(\mem<21><13> ), .B(n1789), .Y(n2709) );
  OAI21X1 U430 ( .A(n1826), .B(n1788), .C(n2708), .Y(n2193) );
  NAND2X1 U431 ( .A(\mem<21><14> ), .B(n1789), .Y(n2708) );
  OAI21X1 U432 ( .A(n1825), .B(n1788), .C(n2707), .Y(n2192) );
  NAND2X1 U433 ( .A(\mem<21><15> ), .B(n1789), .Y(n2707) );
  OAI21X1 U436 ( .A(n1840), .B(n1785), .C(n2706), .Y(n2191) );
  NAND2X1 U437 ( .A(\mem<20><0> ), .B(n1787), .Y(n2706) );
  OAI21X1 U438 ( .A(n1839), .B(n1785), .C(n2705), .Y(n2190) );
  NAND2X1 U439 ( .A(\mem<20><1> ), .B(n1787), .Y(n2705) );
  OAI21X1 U440 ( .A(n1838), .B(n1785), .C(n2704), .Y(n2189) );
  NAND2X1 U441 ( .A(\mem<20><2> ), .B(n1787), .Y(n2704) );
  OAI21X1 U442 ( .A(n1837), .B(n1785), .C(n2703), .Y(n2188) );
  NAND2X1 U443 ( .A(\mem<20><3> ), .B(n1787), .Y(n2703) );
  OAI21X1 U444 ( .A(n1836), .B(n1785), .C(n2702), .Y(n2187) );
  NAND2X1 U445 ( .A(\mem<20><4> ), .B(n1787), .Y(n2702) );
  OAI21X1 U446 ( .A(n1835), .B(n1785), .C(n2701), .Y(n2186) );
  NAND2X1 U447 ( .A(\mem<20><5> ), .B(n1787), .Y(n2701) );
  OAI21X1 U448 ( .A(n1834), .B(n1785), .C(n2700), .Y(n2185) );
  NAND2X1 U449 ( .A(\mem<20><6> ), .B(n1787), .Y(n2700) );
  OAI21X1 U450 ( .A(n1833), .B(n1785), .C(n2699), .Y(n2184) );
  NAND2X1 U451 ( .A(\mem<20><7> ), .B(n1787), .Y(n2699) );
  OAI21X1 U452 ( .A(n1832), .B(n1785), .C(n2698), .Y(n2183) );
  NAND2X1 U453 ( .A(\mem<20><8> ), .B(n1786), .Y(n2698) );
  OAI21X1 U454 ( .A(n1831), .B(n1785), .C(n2697), .Y(n2182) );
  NAND2X1 U455 ( .A(\mem<20><9> ), .B(n1786), .Y(n2697) );
  OAI21X1 U456 ( .A(n1830), .B(n1785), .C(n2696), .Y(n2181) );
  NAND2X1 U457 ( .A(\mem<20><10> ), .B(n1786), .Y(n2696) );
  OAI21X1 U458 ( .A(n1829), .B(n1785), .C(n2695), .Y(n2180) );
  NAND2X1 U459 ( .A(\mem<20><11> ), .B(n1786), .Y(n2695) );
  OAI21X1 U460 ( .A(n1828), .B(n1785), .C(n2694), .Y(n2179) );
  NAND2X1 U461 ( .A(\mem<20><12> ), .B(n1786), .Y(n2694) );
  OAI21X1 U462 ( .A(n1827), .B(n1785), .C(n2693), .Y(n2178) );
  NAND2X1 U463 ( .A(\mem<20><13> ), .B(n1786), .Y(n2693) );
  OAI21X1 U464 ( .A(n1826), .B(n1785), .C(n2692), .Y(n2177) );
  NAND2X1 U465 ( .A(\mem<20><14> ), .B(n1786), .Y(n2692) );
  OAI21X1 U466 ( .A(n1825), .B(n1785), .C(n2691), .Y(n2176) );
  NAND2X1 U467 ( .A(\mem<20><15> ), .B(n1786), .Y(n2691) );
  OAI21X1 U470 ( .A(n1840), .B(n1782), .C(n2690), .Y(n2175) );
  NAND2X1 U471 ( .A(\mem<19><0> ), .B(n1784), .Y(n2690) );
  OAI21X1 U472 ( .A(n1839), .B(n1782), .C(n2689), .Y(n2174) );
  NAND2X1 U473 ( .A(\mem<19><1> ), .B(n1784), .Y(n2689) );
  OAI21X1 U474 ( .A(n1838), .B(n1782), .C(n2688), .Y(n2173) );
  NAND2X1 U475 ( .A(\mem<19><2> ), .B(n1784), .Y(n2688) );
  OAI21X1 U476 ( .A(n1837), .B(n1782), .C(n2687), .Y(n2172) );
  NAND2X1 U477 ( .A(\mem<19><3> ), .B(n1784), .Y(n2687) );
  OAI21X1 U478 ( .A(n1836), .B(n1782), .C(n2686), .Y(n2171) );
  NAND2X1 U479 ( .A(\mem<19><4> ), .B(n1784), .Y(n2686) );
  OAI21X1 U480 ( .A(n1835), .B(n1782), .C(n2685), .Y(n2170) );
  NAND2X1 U481 ( .A(\mem<19><5> ), .B(n1784), .Y(n2685) );
  OAI21X1 U482 ( .A(n1834), .B(n1782), .C(n2684), .Y(n2169) );
  NAND2X1 U483 ( .A(\mem<19><6> ), .B(n1784), .Y(n2684) );
  OAI21X1 U484 ( .A(n1833), .B(n1782), .C(n2683), .Y(n2168) );
  NAND2X1 U485 ( .A(\mem<19><7> ), .B(n1784), .Y(n2683) );
  OAI21X1 U486 ( .A(n1832), .B(n1782), .C(n2682), .Y(n2167) );
  NAND2X1 U487 ( .A(\mem<19><8> ), .B(n1783), .Y(n2682) );
  OAI21X1 U488 ( .A(n1831), .B(n1782), .C(n2681), .Y(n2166) );
  NAND2X1 U489 ( .A(\mem<19><9> ), .B(n1783), .Y(n2681) );
  OAI21X1 U490 ( .A(n1830), .B(n1782), .C(n2680), .Y(n2165) );
  NAND2X1 U491 ( .A(\mem<19><10> ), .B(n1783), .Y(n2680) );
  OAI21X1 U492 ( .A(n1829), .B(n1782), .C(n2679), .Y(n2164) );
  NAND2X1 U493 ( .A(\mem<19><11> ), .B(n1783), .Y(n2679) );
  OAI21X1 U494 ( .A(n1828), .B(n1782), .C(n2678), .Y(n2163) );
  NAND2X1 U495 ( .A(\mem<19><12> ), .B(n1783), .Y(n2678) );
  OAI21X1 U496 ( .A(n1827), .B(n1782), .C(n2677), .Y(n2162) );
  NAND2X1 U497 ( .A(\mem<19><13> ), .B(n1783), .Y(n2677) );
  OAI21X1 U498 ( .A(n1826), .B(n1782), .C(n2676), .Y(n2161) );
  NAND2X1 U499 ( .A(\mem<19><14> ), .B(n1783), .Y(n2676) );
  OAI21X1 U500 ( .A(n1825), .B(n1782), .C(n2675), .Y(n2160) );
  NAND2X1 U501 ( .A(\mem<19><15> ), .B(n1783), .Y(n2675) );
  OAI21X1 U504 ( .A(n1840), .B(n1779), .C(n2674), .Y(n2159) );
  NAND2X1 U505 ( .A(\mem<18><0> ), .B(n1781), .Y(n2674) );
  OAI21X1 U506 ( .A(n1839), .B(n1779), .C(n2673), .Y(n2158) );
  NAND2X1 U507 ( .A(\mem<18><1> ), .B(n1781), .Y(n2673) );
  OAI21X1 U508 ( .A(n1838), .B(n1779), .C(n2672), .Y(n2157) );
  NAND2X1 U509 ( .A(\mem<18><2> ), .B(n1781), .Y(n2672) );
  OAI21X1 U510 ( .A(n1837), .B(n1779), .C(n2671), .Y(n2156) );
  NAND2X1 U511 ( .A(\mem<18><3> ), .B(n1781), .Y(n2671) );
  OAI21X1 U512 ( .A(n1836), .B(n1779), .C(n2670), .Y(n2155) );
  NAND2X1 U513 ( .A(\mem<18><4> ), .B(n1781), .Y(n2670) );
  OAI21X1 U514 ( .A(n1835), .B(n1779), .C(n2669), .Y(n2154) );
  NAND2X1 U515 ( .A(\mem<18><5> ), .B(n1781), .Y(n2669) );
  OAI21X1 U516 ( .A(n1834), .B(n1779), .C(n2668), .Y(n2153) );
  NAND2X1 U517 ( .A(\mem<18><6> ), .B(n1781), .Y(n2668) );
  OAI21X1 U518 ( .A(n1833), .B(n1779), .C(n2667), .Y(n2152) );
  NAND2X1 U519 ( .A(\mem<18><7> ), .B(n1781), .Y(n2667) );
  OAI21X1 U520 ( .A(n1832), .B(n1779), .C(n2666), .Y(n2151) );
  NAND2X1 U521 ( .A(\mem<18><8> ), .B(n1780), .Y(n2666) );
  OAI21X1 U522 ( .A(n1831), .B(n1779), .C(n2665), .Y(n2150) );
  NAND2X1 U523 ( .A(\mem<18><9> ), .B(n1780), .Y(n2665) );
  OAI21X1 U524 ( .A(n1830), .B(n1779), .C(n2664), .Y(n2149) );
  NAND2X1 U525 ( .A(\mem<18><10> ), .B(n1780), .Y(n2664) );
  OAI21X1 U526 ( .A(n1829), .B(n1779), .C(n2663), .Y(n2148) );
  NAND2X1 U527 ( .A(\mem<18><11> ), .B(n1780), .Y(n2663) );
  OAI21X1 U528 ( .A(n1828), .B(n1779), .C(n2662), .Y(n2147) );
  NAND2X1 U529 ( .A(\mem<18><12> ), .B(n1780), .Y(n2662) );
  OAI21X1 U530 ( .A(n1827), .B(n1779), .C(n2661), .Y(n2146) );
  NAND2X1 U531 ( .A(\mem<18><13> ), .B(n1780), .Y(n2661) );
  OAI21X1 U532 ( .A(n1826), .B(n1779), .C(n2660), .Y(n2145) );
  NAND2X1 U533 ( .A(\mem<18><14> ), .B(n1780), .Y(n2660) );
  OAI21X1 U534 ( .A(n1825), .B(n1779), .C(n2659), .Y(n2144) );
  NAND2X1 U535 ( .A(\mem<18><15> ), .B(n1780), .Y(n2659) );
  OAI21X1 U538 ( .A(n1840), .B(n1776), .C(n2658), .Y(n2143) );
  NAND2X1 U539 ( .A(\mem<17><0> ), .B(n1778), .Y(n2658) );
  OAI21X1 U540 ( .A(n1839), .B(n1776), .C(n2657), .Y(n2142) );
  NAND2X1 U541 ( .A(\mem<17><1> ), .B(n1778), .Y(n2657) );
  OAI21X1 U542 ( .A(n1838), .B(n1776), .C(n2656), .Y(n2141) );
  NAND2X1 U543 ( .A(\mem<17><2> ), .B(n1778), .Y(n2656) );
  OAI21X1 U544 ( .A(n1837), .B(n1776), .C(n2655), .Y(n2140) );
  NAND2X1 U545 ( .A(\mem<17><3> ), .B(n1778), .Y(n2655) );
  OAI21X1 U546 ( .A(n1836), .B(n1776), .C(n2654), .Y(n2139) );
  NAND2X1 U547 ( .A(\mem<17><4> ), .B(n1778), .Y(n2654) );
  OAI21X1 U548 ( .A(n1835), .B(n1776), .C(n2653), .Y(n2138) );
  NAND2X1 U549 ( .A(\mem<17><5> ), .B(n1778), .Y(n2653) );
  OAI21X1 U550 ( .A(n1834), .B(n1776), .C(n2652), .Y(n2137) );
  NAND2X1 U551 ( .A(\mem<17><6> ), .B(n1778), .Y(n2652) );
  OAI21X1 U552 ( .A(n1833), .B(n1776), .C(n2651), .Y(n2136) );
  NAND2X1 U553 ( .A(\mem<17><7> ), .B(n1778), .Y(n2651) );
  OAI21X1 U554 ( .A(n1832), .B(n1776), .C(n2650), .Y(n2135) );
  NAND2X1 U555 ( .A(\mem<17><8> ), .B(n1777), .Y(n2650) );
  OAI21X1 U556 ( .A(n1831), .B(n1776), .C(n2649), .Y(n2134) );
  NAND2X1 U557 ( .A(\mem<17><9> ), .B(n1777), .Y(n2649) );
  OAI21X1 U558 ( .A(n1830), .B(n1776), .C(n2648), .Y(n2133) );
  NAND2X1 U559 ( .A(\mem<17><10> ), .B(n1777), .Y(n2648) );
  OAI21X1 U560 ( .A(n1829), .B(n1776), .C(n2647), .Y(n2132) );
  NAND2X1 U561 ( .A(\mem<17><11> ), .B(n1777), .Y(n2647) );
  OAI21X1 U562 ( .A(n1828), .B(n1776), .C(n2646), .Y(n2131) );
  NAND2X1 U563 ( .A(\mem<17><12> ), .B(n1777), .Y(n2646) );
  OAI21X1 U564 ( .A(n1827), .B(n1776), .C(n2645), .Y(n2130) );
  NAND2X1 U565 ( .A(\mem<17><13> ), .B(n1777), .Y(n2645) );
  OAI21X1 U566 ( .A(n1826), .B(n1776), .C(n2644), .Y(n2129) );
  NAND2X1 U567 ( .A(\mem<17><14> ), .B(n1777), .Y(n2644) );
  OAI21X1 U568 ( .A(n1825), .B(n1776), .C(n2643), .Y(n2128) );
  NAND2X1 U569 ( .A(\mem<17><15> ), .B(n1777), .Y(n2643) );
  OAI21X1 U572 ( .A(n1840), .B(n1773), .C(n2642), .Y(n2127) );
  NAND2X1 U573 ( .A(\mem<16><0> ), .B(n1775), .Y(n2642) );
  OAI21X1 U574 ( .A(n1839), .B(n1773), .C(n2641), .Y(n2126) );
  NAND2X1 U575 ( .A(\mem<16><1> ), .B(n1775), .Y(n2641) );
  OAI21X1 U576 ( .A(n1838), .B(n1773), .C(n2640), .Y(n2125) );
  NAND2X1 U577 ( .A(\mem<16><2> ), .B(n1775), .Y(n2640) );
  OAI21X1 U578 ( .A(n1837), .B(n1773), .C(n2639), .Y(n2124) );
  NAND2X1 U579 ( .A(\mem<16><3> ), .B(n1775), .Y(n2639) );
  OAI21X1 U580 ( .A(n1836), .B(n1773), .C(n2638), .Y(n2123) );
  NAND2X1 U581 ( .A(\mem<16><4> ), .B(n1775), .Y(n2638) );
  OAI21X1 U582 ( .A(n1835), .B(n1773), .C(n2637), .Y(n2122) );
  NAND2X1 U583 ( .A(\mem<16><5> ), .B(n1775), .Y(n2637) );
  OAI21X1 U584 ( .A(n1834), .B(n1773), .C(n2636), .Y(n2121) );
  NAND2X1 U585 ( .A(\mem<16><6> ), .B(n1775), .Y(n2636) );
  OAI21X1 U586 ( .A(n1833), .B(n1773), .C(n2635), .Y(n2120) );
  NAND2X1 U587 ( .A(\mem<16><7> ), .B(n1775), .Y(n2635) );
  OAI21X1 U588 ( .A(n1832), .B(n1773), .C(n2634), .Y(n2119) );
  NAND2X1 U589 ( .A(\mem<16><8> ), .B(n1774), .Y(n2634) );
  OAI21X1 U590 ( .A(n1831), .B(n1773), .C(n2633), .Y(n2118) );
  NAND2X1 U591 ( .A(\mem<16><9> ), .B(n1774), .Y(n2633) );
  OAI21X1 U592 ( .A(n1830), .B(n1773), .C(n2632), .Y(n2117) );
  NAND2X1 U593 ( .A(\mem<16><10> ), .B(n1774), .Y(n2632) );
  OAI21X1 U594 ( .A(n1829), .B(n1773), .C(n2631), .Y(n2116) );
  NAND2X1 U595 ( .A(\mem<16><11> ), .B(n1774), .Y(n2631) );
  OAI21X1 U596 ( .A(n1828), .B(n1773), .C(n2630), .Y(n2115) );
  NAND2X1 U597 ( .A(\mem<16><12> ), .B(n1774), .Y(n2630) );
  OAI21X1 U598 ( .A(n1827), .B(n1773), .C(n2629), .Y(n2114) );
  NAND2X1 U599 ( .A(\mem<16><13> ), .B(n1774), .Y(n2629) );
  OAI21X1 U600 ( .A(n1826), .B(n1773), .C(n2628), .Y(n2113) );
  NAND2X1 U601 ( .A(\mem<16><14> ), .B(n1774), .Y(n2628) );
  OAI21X1 U602 ( .A(n1825), .B(n1773), .C(n2627), .Y(n2112) );
  NAND2X1 U603 ( .A(\mem<16><15> ), .B(n1774), .Y(n2627) );
  NAND3X1 U606 ( .A(n2755), .B(n1847), .C(n1848), .Y(n2626) );
  OAI21X1 U607 ( .A(n1840), .B(n1770), .C(n2625), .Y(n2111) );
  NAND2X1 U608 ( .A(\mem<15><0> ), .B(n1772), .Y(n2625) );
  OAI21X1 U609 ( .A(n1839), .B(n1770), .C(n2624), .Y(n2110) );
  NAND2X1 U610 ( .A(\mem<15><1> ), .B(n1772), .Y(n2624) );
  OAI21X1 U611 ( .A(n1838), .B(n1770), .C(n2623), .Y(n2109) );
  NAND2X1 U612 ( .A(\mem<15><2> ), .B(n1772), .Y(n2623) );
  OAI21X1 U613 ( .A(n1837), .B(n1770), .C(n2622), .Y(n2108) );
  NAND2X1 U614 ( .A(\mem<15><3> ), .B(n1772), .Y(n2622) );
  OAI21X1 U615 ( .A(n1836), .B(n1770), .C(n2621), .Y(n2107) );
  NAND2X1 U616 ( .A(\mem<15><4> ), .B(n1772), .Y(n2621) );
  OAI21X1 U617 ( .A(n1835), .B(n1770), .C(n2620), .Y(n2106) );
  NAND2X1 U618 ( .A(\mem<15><5> ), .B(n1772), .Y(n2620) );
  OAI21X1 U619 ( .A(n1834), .B(n1770), .C(n2619), .Y(n2105) );
  NAND2X1 U620 ( .A(\mem<15><6> ), .B(n1772), .Y(n2619) );
  OAI21X1 U621 ( .A(n1833), .B(n1770), .C(n2618), .Y(n2104) );
  NAND2X1 U622 ( .A(\mem<15><7> ), .B(n1772), .Y(n2618) );
  OAI21X1 U623 ( .A(n1832), .B(n1770), .C(n2617), .Y(n2103) );
  NAND2X1 U624 ( .A(\mem<15><8> ), .B(n1771), .Y(n2617) );
  OAI21X1 U625 ( .A(n1831), .B(n1770), .C(n2616), .Y(n2102) );
  NAND2X1 U626 ( .A(\mem<15><9> ), .B(n1771), .Y(n2616) );
  OAI21X1 U627 ( .A(n1830), .B(n1770), .C(n2615), .Y(n2101) );
  NAND2X1 U628 ( .A(\mem<15><10> ), .B(n1771), .Y(n2615) );
  OAI21X1 U629 ( .A(n1829), .B(n1770), .C(n2614), .Y(n2100) );
  NAND2X1 U630 ( .A(\mem<15><11> ), .B(n1771), .Y(n2614) );
  OAI21X1 U631 ( .A(n1828), .B(n1770), .C(n2613), .Y(n2099) );
  NAND2X1 U632 ( .A(\mem<15><12> ), .B(n1771), .Y(n2613) );
  OAI21X1 U633 ( .A(n1827), .B(n1770), .C(n2612), .Y(n2098) );
  NAND2X1 U634 ( .A(\mem<15><13> ), .B(n1771), .Y(n2612) );
  OAI21X1 U635 ( .A(n1826), .B(n1770), .C(n2611), .Y(n2097) );
  NAND2X1 U636 ( .A(\mem<15><14> ), .B(n1771), .Y(n2611) );
  OAI21X1 U637 ( .A(n1825), .B(n1770), .C(n2610), .Y(n2096) );
  NAND2X1 U638 ( .A(\mem<15><15> ), .B(n1771), .Y(n2610) );
  OAI21X1 U641 ( .A(n1840), .B(n1767), .C(n2609), .Y(n2095) );
  NAND2X1 U642 ( .A(\mem<14><0> ), .B(n1769), .Y(n2609) );
  OAI21X1 U643 ( .A(n1839), .B(n1767), .C(n2608), .Y(n2094) );
  NAND2X1 U644 ( .A(\mem<14><1> ), .B(n1769), .Y(n2608) );
  OAI21X1 U645 ( .A(n1838), .B(n1767), .C(n2607), .Y(n2093) );
  NAND2X1 U646 ( .A(\mem<14><2> ), .B(n1769), .Y(n2607) );
  OAI21X1 U647 ( .A(n1837), .B(n1767), .C(n2606), .Y(n2092) );
  NAND2X1 U648 ( .A(\mem<14><3> ), .B(n1769), .Y(n2606) );
  OAI21X1 U649 ( .A(n1836), .B(n1767), .C(n2605), .Y(n2091) );
  NAND2X1 U650 ( .A(\mem<14><4> ), .B(n1769), .Y(n2605) );
  OAI21X1 U651 ( .A(n1835), .B(n1767), .C(n2604), .Y(n2090) );
  NAND2X1 U652 ( .A(\mem<14><5> ), .B(n1769), .Y(n2604) );
  OAI21X1 U653 ( .A(n1834), .B(n1767), .C(n2603), .Y(n2089) );
  NAND2X1 U654 ( .A(\mem<14><6> ), .B(n1769), .Y(n2603) );
  OAI21X1 U655 ( .A(n1833), .B(n1767), .C(n2602), .Y(n2088) );
  NAND2X1 U656 ( .A(\mem<14><7> ), .B(n1769), .Y(n2602) );
  OAI21X1 U657 ( .A(n1832), .B(n1767), .C(n2601), .Y(n2087) );
  NAND2X1 U658 ( .A(\mem<14><8> ), .B(n1768), .Y(n2601) );
  OAI21X1 U659 ( .A(n1831), .B(n1767), .C(n2600), .Y(n2086) );
  NAND2X1 U660 ( .A(\mem<14><9> ), .B(n1768), .Y(n2600) );
  OAI21X1 U661 ( .A(n1830), .B(n1767), .C(n2599), .Y(n2085) );
  NAND2X1 U662 ( .A(\mem<14><10> ), .B(n1768), .Y(n2599) );
  OAI21X1 U663 ( .A(n1829), .B(n1767), .C(n2598), .Y(n2084) );
  NAND2X1 U664 ( .A(\mem<14><11> ), .B(n1768), .Y(n2598) );
  OAI21X1 U665 ( .A(n1828), .B(n1767), .C(n2597), .Y(n2083) );
  NAND2X1 U666 ( .A(\mem<14><12> ), .B(n1768), .Y(n2597) );
  OAI21X1 U667 ( .A(n1827), .B(n1767), .C(n2596), .Y(n2082) );
  NAND2X1 U668 ( .A(\mem<14><13> ), .B(n1768), .Y(n2596) );
  OAI21X1 U669 ( .A(n1826), .B(n1767), .C(n2595), .Y(n2081) );
  NAND2X1 U670 ( .A(\mem<14><14> ), .B(n1768), .Y(n2595) );
  OAI21X1 U671 ( .A(n1825), .B(n1767), .C(n2594), .Y(n2080) );
  NAND2X1 U672 ( .A(\mem<14><15> ), .B(n1768), .Y(n2594) );
  OAI21X1 U675 ( .A(n1840), .B(n1764), .C(n2593), .Y(n2079) );
  NAND2X1 U676 ( .A(\mem<13><0> ), .B(n1766), .Y(n2593) );
  OAI21X1 U677 ( .A(n1839), .B(n1764), .C(n2592), .Y(n2078) );
  NAND2X1 U678 ( .A(\mem<13><1> ), .B(n1766), .Y(n2592) );
  OAI21X1 U679 ( .A(n1838), .B(n1764), .C(n2591), .Y(n2077) );
  NAND2X1 U680 ( .A(\mem<13><2> ), .B(n1766), .Y(n2591) );
  OAI21X1 U681 ( .A(n1837), .B(n1764), .C(n2590), .Y(n2076) );
  NAND2X1 U682 ( .A(\mem<13><3> ), .B(n1766), .Y(n2590) );
  OAI21X1 U683 ( .A(n1836), .B(n1764), .C(n2589), .Y(n2075) );
  NAND2X1 U684 ( .A(\mem<13><4> ), .B(n1766), .Y(n2589) );
  OAI21X1 U685 ( .A(n1835), .B(n1764), .C(n2588), .Y(n2074) );
  NAND2X1 U686 ( .A(\mem<13><5> ), .B(n1766), .Y(n2588) );
  OAI21X1 U687 ( .A(n1834), .B(n1764), .C(n2587), .Y(n2073) );
  NAND2X1 U688 ( .A(\mem<13><6> ), .B(n1766), .Y(n2587) );
  OAI21X1 U689 ( .A(n1833), .B(n1764), .C(n2586), .Y(n2072) );
  NAND2X1 U690 ( .A(\mem<13><7> ), .B(n1766), .Y(n2586) );
  OAI21X1 U691 ( .A(n1832), .B(n1764), .C(n2585), .Y(n2071) );
  NAND2X1 U692 ( .A(\mem<13><8> ), .B(n1765), .Y(n2585) );
  OAI21X1 U693 ( .A(n1831), .B(n1764), .C(n2584), .Y(n2070) );
  NAND2X1 U694 ( .A(\mem<13><9> ), .B(n1765), .Y(n2584) );
  OAI21X1 U695 ( .A(n1830), .B(n1764), .C(n2583), .Y(n2069) );
  NAND2X1 U696 ( .A(\mem<13><10> ), .B(n1765), .Y(n2583) );
  OAI21X1 U697 ( .A(n1829), .B(n1764), .C(n2582), .Y(n2068) );
  NAND2X1 U698 ( .A(\mem<13><11> ), .B(n1765), .Y(n2582) );
  OAI21X1 U699 ( .A(n1828), .B(n1764), .C(n2581), .Y(n2067) );
  NAND2X1 U700 ( .A(\mem<13><12> ), .B(n1765), .Y(n2581) );
  OAI21X1 U701 ( .A(n1827), .B(n1764), .C(n2580), .Y(n2066) );
  NAND2X1 U702 ( .A(\mem<13><13> ), .B(n1765), .Y(n2580) );
  OAI21X1 U703 ( .A(n1826), .B(n1764), .C(n2579), .Y(n2065) );
  NAND2X1 U704 ( .A(\mem<13><14> ), .B(n1765), .Y(n2579) );
  OAI21X1 U705 ( .A(n1825), .B(n1764), .C(n2578), .Y(n2064) );
  NAND2X1 U706 ( .A(\mem<13><15> ), .B(n1765), .Y(n2578) );
  OAI21X1 U709 ( .A(n1840), .B(n1761), .C(n2577), .Y(n2063) );
  NAND2X1 U710 ( .A(\mem<12><0> ), .B(n1763), .Y(n2577) );
  OAI21X1 U711 ( .A(n1839), .B(n1761), .C(n2576), .Y(n2062) );
  NAND2X1 U712 ( .A(\mem<12><1> ), .B(n1763), .Y(n2576) );
  OAI21X1 U713 ( .A(n1838), .B(n1761), .C(n2575), .Y(n2061) );
  NAND2X1 U714 ( .A(\mem<12><2> ), .B(n1763), .Y(n2575) );
  OAI21X1 U715 ( .A(n1837), .B(n1761), .C(n2574), .Y(n2060) );
  NAND2X1 U716 ( .A(\mem<12><3> ), .B(n1763), .Y(n2574) );
  OAI21X1 U717 ( .A(n1836), .B(n1761), .C(n2573), .Y(n2059) );
  NAND2X1 U718 ( .A(\mem<12><4> ), .B(n1763), .Y(n2573) );
  OAI21X1 U719 ( .A(n1835), .B(n1761), .C(n2572), .Y(n2058) );
  NAND2X1 U720 ( .A(\mem<12><5> ), .B(n1763), .Y(n2572) );
  OAI21X1 U721 ( .A(n1834), .B(n1761), .C(n2571), .Y(n2057) );
  NAND2X1 U722 ( .A(\mem<12><6> ), .B(n1763), .Y(n2571) );
  OAI21X1 U723 ( .A(n1833), .B(n1761), .C(n2570), .Y(n2056) );
  NAND2X1 U724 ( .A(\mem<12><7> ), .B(n1763), .Y(n2570) );
  OAI21X1 U725 ( .A(n1832), .B(n1761), .C(n2569), .Y(n2055) );
  NAND2X1 U726 ( .A(\mem<12><8> ), .B(n1762), .Y(n2569) );
  OAI21X1 U727 ( .A(n1831), .B(n1761), .C(n2568), .Y(n2054) );
  NAND2X1 U728 ( .A(\mem<12><9> ), .B(n1762), .Y(n2568) );
  OAI21X1 U729 ( .A(n1830), .B(n1761), .C(n2567), .Y(n2053) );
  NAND2X1 U730 ( .A(\mem<12><10> ), .B(n1762), .Y(n2567) );
  OAI21X1 U731 ( .A(n1829), .B(n1761), .C(n2566), .Y(n2052) );
  NAND2X1 U732 ( .A(\mem<12><11> ), .B(n1762), .Y(n2566) );
  OAI21X1 U733 ( .A(n1828), .B(n1761), .C(n2565), .Y(n2051) );
  NAND2X1 U734 ( .A(\mem<12><12> ), .B(n1762), .Y(n2565) );
  OAI21X1 U735 ( .A(n1827), .B(n1761), .C(n2564), .Y(n2050) );
  NAND2X1 U736 ( .A(\mem<12><13> ), .B(n1762), .Y(n2564) );
  OAI21X1 U737 ( .A(n1826), .B(n1761), .C(n2563), .Y(n2049) );
  NAND2X1 U738 ( .A(\mem<12><14> ), .B(n1762), .Y(n2563) );
  OAI21X1 U739 ( .A(n1825), .B(n1761), .C(n2562), .Y(n2048) );
  NAND2X1 U740 ( .A(\mem<12><15> ), .B(n1762), .Y(n2562) );
  OAI21X1 U743 ( .A(n1840), .B(n1758), .C(n2561), .Y(n2047) );
  NAND2X1 U744 ( .A(\mem<11><0> ), .B(n1760), .Y(n2561) );
  OAI21X1 U745 ( .A(n1839), .B(n1758), .C(n2560), .Y(n2046) );
  NAND2X1 U746 ( .A(\mem<11><1> ), .B(n1760), .Y(n2560) );
  OAI21X1 U747 ( .A(n1838), .B(n1758), .C(n2559), .Y(n2045) );
  NAND2X1 U748 ( .A(\mem<11><2> ), .B(n1760), .Y(n2559) );
  OAI21X1 U749 ( .A(n1837), .B(n1758), .C(n2558), .Y(n2044) );
  NAND2X1 U750 ( .A(\mem<11><3> ), .B(n1760), .Y(n2558) );
  OAI21X1 U751 ( .A(n1836), .B(n1758), .C(n2557), .Y(n2043) );
  NAND2X1 U752 ( .A(\mem<11><4> ), .B(n1760), .Y(n2557) );
  OAI21X1 U753 ( .A(n1835), .B(n1758), .C(n2556), .Y(n2042) );
  NAND2X1 U754 ( .A(\mem<11><5> ), .B(n1760), .Y(n2556) );
  OAI21X1 U755 ( .A(n1834), .B(n1758), .C(n2555), .Y(n2041) );
  NAND2X1 U756 ( .A(\mem<11><6> ), .B(n1760), .Y(n2555) );
  OAI21X1 U757 ( .A(n1833), .B(n1758), .C(n2554), .Y(n2040) );
  NAND2X1 U758 ( .A(\mem<11><7> ), .B(n1760), .Y(n2554) );
  OAI21X1 U759 ( .A(n1832), .B(n1758), .C(n2553), .Y(n2039) );
  NAND2X1 U760 ( .A(\mem<11><8> ), .B(n1759), .Y(n2553) );
  OAI21X1 U761 ( .A(n1831), .B(n1758), .C(n2552), .Y(n2038) );
  NAND2X1 U762 ( .A(\mem<11><9> ), .B(n1759), .Y(n2552) );
  OAI21X1 U763 ( .A(n1830), .B(n1758), .C(n2551), .Y(n2037) );
  NAND2X1 U764 ( .A(\mem<11><10> ), .B(n1759), .Y(n2551) );
  OAI21X1 U765 ( .A(n1829), .B(n1758), .C(n2550), .Y(n2036) );
  NAND2X1 U766 ( .A(\mem<11><11> ), .B(n1759), .Y(n2550) );
  OAI21X1 U767 ( .A(n1828), .B(n1758), .C(n2549), .Y(n2035) );
  NAND2X1 U768 ( .A(\mem<11><12> ), .B(n1759), .Y(n2549) );
  OAI21X1 U769 ( .A(n1827), .B(n1758), .C(n2548), .Y(n2034) );
  NAND2X1 U770 ( .A(\mem<11><13> ), .B(n1759), .Y(n2548) );
  OAI21X1 U771 ( .A(n1826), .B(n1758), .C(n2547), .Y(n2033) );
  NAND2X1 U772 ( .A(\mem<11><14> ), .B(n1759), .Y(n2547) );
  OAI21X1 U773 ( .A(n1825), .B(n1758), .C(n2546), .Y(n2032) );
  NAND2X1 U774 ( .A(\mem<11><15> ), .B(n1759), .Y(n2546) );
  OAI21X1 U777 ( .A(n1840), .B(n1755), .C(n2545), .Y(n2031) );
  NAND2X1 U778 ( .A(\mem<10><0> ), .B(n1757), .Y(n2545) );
  OAI21X1 U779 ( .A(n1839), .B(n1755), .C(n2544), .Y(n2030) );
  NAND2X1 U780 ( .A(\mem<10><1> ), .B(n1757), .Y(n2544) );
  OAI21X1 U781 ( .A(n1838), .B(n1755), .C(n2543), .Y(n2029) );
  NAND2X1 U782 ( .A(\mem<10><2> ), .B(n1757), .Y(n2543) );
  OAI21X1 U783 ( .A(n1837), .B(n1755), .C(n2542), .Y(n2028) );
  NAND2X1 U784 ( .A(\mem<10><3> ), .B(n1757), .Y(n2542) );
  OAI21X1 U785 ( .A(n1836), .B(n1755), .C(n2541), .Y(n2027) );
  NAND2X1 U786 ( .A(\mem<10><4> ), .B(n1757), .Y(n2541) );
  OAI21X1 U787 ( .A(n1835), .B(n1755), .C(n2540), .Y(n2026) );
  NAND2X1 U788 ( .A(\mem<10><5> ), .B(n1757), .Y(n2540) );
  OAI21X1 U789 ( .A(n1834), .B(n1755), .C(n2539), .Y(n2025) );
  NAND2X1 U790 ( .A(\mem<10><6> ), .B(n1757), .Y(n2539) );
  OAI21X1 U791 ( .A(n1833), .B(n1755), .C(n2538), .Y(n2024) );
  NAND2X1 U792 ( .A(\mem<10><7> ), .B(n1757), .Y(n2538) );
  OAI21X1 U793 ( .A(n1832), .B(n1755), .C(n2537), .Y(n2023) );
  NAND2X1 U794 ( .A(\mem<10><8> ), .B(n1756), .Y(n2537) );
  OAI21X1 U795 ( .A(n1831), .B(n1755), .C(n2536), .Y(n2022) );
  NAND2X1 U796 ( .A(\mem<10><9> ), .B(n1756), .Y(n2536) );
  OAI21X1 U797 ( .A(n1830), .B(n1755), .C(n2535), .Y(n2021) );
  NAND2X1 U798 ( .A(\mem<10><10> ), .B(n1756), .Y(n2535) );
  OAI21X1 U799 ( .A(n1829), .B(n1755), .C(n2534), .Y(n2020) );
  NAND2X1 U800 ( .A(\mem<10><11> ), .B(n1756), .Y(n2534) );
  OAI21X1 U801 ( .A(n1828), .B(n1755), .C(n2533), .Y(n2019) );
  NAND2X1 U802 ( .A(\mem<10><12> ), .B(n1756), .Y(n2533) );
  OAI21X1 U803 ( .A(n1827), .B(n1755), .C(n2532), .Y(n2018) );
  NAND2X1 U804 ( .A(\mem<10><13> ), .B(n1756), .Y(n2532) );
  OAI21X1 U805 ( .A(n1826), .B(n1755), .C(n2531), .Y(n2017) );
  NAND2X1 U806 ( .A(\mem<10><14> ), .B(n1756), .Y(n2531) );
  OAI21X1 U807 ( .A(n1825), .B(n1755), .C(n2530), .Y(n2016) );
  NAND2X1 U808 ( .A(\mem<10><15> ), .B(n1756), .Y(n2530) );
  OAI21X1 U811 ( .A(n1840), .B(n1752), .C(n2529), .Y(n2015) );
  NAND2X1 U812 ( .A(\mem<9><0> ), .B(n1754), .Y(n2529) );
  OAI21X1 U813 ( .A(n1839), .B(n1752), .C(n2528), .Y(n2014) );
  NAND2X1 U814 ( .A(\mem<9><1> ), .B(n1754), .Y(n2528) );
  OAI21X1 U815 ( .A(n1838), .B(n1752), .C(n2527), .Y(n2013) );
  NAND2X1 U816 ( .A(\mem<9><2> ), .B(n1754), .Y(n2527) );
  OAI21X1 U817 ( .A(n1837), .B(n1752), .C(n2526), .Y(n2012) );
  NAND2X1 U818 ( .A(\mem<9><3> ), .B(n1754), .Y(n2526) );
  OAI21X1 U819 ( .A(n1836), .B(n1752), .C(n2525), .Y(n2011) );
  NAND2X1 U820 ( .A(\mem<9><4> ), .B(n1754), .Y(n2525) );
  OAI21X1 U821 ( .A(n1835), .B(n1752), .C(n2524), .Y(n2010) );
  NAND2X1 U822 ( .A(\mem<9><5> ), .B(n1754), .Y(n2524) );
  OAI21X1 U823 ( .A(n1834), .B(n1752), .C(n2523), .Y(n2009) );
  NAND2X1 U824 ( .A(\mem<9><6> ), .B(n1754), .Y(n2523) );
  OAI21X1 U825 ( .A(n1833), .B(n1752), .C(n2522), .Y(n2008) );
  NAND2X1 U826 ( .A(\mem<9><7> ), .B(n1754), .Y(n2522) );
  OAI21X1 U827 ( .A(n1832), .B(n1752), .C(n2521), .Y(n2007) );
  NAND2X1 U828 ( .A(\mem<9><8> ), .B(n1753), .Y(n2521) );
  OAI21X1 U829 ( .A(n1831), .B(n1752), .C(n2520), .Y(n2006) );
  NAND2X1 U830 ( .A(\mem<9><9> ), .B(n1753), .Y(n2520) );
  OAI21X1 U831 ( .A(n1830), .B(n1752), .C(n2519), .Y(n2005) );
  NAND2X1 U832 ( .A(\mem<9><10> ), .B(n1753), .Y(n2519) );
  OAI21X1 U833 ( .A(n1829), .B(n1752), .C(n2518), .Y(n2004) );
  NAND2X1 U834 ( .A(\mem<9><11> ), .B(n1753), .Y(n2518) );
  OAI21X1 U835 ( .A(n1828), .B(n1752), .C(n2517), .Y(n2003) );
  NAND2X1 U836 ( .A(\mem<9><12> ), .B(n1753), .Y(n2517) );
  OAI21X1 U837 ( .A(n1827), .B(n1752), .C(n2516), .Y(n2002) );
  NAND2X1 U838 ( .A(\mem<9><13> ), .B(n1753), .Y(n2516) );
  OAI21X1 U839 ( .A(n1826), .B(n1752), .C(n2515), .Y(n2001) );
  NAND2X1 U840 ( .A(\mem<9><14> ), .B(n1753), .Y(n2515) );
  OAI21X1 U841 ( .A(n1825), .B(n1752), .C(n2514), .Y(n2000) );
  NAND2X1 U842 ( .A(\mem<9><15> ), .B(n1753), .Y(n2514) );
  OAI21X1 U845 ( .A(n1840), .B(n1749), .C(n2513), .Y(n1999) );
  NAND2X1 U846 ( .A(\mem<8><0> ), .B(n1751), .Y(n2513) );
  OAI21X1 U847 ( .A(n1839), .B(n1749), .C(n2512), .Y(n1998) );
  NAND2X1 U848 ( .A(\mem<8><1> ), .B(n1751), .Y(n2512) );
  OAI21X1 U849 ( .A(n1838), .B(n1749), .C(n2511), .Y(n1997) );
  NAND2X1 U850 ( .A(\mem<8><2> ), .B(n1751), .Y(n2511) );
  OAI21X1 U851 ( .A(n1837), .B(n1749), .C(n2510), .Y(n1996) );
  NAND2X1 U852 ( .A(\mem<8><3> ), .B(n1751), .Y(n2510) );
  OAI21X1 U853 ( .A(n1836), .B(n1749), .C(n2509), .Y(n1995) );
  NAND2X1 U854 ( .A(\mem<8><4> ), .B(n1751), .Y(n2509) );
  OAI21X1 U855 ( .A(n1835), .B(n1749), .C(n2508), .Y(n1994) );
  NAND2X1 U856 ( .A(\mem<8><5> ), .B(n1751), .Y(n2508) );
  OAI21X1 U857 ( .A(n1834), .B(n1749), .C(n2507), .Y(n1993) );
  NAND2X1 U858 ( .A(\mem<8><6> ), .B(n1751), .Y(n2507) );
  OAI21X1 U859 ( .A(n1833), .B(n1749), .C(n2506), .Y(n1992) );
  NAND2X1 U860 ( .A(\mem<8><7> ), .B(n1751), .Y(n2506) );
  OAI21X1 U861 ( .A(n1832), .B(n1749), .C(n2505), .Y(n1991) );
  NAND2X1 U862 ( .A(\mem<8><8> ), .B(n1750), .Y(n2505) );
  OAI21X1 U863 ( .A(n1831), .B(n1749), .C(n2504), .Y(n1990) );
  NAND2X1 U864 ( .A(\mem<8><9> ), .B(n1750), .Y(n2504) );
  OAI21X1 U865 ( .A(n1830), .B(n1749), .C(n2503), .Y(n1989) );
  NAND2X1 U866 ( .A(\mem<8><10> ), .B(n1750), .Y(n2503) );
  OAI21X1 U867 ( .A(n1829), .B(n1749), .C(n2502), .Y(n1988) );
  NAND2X1 U868 ( .A(\mem<8><11> ), .B(n1750), .Y(n2502) );
  OAI21X1 U869 ( .A(n1828), .B(n1749), .C(n2501), .Y(n1987) );
  NAND2X1 U870 ( .A(\mem<8><12> ), .B(n1750), .Y(n2501) );
  OAI21X1 U871 ( .A(n1827), .B(n1749), .C(n2500), .Y(n1986) );
  NAND2X1 U872 ( .A(\mem<8><13> ), .B(n1750), .Y(n2500) );
  OAI21X1 U873 ( .A(n1826), .B(n1749), .C(n2499), .Y(n1985) );
  NAND2X1 U874 ( .A(\mem<8><14> ), .B(n1750), .Y(n2499) );
  OAI21X1 U875 ( .A(n1825), .B(n1749), .C(n2498), .Y(n1984) );
  NAND2X1 U876 ( .A(\mem<8><15> ), .B(n1750), .Y(n2498) );
  NAND3X1 U879 ( .A(n2755), .B(n1849), .C(n1846), .Y(n2497) );
  OAI21X1 U880 ( .A(n1840), .B(n1746), .C(n2496), .Y(n1983) );
  NAND2X1 U881 ( .A(\mem<7><0> ), .B(n1748), .Y(n2496) );
  OAI21X1 U882 ( .A(n1839), .B(n1746), .C(n2495), .Y(n1982) );
  NAND2X1 U883 ( .A(\mem<7><1> ), .B(n1748), .Y(n2495) );
  OAI21X1 U884 ( .A(n1838), .B(n1746), .C(n2494), .Y(n1981) );
  NAND2X1 U885 ( .A(\mem<7><2> ), .B(n1748), .Y(n2494) );
  OAI21X1 U886 ( .A(n1837), .B(n1746), .C(n2493), .Y(n1980) );
  NAND2X1 U887 ( .A(\mem<7><3> ), .B(n1748), .Y(n2493) );
  OAI21X1 U888 ( .A(n1836), .B(n1746), .C(n2492), .Y(n1979) );
  NAND2X1 U889 ( .A(\mem<7><4> ), .B(n1748), .Y(n2492) );
  OAI21X1 U890 ( .A(n1835), .B(n1746), .C(n2491), .Y(n1978) );
  NAND2X1 U891 ( .A(\mem<7><5> ), .B(n1748), .Y(n2491) );
  OAI21X1 U892 ( .A(n1834), .B(n1746), .C(n2490), .Y(n1977) );
  NAND2X1 U893 ( .A(\mem<7><6> ), .B(n1748), .Y(n2490) );
  OAI21X1 U894 ( .A(n1833), .B(n1746), .C(n2489), .Y(n1976) );
  NAND2X1 U895 ( .A(\mem<7><7> ), .B(n1748), .Y(n2489) );
  OAI21X1 U896 ( .A(n1832), .B(n1746), .C(n2488), .Y(n1975) );
  NAND2X1 U897 ( .A(\mem<7><8> ), .B(n1747), .Y(n2488) );
  OAI21X1 U898 ( .A(n1831), .B(n1746), .C(n2487), .Y(n1974) );
  NAND2X1 U899 ( .A(\mem<7><9> ), .B(n1747), .Y(n2487) );
  OAI21X1 U900 ( .A(n1830), .B(n1746), .C(n2486), .Y(n1973) );
  NAND2X1 U901 ( .A(\mem<7><10> ), .B(n1747), .Y(n2486) );
  OAI21X1 U902 ( .A(n1829), .B(n1746), .C(n2485), .Y(n1972) );
  NAND2X1 U903 ( .A(\mem<7><11> ), .B(n1747), .Y(n2485) );
  OAI21X1 U904 ( .A(n1828), .B(n1746), .C(n2484), .Y(n1971) );
  NAND2X1 U905 ( .A(\mem<7><12> ), .B(n1747), .Y(n2484) );
  OAI21X1 U906 ( .A(n1827), .B(n1746), .C(n2483), .Y(n1970) );
  NAND2X1 U907 ( .A(\mem<7><13> ), .B(n1747), .Y(n2483) );
  OAI21X1 U908 ( .A(n1826), .B(n1746), .C(n2482), .Y(n1969) );
  NAND2X1 U909 ( .A(\mem<7><14> ), .B(n1747), .Y(n2482) );
  OAI21X1 U910 ( .A(n1825), .B(n1746), .C(n2481), .Y(n1968) );
  NAND2X1 U911 ( .A(\mem<7><15> ), .B(n1747), .Y(n2481) );
  NOR3X1 U914 ( .A(n1844), .B(n1842), .C(n1845), .Y(n2876) );
  OAI21X1 U915 ( .A(n1840), .B(n1743), .C(n2480), .Y(n1967) );
  NAND2X1 U916 ( .A(\mem<6><0> ), .B(n1745), .Y(n2480) );
  OAI21X1 U917 ( .A(n1839), .B(n1743), .C(n2479), .Y(n1966) );
  NAND2X1 U918 ( .A(\mem<6><1> ), .B(n1745), .Y(n2479) );
  OAI21X1 U919 ( .A(n1838), .B(n1743), .C(n2478), .Y(n1965) );
  NAND2X1 U920 ( .A(\mem<6><2> ), .B(n1745), .Y(n2478) );
  OAI21X1 U921 ( .A(n1837), .B(n1743), .C(n2477), .Y(n1964) );
  NAND2X1 U922 ( .A(\mem<6><3> ), .B(n1745), .Y(n2477) );
  OAI21X1 U923 ( .A(n1836), .B(n1743), .C(n2476), .Y(n1963) );
  NAND2X1 U924 ( .A(\mem<6><4> ), .B(n1745), .Y(n2476) );
  OAI21X1 U925 ( .A(n1835), .B(n1743), .C(n2475), .Y(n1962) );
  NAND2X1 U926 ( .A(\mem<6><5> ), .B(n1745), .Y(n2475) );
  OAI21X1 U927 ( .A(n1834), .B(n1743), .C(n2474), .Y(n1961) );
  NAND2X1 U928 ( .A(\mem<6><6> ), .B(n1745), .Y(n2474) );
  OAI21X1 U929 ( .A(n1833), .B(n1743), .C(n2473), .Y(n1960) );
  NAND2X1 U930 ( .A(\mem<6><7> ), .B(n1745), .Y(n2473) );
  OAI21X1 U931 ( .A(n1832), .B(n1743), .C(n2472), .Y(n1959) );
  NAND2X1 U932 ( .A(\mem<6><8> ), .B(n1744), .Y(n2472) );
  OAI21X1 U933 ( .A(n1831), .B(n1743), .C(n2471), .Y(n1958) );
  NAND2X1 U934 ( .A(\mem<6><9> ), .B(n1744), .Y(n2471) );
  OAI21X1 U935 ( .A(n1830), .B(n1743), .C(n2470), .Y(n1957) );
  NAND2X1 U936 ( .A(\mem<6><10> ), .B(n1744), .Y(n2470) );
  OAI21X1 U937 ( .A(n1829), .B(n1743), .C(n2469), .Y(n1956) );
  NAND2X1 U938 ( .A(\mem<6><11> ), .B(n1744), .Y(n2469) );
  OAI21X1 U939 ( .A(n1828), .B(n1743), .C(n2468), .Y(n1955) );
  NAND2X1 U940 ( .A(\mem<6><12> ), .B(n1744), .Y(n2468) );
  OAI21X1 U941 ( .A(n1827), .B(n1743), .C(n2467), .Y(n1954) );
  NAND2X1 U942 ( .A(\mem<6><13> ), .B(n1744), .Y(n2467) );
  OAI21X1 U943 ( .A(n1826), .B(n1743), .C(n2466), .Y(n1953) );
  NAND2X1 U944 ( .A(\mem<6><14> ), .B(n1744), .Y(n2466) );
  OAI21X1 U945 ( .A(n1825), .B(n1743), .C(n2465), .Y(n1952) );
  NAND2X1 U946 ( .A(\mem<6><15> ), .B(n1744), .Y(n2465) );
  NOR3X1 U949 ( .A(n1844), .B(n1841), .C(n1845), .Y(n2859) );
  OAI21X1 U950 ( .A(n1840), .B(n1740), .C(n2464), .Y(n1951) );
  NAND2X1 U951 ( .A(\mem<5><0> ), .B(n1742), .Y(n2464) );
  OAI21X1 U952 ( .A(n1839), .B(n1740), .C(n2463), .Y(n1950) );
  NAND2X1 U953 ( .A(\mem<5><1> ), .B(n1742), .Y(n2463) );
  OAI21X1 U954 ( .A(n1838), .B(n1740), .C(n2462), .Y(n1949) );
  NAND2X1 U955 ( .A(\mem<5><2> ), .B(n1742), .Y(n2462) );
  OAI21X1 U956 ( .A(n1837), .B(n1740), .C(n2461), .Y(n1948) );
  NAND2X1 U957 ( .A(\mem<5><3> ), .B(n1742), .Y(n2461) );
  OAI21X1 U958 ( .A(n1836), .B(n1740), .C(n2460), .Y(n1947) );
  NAND2X1 U959 ( .A(\mem<5><4> ), .B(n1742), .Y(n2460) );
  OAI21X1 U960 ( .A(n1835), .B(n1740), .C(n2459), .Y(n1946) );
  NAND2X1 U961 ( .A(\mem<5><5> ), .B(n1742), .Y(n2459) );
  OAI21X1 U962 ( .A(n1834), .B(n1740), .C(n2458), .Y(n1945) );
  NAND2X1 U963 ( .A(\mem<5><6> ), .B(n1742), .Y(n2458) );
  OAI21X1 U964 ( .A(n1833), .B(n1740), .C(n2457), .Y(n1944) );
  NAND2X1 U965 ( .A(\mem<5><7> ), .B(n1742), .Y(n2457) );
  OAI21X1 U966 ( .A(n1832), .B(n1740), .C(n2456), .Y(n1943) );
  NAND2X1 U967 ( .A(\mem<5><8> ), .B(n1741), .Y(n2456) );
  OAI21X1 U968 ( .A(n1831), .B(n1740), .C(n2455), .Y(n1942) );
  NAND2X1 U969 ( .A(\mem<5><9> ), .B(n1741), .Y(n2455) );
  OAI21X1 U970 ( .A(n1830), .B(n1740), .C(n2454), .Y(n1941) );
  NAND2X1 U971 ( .A(\mem<5><10> ), .B(n1741), .Y(n2454) );
  OAI21X1 U972 ( .A(n1829), .B(n1740), .C(n2453), .Y(n1940) );
  NAND2X1 U973 ( .A(\mem<5><11> ), .B(n1741), .Y(n2453) );
  OAI21X1 U974 ( .A(n1828), .B(n1740), .C(n2452), .Y(n1939) );
  NAND2X1 U975 ( .A(\mem<5><12> ), .B(n1741), .Y(n2452) );
  OAI21X1 U976 ( .A(n1827), .B(n1740), .C(n2451), .Y(n1938) );
  NAND2X1 U977 ( .A(\mem<5><13> ), .B(n1741), .Y(n2451) );
  OAI21X1 U978 ( .A(n1826), .B(n1740), .C(n2450), .Y(n1937) );
  NAND2X1 U979 ( .A(\mem<5><14> ), .B(n1741), .Y(n2450) );
  OAI21X1 U980 ( .A(n1825), .B(n1740), .C(n2449), .Y(n1936) );
  NAND2X1 U981 ( .A(\mem<5><15> ), .B(n1741), .Y(n2449) );
  NOR3X1 U984 ( .A(n1842), .B(n1843), .C(n1845), .Y(n2842) );
  OAI21X1 U985 ( .A(n1840), .B(n1737), .C(n2448), .Y(n1935) );
  NAND2X1 U986 ( .A(\mem<4><0> ), .B(n1739), .Y(n2448) );
  OAI21X1 U987 ( .A(n1839), .B(n1737), .C(n2447), .Y(n1934) );
  NAND2X1 U988 ( .A(\mem<4><1> ), .B(n1739), .Y(n2447) );
  OAI21X1 U989 ( .A(n1838), .B(n1737), .C(n2446), .Y(n1933) );
  NAND2X1 U990 ( .A(\mem<4><2> ), .B(n1739), .Y(n2446) );
  OAI21X1 U991 ( .A(n1837), .B(n1737), .C(n2445), .Y(n1932) );
  NAND2X1 U992 ( .A(\mem<4><3> ), .B(n1739), .Y(n2445) );
  OAI21X1 U993 ( .A(n1836), .B(n1737), .C(n2444), .Y(n1931) );
  NAND2X1 U994 ( .A(\mem<4><4> ), .B(n1739), .Y(n2444) );
  OAI21X1 U995 ( .A(n1835), .B(n1737), .C(n2443), .Y(n1930) );
  NAND2X1 U996 ( .A(\mem<4><5> ), .B(n1739), .Y(n2443) );
  OAI21X1 U997 ( .A(n1834), .B(n1737), .C(n2442), .Y(n1929) );
  NAND2X1 U998 ( .A(\mem<4><6> ), .B(n1739), .Y(n2442) );
  OAI21X1 U999 ( .A(n1833), .B(n1737), .C(n2441), .Y(n1928) );
  NAND2X1 U1000 ( .A(\mem<4><7> ), .B(n1739), .Y(n2441) );
  OAI21X1 U1001 ( .A(n1832), .B(n1737), .C(n2440), .Y(n1927) );
  NAND2X1 U1002 ( .A(\mem<4><8> ), .B(n1738), .Y(n2440) );
  OAI21X1 U1003 ( .A(n1831), .B(n1737), .C(n2439), .Y(n1926) );
  NAND2X1 U1004 ( .A(\mem<4><9> ), .B(n1738), .Y(n2439) );
  OAI21X1 U1005 ( .A(n1830), .B(n1737), .C(n2438), .Y(n1925) );
  NAND2X1 U1006 ( .A(\mem<4><10> ), .B(n1738), .Y(n2438) );
  OAI21X1 U1007 ( .A(n1829), .B(n1737), .C(n2437), .Y(n1924) );
  NAND2X1 U1008 ( .A(\mem<4><11> ), .B(n1738), .Y(n2437) );
  OAI21X1 U1009 ( .A(n1828), .B(n1737), .C(n2436), .Y(n1923) );
  NAND2X1 U1010 ( .A(\mem<4><12> ), .B(n1738), .Y(n2436) );
  OAI21X1 U1011 ( .A(n1827), .B(n1737), .C(n2435), .Y(n1922) );
  NAND2X1 U1012 ( .A(\mem<4><13> ), .B(n1738), .Y(n2435) );
  OAI21X1 U1013 ( .A(n1826), .B(n1737), .C(n2434), .Y(n1921) );
  NAND2X1 U1014 ( .A(\mem<4><14> ), .B(n1738), .Y(n2434) );
  OAI21X1 U1015 ( .A(n1825), .B(n1737), .C(n2433), .Y(n1920) );
  NAND2X1 U1016 ( .A(\mem<4><15> ), .B(n1738), .Y(n2433) );
  NOR3X1 U1019 ( .A(n1841), .B(n1843), .C(n1845), .Y(n2825) );
  OAI21X1 U1020 ( .A(n1840), .B(n1734), .C(n2432), .Y(n1919) );
  NAND2X1 U1021 ( .A(\mem<3><0> ), .B(n1736), .Y(n2432) );
  OAI21X1 U1022 ( .A(n1839), .B(n1734), .C(n2431), .Y(n1918) );
  NAND2X1 U1023 ( .A(\mem<3><1> ), .B(n1736), .Y(n2431) );
  OAI21X1 U1024 ( .A(n1838), .B(n1734), .C(n2430), .Y(n1917) );
  NAND2X1 U1025 ( .A(\mem<3><2> ), .B(n1736), .Y(n2430) );
  OAI21X1 U1026 ( .A(n1837), .B(n1734), .C(n2429), .Y(n1916) );
  NAND2X1 U1027 ( .A(\mem<3><3> ), .B(n1736), .Y(n2429) );
  OAI21X1 U1028 ( .A(n1836), .B(n1734), .C(n2428), .Y(n1915) );
  NAND2X1 U1029 ( .A(\mem<3><4> ), .B(n1736), .Y(n2428) );
  OAI21X1 U1030 ( .A(n1835), .B(n1734), .C(n2427), .Y(n1914) );
  NAND2X1 U1031 ( .A(\mem<3><5> ), .B(n1736), .Y(n2427) );
  OAI21X1 U1032 ( .A(n1834), .B(n1734), .C(n2426), .Y(n1913) );
  NAND2X1 U1033 ( .A(\mem<3><6> ), .B(n1736), .Y(n2426) );
  OAI21X1 U1034 ( .A(n1833), .B(n1734), .C(n2425), .Y(n1912) );
  NAND2X1 U1035 ( .A(\mem<3><7> ), .B(n1736), .Y(n2425) );
  OAI21X1 U1036 ( .A(n1832), .B(n1734), .C(n2424), .Y(n1911) );
  NAND2X1 U1037 ( .A(\mem<3><8> ), .B(n1735), .Y(n2424) );
  OAI21X1 U1038 ( .A(n1831), .B(n1734), .C(n2423), .Y(n1910) );
  NAND2X1 U1039 ( .A(\mem<3><9> ), .B(n1735), .Y(n2423) );
  OAI21X1 U1040 ( .A(n1830), .B(n1734), .C(n2422), .Y(n1909) );
  NAND2X1 U1041 ( .A(\mem<3><10> ), .B(n1735), .Y(n2422) );
  OAI21X1 U1042 ( .A(n1829), .B(n1734), .C(n2421), .Y(n1908) );
  NAND2X1 U1043 ( .A(\mem<3><11> ), .B(n1735), .Y(n2421) );
  OAI21X1 U1044 ( .A(n1828), .B(n1734), .C(n2420), .Y(n1907) );
  NAND2X1 U1045 ( .A(\mem<3><12> ), .B(n1735), .Y(n2420) );
  OAI21X1 U1046 ( .A(n1827), .B(n1734), .C(n2419), .Y(n1906) );
  NAND2X1 U1047 ( .A(\mem<3><13> ), .B(n1735), .Y(n2419) );
  OAI21X1 U1048 ( .A(n1826), .B(n1734), .C(n2418), .Y(n1905) );
  NAND2X1 U1049 ( .A(\mem<3><14> ), .B(n1735), .Y(n2418) );
  OAI21X1 U1050 ( .A(n1825), .B(n1734), .C(n2417), .Y(n1904) );
  NAND2X1 U1051 ( .A(\mem<3><15> ), .B(n1735), .Y(n2417) );
  NOR3X1 U1054 ( .A(n1842), .B(n1688), .C(n1844), .Y(n2808) );
  OAI21X1 U1055 ( .A(n1840), .B(n1731), .C(n2416), .Y(n1903) );
  NAND2X1 U1056 ( .A(\mem<2><0> ), .B(n1733), .Y(n2416) );
  OAI21X1 U1057 ( .A(n1839), .B(n1731), .C(n2415), .Y(n1902) );
  NAND2X1 U1058 ( .A(\mem<2><1> ), .B(n1733), .Y(n2415) );
  OAI21X1 U1059 ( .A(n1838), .B(n1731), .C(n2414), .Y(n1901) );
  NAND2X1 U1060 ( .A(\mem<2><2> ), .B(n1733), .Y(n2414) );
  OAI21X1 U1061 ( .A(n1837), .B(n1731), .C(n2413), .Y(n1900) );
  NAND2X1 U1062 ( .A(\mem<2><3> ), .B(n1733), .Y(n2413) );
  OAI21X1 U1063 ( .A(n1836), .B(n1731), .C(n2412), .Y(n1899) );
  NAND2X1 U1064 ( .A(\mem<2><4> ), .B(n1733), .Y(n2412) );
  OAI21X1 U1065 ( .A(n1835), .B(n1731), .C(n2411), .Y(n1898) );
  NAND2X1 U1066 ( .A(\mem<2><5> ), .B(n1733), .Y(n2411) );
  OAI21X1 U1067 ( .A(n1834), .B(n1731), .C(n2410), .Y(n1897) );
  NAND2X1 U1068 ( .A(\mem<2><6> ), .B(n1733), .Y(n2410) );
  OAI21X1 U1069 ( .A(n1833), .B(n1731), .C(n2409), .Y(n1896) );
  NAND2X1 U1070 ( .A(\mem<2><7> ), .B(n1733), .Y(n2409) );
  OAI21X1 U1071 ( .A(n1832), .B(n1731), .C(n2408), .Y(n1895) );
  NAND2X1 U1072 ( .A(\mem<2><8> ), .B(n1732), .Y(n2408) );
  OAI21X1 U1073 ( .A(n1831), .B(n1731), .C(n2407), .Y(n1894) );
  NAND2X1 U1074 ( .A(\mem<2><9> ), .B(n1732), .Y(n2407) );
  OAI21X1 U1075 ( .A(n1830), .B(n1731), .C(n2406), .Y(n1893) );
  NAND2X1 U1076 ( .A(\mem<2><10> ), .B(n1732), .Y(n2406) );
  OAI21X1 U1077 ( .A(n1829), .B(n1731), .C(n2405), .Y(n1892) );
  NAND2X1 U1078 ( .A(\mem<2><11> ), .B(n1732), .Y(n2405) );
  OAI21X1 U1079 ( .A(n1828), .B(n1731), .C(n2404), .Y(n1891) );
  NAND2X1 U1080 ( .A(\mem<2><12> ), .B(n1732), .Y(n2404) );
  OAI21X1 U1081 ( .A(n1827), .B(n1731), .C(n2403), .Y(n1890) );
  NAND2X1 U1082 ( .A(\mem<2><13> ), .B(n1732), .Y(n2403) );
  OAI21X1 U1083 ( .A(n1826), .B(n1731), .C(n2402), .Y(n1889) );
  NAND2X1 U1084 ( .A(\mem<2><14> ), .B(n1732), .Y(n2402) );
  OAI21X1 U1085 ( .A(n1825), .B(n1731), .C(n2401), .Y(n1888) );
  NAND2X1 U1086 ( .A(\mem<2><15> ), .B(n1732), .Y(n2401) );
  NOR3X1 U1089 ( .A(n1841), .B(n1688), .C(n1844), .Y(n2791) );
  OAI21X1 U1090 ( .A(n1840), .B(n1728), .C(n2400), .Y(n1887) );
  NAND2X1 U1091 ( .A(\mem<1><0> ), .B(n1730), .Y(n2400) );
  OAI21X1 U1092 ( .A(n1839), .B(n1728), .C(n2399), .Y(n1886) );
  NAND2X1 U1093 ( .A(\mem<1><1> ), .B(n1730), .Y(n2399) );
  OAI21X1 U1094 ( .A(n1838), .B(n1728), .C(n2398), .Y(n1885) );
  NAND2X1 U1095 ( .A(\mem<1><2> ), .B(n1730), .Y(n2398) );
  OAI21X1 U1096 ( .A(n1837), .B(n1728), .C(n2397), .Y(n1884) );
  NAND2X1 U1097 ( .A(\mem<1><3> ), .B(n1730), .Y(n2397) );
  OAI21X1 U1098 ( .A(n1836), .B(n1728), .C(n2396), .Y(n1883) );
  NAND2X1 U1099 ( .A(\mem<1><4> ), .B(n1730), .Y(n2396) );
  OAI21X1 U1100 ( .A(n1835), .B(n1728), .C(n2395), .Y(n1882) );
  NAND2X1 U1101 ( .A(\mem<1><5> ), .B(n1730), .Y(n2395) );
  OAI21X1 U1102 ( .A(n1834), .B(n1728), .C(n2394), .Y(n1881) );
  NAND2X1 U1103 ( .A(\mem<1><6> ), .B(n1730), .Y(n2394) );
  OAI21X1 U1104 ( .A(n1833), .B(n1728), .C(n2393), .Y(n1880) );
  NAND2X1 U1105 ( .A(\mem<1><7> ), .B(n1730), .Y(n2393) );
  OAI21X1 U1106 ( .A(n1832), .B(n1728), .C(n2392), .Y(n1879) );
  NAND2X1 U1107 ( .A(\mem<1><8> ), .B(n1729), .Y(n2392) );
  OAI21X1 U1108 ( .A(n1831), .B(n1728), .C(n2391), .Y(n1878) );
  NAND2X1 U1109 ( .A(\mem<1><9> ), .B(n1729), .Y(n2391) );
  OAI21X1 U1110 ( .A(n1830), .B(n1728), .C(n2390), .Y(n1877) );
  NAND2X1 U1111 ( .A(\mem<1><10> ), .B(n1729), .Y(n2390) );
  OAI21X1 U1112 ( .A(n1829), .B(n1728), .C(n2389), .Y(n1876) );
  NAND2X1 U1113 ( .A(\mem<1><11> ), .B(n1729), .Y(n2389) );
  OAI21X1 U1114 ( .A(n1828), .B(n1728), .C(n2388), .Y(n1875) );
  NAND2X1 U1115 ( .A(\mem<1><12> ), .B(n1729), .Y(n2388) );
  OAI21X1 U1116 ( .A(n1827), .B(n1728), .C(n2387), .Y(n1874) );
  NAND2X1 U1117 ( .A(\mem<1><13> ), .B(n1729), .Y(n2387) );
  OAI21X1 U1118 ( .A(n1826), .B(n1728), .C(n2386), .Y(n1873) );
  NAND2X1 U1119 ( .A(\mem<1><14> ), .B(n1729), .Y(n2386) );
  OAI21X1 U1120 ( .A(n1825), .B(n1728), .C(n2385), .Y(n1872) );
  NAND2X1 U1121 ( .A(\mem<1><15> ), .B(n1729), .Y(n2385) );
  NOR3X1 U1124 ( .A(n1843), .B(n1688), .C(n1842), .Y(n2774) );
  OAI21X1 U1125 ( .A(n1840), .B(n1725), .C(n2384), .Y(n1871) );
  NAND2X1 U1126 ( .A(\mem<0><0> ), .B(n1727), .Y(n2384) );
  OAI21X1 U1128 ( .A(n1839), .B(n1725), .C(n2383), .Y(n1870) );
  NAND2X1 U1129 ( .A(\mem<0><1> ), .B(n1727), .Y(n2383) );
  OAI21X1 U1131 ( .A(n1838), .B(n1725), .C(n2382), .Y(n1869) );
  NAND2X1 U1132 ( .A(\mem<0><2> ), .B(n1727), .Y(n2382) );
  OAI21X1 U1134 ( .A(n1837), .B(n1725), .C(n2381), .Y(n1868) );
  NAND2X1 U1135 ( .A(\mem<0><3> ), .B(n1727), .Y(n2381) );
  OAI21X1 U1137 ( .A(n1836), .B(n1725), .C(n2380), .Y(n1867) );
  NAND2X1 U1138 ( .A(\mem<0><4> ), .B(n1727), .Y(n2380) );
  OAI21X1 U1140 ( .A(n1835), .B(n1725), .C(n2379), .Y(n1866) );
  NAND2X1 U1141 ( .A(\mem<0><5> ), .B(n1727), .Y(n2379) );
  OAI21X1 U1143 ( .A(n1834), .B(n1725), .C(n2378), .Y(n1865) );
  NAND2X1 U1144 ( .A(\mem<0><6> ), .B(n1727), .Y(n2378) );
  OAI21X1 U1146 ( .A(n1833), .B(n1725), .C(n2377), .Y(n1864) );
  NAND2X1 U1147 ( .A(\mem<0><7> ), .B(n1727), .Y(n2377) );
  OAI21X1 U1149 ( .A(n1832), .B(n1725), .C(n2376), .Y(n1863) );
  NAND2X1 U1150 ( .A(\mem<0><8> ), .B(n1726), .Y(n2376) );
  OAI21X1 U1152 ( .A(n1831), .B(n1725), .C(n2375), .Y(n1862) );
  NAND2X1 U1153 ( .A(\mem<0><9> ), .B(n1726), .Y(n2375) );
  OAI21X1 U1155 ( .A(n1830), .B(n1725), .C(n2374), .Y(n1861) );
  NAND2X1 U1156 ( .A(\mem<0><10> ), .B(n1726), .Y(n2374) );
  OAI21X1 U1158 ( .A(n1829), .B(n1725), .C(n2373), .Y(n1860) );
  NAND2X1 U1159 ( .A(\mem<0><11> ), .B(n1726), .Y(n2373) );
  OAI21X1 U1161 ( .A(n1828), .B(n1725), .C(n2372), .Y(n1859) );
  NAND2X1 U1162 ( .A(\mem<0><12> ), .B(n1726), .Y(n2372) );
  OAI21X1 U1164 ( .A(n1827), .B(n1725), .C(n2371), .Y(n1858) );
  NAND2X1 U1165 ( .A(\mem<0><13> ), .B(n1726), .Y(n2371) );
  OAI21X1 U1167 ( .A(n1826), .B(n1725), .C(n2370), .Y(n1857) );
  NAND2X1 U1168 ( .A(\mem<0><14> ), .B(n1726), .Y(n2370) );
  OAI21X1 U1170 ( .A(n1825), .B(n1725), .C(n2369), .Y(n1856) );
  NAND2X1 U1171 ( .A(\mem<0><15> ), .B(n1726), .Y(n2369) );
  NOR3X1 U1174 ( .A(n1843), .B(n1688), .C(n1841), .Y(n2757) );
  NAND3X1 U1175 ( .A(n1847), .B(n1849), .C(n2755), .Y(n2368) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2755) );
  AND2X2 U3 ( .A(\data_in<9> ), .B(n1821), .Y(n47) );
  AND2X2 U4 ( .A(\data_in<15> ), .B(n1821), .Y(n39) );
  AND2X2 U5 ( .A(\data_in<0> ), .B(n1823), .Y(n64) );
  INVX8 U6 ( .A(n64), .Y(n1840) );
  AND2X2 U7 ( .A(\data_in<2> ), .B(n1823), .Y(n60) );
  INVX8 U8 ( .A(n60), .Y(n1838) );
  AND2X2 U9 ( .A(\data_in<3> ), .B(n1823), .Y(n58) );
  AND2X2 U10 ( .A(\data_in<4> ), .B(n1823), .Y(n56) );
  INVX8 U11 ( .A(n56), .Y(n1836) );
  AND2X2 U12 ( .A(\data_in<5> ), .B(n1823), .Y(n54) );
  AND2X2 U13 ( .A(\data_in<6> ), .B(n1823), .Y(n52) );
  INVX8 U14 ( .A(n52), .Y(n1834) );
  AND2X2 U15 ( .A(\data_in<7> ), .B(n1823), .Y(n50) );
  AND2X2 U16 ( .A(\data_in<13> ), .B(n1823), .Y(n42) );
  AND2X2 U17 ( .A(\data_in<11> ), .B(n1822), .Y(n44) );
  INVX2 U18 ( .A(n1708), .Y(n1711) );
  INVX2 U19 ( .A(n1708), .Y(n1710) );
  INVX1 U20 ( .A(n1842), .Y(n1718) );
  INVX1 U21 ( .A(n1842), .Y(n1719) );
  INVX1 U22 ( .A(n1842), .Y(n1720) );
  INVX1 U23 ( .A(n1841), .Y(n1707) );
  INVX1 U24 ( .A(n1842), .Y(n1724) );
  INVX2 U25 ( .A(n1708), .Y(n1709) );
  INVX2 U26 ( .A(n1841), .Y(n1708) );
  INVX1 U27 ( .A(n1695), .Y(n1698) );
  INVX2 U28 ( .A(n1706), .Y(n1715) );
  INVX1 U29 ( .A(n1695), .Y(n1699) );
  INVX2 U30 ( .A(n1706), .Y(n1717) );
  INVX1 U31 ( .A(n1694), .Y(n1701) );
  INVX2 U32 ( .A(n1706), .Y(n1721) );
  INVX2 U33 ( .A(n1706), .Y(n1722) );
  INVX1 U34 ( .A(n1695), .Y(n1704) );
  INVX1 U35 ( .A(n1724), .Y(n1706) );
  INVX2 U36 ( .A(n1706), .Y(n1723) );
  INVX1 U37 ( .A(n1694), .Y(n1705) );
  INVX1 U38 ( .A(n1845), .Y(n1693) );
  INVX1 U39 ( .A(n1844), .Y(n1697) );
  INVX2 U40 ( .A(n1845), .Y(n1692) );
  INVX2 U41 ( .A(n1706), .Y(n1716) );
  INVX2 U42 ( .A(n1695), .Y(n1700) );
  INVX2 U43 ( .A(n1845), .Y(n1691) );
  INVX1 U44 ( .A(n1694), .Y(n1702) );
  INVX2 U45 ( .A(n1694), .Y(n1703) );
  INVX2 U46 ( .A(n1845), .Y(n1690) );
  INVX2 U47 ( .A(n1851), .Y(n1) );
  BUFX2 U48 ( .A(n1188), .Y(n1820) );
  BUFX2 U49 ( .A(n1188), .Y(n1819) );
  BUFX2 U50 ( .A(n1186), .Y(n1817) );
  BUFX2 U51 ( .A(n1186), .Y(n1816) );
  BUFX2 U52 ( .A(n1184), .Y(n1814) );
  BUFX2 U53 ( .A(n1184), .Y(n1813) );
  BUFX2 U54 ( .A(n1182), .Y(n1811) );
  BUFX2 U55 ( .A(n1182), .Y(n1810) );
  BUFX2 U56 ( .A(n1180), .Y(n1808) );
  BUFX2 U57 ( .A(n1180), .Y(n1807) );
  BUFX2 U58 ( .A(n1178), .Y(n1805) );
  BUFX2 U59 ( .A(n1178), .Y(n1804) );
  BUFX2 U60 ( .A(n1176), .Y(n1802) );
  BUFX2 U93 ( .A(n1176), .Y(n1801) );
  BUFX2 U94 ( .A(n1174), .Y(n1799) );
  BUFX2 U127 ( .A(n1174), .Y(n1798) );
  BUFX2 U128 ( .A(n1172), .Y(n1796) );
  BUFX2 U161 ( .A(n1172), .Y(n1795) );
  BUFX2 U162 ( .A(n1170), .Y(n1793) );
  BUFX2 U195 ( .A(n1170), .Y(n1792) );
  BUFX2 U196 ( .A(n1168), .Y(n1790) );
  BUFX2 U229 ( .A(n1168), .Y(n1789) );
  BUFX2 U230 ( .A(n1166), .Y(n1787) );
  BUFX2 U263 ( .A(n1166), .Y(n1786) );
  BUFX2 U264 ( .A(n1164), .Y(n1784) );
  BUFX2 U297 ( .A(n1164), .Y(n1783) );
  BUFX2 U298 ( .A(n650), .Y(n1781) );
  BUFX2 U331 ( .A(n650), .Y(n1780) );
  BUFX2 U332 ( .A(n631), .Y(n1778) );
  BUFX2 U366 ( .A(n631), .Y(n1777) );
  BUFX2 U367 ( .A(n613), .Y(n1775) );
  BUFX2 U400 ( .A(n613), .Y(n1774) );
  BUFX2 U401 ( .A(n595), .Y(n1772) );
  BUFX2 U434 ( .A(n595), .Y(n1771) );
  BUFX2 U435 ( .A(n577), .Y(n1769) );
  BUFX2 U468 ( .A(n577), .Y(n1768) );
  BUFX2 U469 ( .A(n559), .Y(n1766) );
  BUFX2 U502 ( .A(n559), .Y(n1765) );
  BUFX2 U503 ( .A(n541), .Y(n1763) );
  BUFX2 U536 ( .A(n541), .Y(n1762) );
  BUFX2 U537 ( .A(n523), .Y(n1760) );
  BUFX2 U570 ( .A(n523), .Y(n1759) );
  BUFX2 U571 ( .A(n505), .Y(n1757) );
  BUFX2 U604 ( .A(n505), .Y(n1756) );
  BUFX2 U605 ( .A(n486), .Y(n1754) );
  BUFX2 U639 ( .A(n486), .Y(n1753) );
  BUFX2 U640 ( .A(n468), .Y(n1751) );
  BUFX2 U673 ( .A(n468), .Y(n1750) );
  BUFX2 U674 ( .A(n450), .Y(n1748) );
  BUFX2 U707 ( .A(n450), .Y(n1747) );
  BUFX2 U708 ( .A(n432), .Y(n1745) );
  BUFX2 U741 ( .A(n432), .Y(n1744) );
  BUFX2 U742 ( .A(n414), .Y(n1742) );
  BUFX2 U775 ( .A(n414), .Y(n1741) );
  BUFX2 U776 ( .A(n396), .Y(n1739) );
  BUFX2 U809 ( .A(n396), .Y(n1738) );
  BUFX2 U810 ( .A(n378), .Y(n1736) );
  BUFX2 U843 ( .A(n378), .Y(n1735) );
  BUFX2 U844 ( .A(n360), .Y(n1733) );
  BUFX2 U877 ( .A(n360), .Y(n1732) );
  BUFX2 U878 ( .A(n341), .Y(n1730) );
  BUFX2 U912 ( .A(n341), .Y(n1729) );
  BUFX2 U913 ( .A(n323), .Y(n1727) );
  BUFX2 U947 ( .A(n323), .Y(n1726) );
  INVX2 U948 ( .A(n1845), .Y(n1688) );
  INVX1 U982 ( .A(n1844), .Y(n1696) );
  INVX1 U983 ( .A(n1842), .Y(n1841) );
  INVX1 U1017 ( .A(N12), .Y(n1845) );
  INVX1 U1018 ( .A(N14), .Y(n1849) );
  INVX1 U1052 ( .A(n1849), .Y(n1685) );
  INVX8 U1053 ( .A(n41), .Y(n1826) );
  INVX8 U1087 ( .A(n43), .Y(n1828) );
  INVX8 U1088 ( .A(n45), .Y(n1830) );
  INVX8 U1122 ( .A(n48), .Y(n1832) );
  INVX1 U1123 ( .A(rst), .Y(n1850) );
  INVX1 U1127 ( .A(N13), .Y(n1847) );
  INVX1 U1130 ( .A(n1844), .Y(n1843) );
  INVX1 U1133 ( .A(n40), .Y(n1725) );
  INVX1 U1136 ( .A(n1847), .Y(n1687) );
  INVX1 U1139 ( .A(n1847), .Y(n1686) );
  INVX1 U1142 ( .A(n66), .Y(n1728) );
  INVX1 U1145 ( .A(n99), .Y(n1752) );
  INVX1 U1148 ( .A(n175), .Y(n1776) );
  INVX1 U1151 ( .A(n68), .Y(n1731) );
  INVX1 U1154 ( .A(n70), .Y(n1734) );
  INVX1 U1157 ( .A(n72), .Y(n1737) );
  INVX1 U1160 ( .A(n74), .Y(n1740) );
  INVX1 U1163 ( .A(n76), .Y(n1743) );
  INVX1 U1166 ( .A(n80), .Y(n1746) );
  INVX1 U1169 ( .A(n82), .Y(n1749) );
  INVX1 U1172 ( .A(n101), .Y(n1755) );
  INVX1 U1173 ( .A(n118), .Y(n1758) );
  INVX1 U1177 ( .A(n120), .Y(n1761) );
  INVX1 U1178 ( .A(n137), .Y(n1764) );
  INVX1 U1179 ( .A(n139), .Y(n1767) );
  INVX1 U1180 ( .A(n156), .Y(n1770) );
  INVX1 U1181 ( .A(n158), .Y(n1773) );
  INVX1 U1182 ( .A(n177), .Y(n1779) );
  INVX1 U1183 ( .A(n194), .Y(n1782) );
  INVX1 U1184 ( .A(n196), .Y(n1785) );
  INVX1 U1185 ( .A(n215), .Y(n1788) );
  INVX1 U1186 ( .A(n217), .Y(n1791) );
  INVX1 U1187 ( .A(n233), .Y(n1794) );
  INVX1 U1188 ( .A(n235), .Y(n1797) );
  INVX1 U1189 ( .A(n251), .Y(n1800) );
  INVX1 U1190 ( .A(n253), .Y(n1803) );
  INVX1 U1191 ( .A(n269), .Y(n1806) );
  INVX1 U1192 ( .A(n271), .Y(n1809) );
  INVX1 U1193 ( .A(n287), .Y(n1812) );
  INVX1 U1194 ( .A(n289), .Y(n1815) );
  INVX1 U1195 ( .A(n305), .Y(n1818) );
  INVX1 U1196 ( .A(n1843), .Y(n1694) );
  INVX1 U1197 ( .A(n1843), .Y(n1695) );
  OR2X2 U1198 ( .A(n2), .B(n1682), .Y(n29) );
  OR2X2 U1199 ( .A(n2), .B(n1684), .Y(n33) );
  OR2X2 U1200 ( .A(n2), .B(n1679), .Y(n23) );
  OR2X2 U1201 ( .A(n2), .B(n1677), .Y(n19) );
  OR2X2 U1202 ( .A(n2), .B(n1669), .Y(n3) );
  OR2X2 U1203 ( .A(n2), .B(n1671), .Y(n7) );
  OR2X2 U1204 ( .A(n2), .B(n1673), .Y(n11) );
  OR2X2 U1205 ( .A(n2), .B(n1675), .Y(n15) );
  OR2X2 U1206 ( .A(n2), .B(n1683), .Y(n31) );
  OR2X2 U1207 ( .A(n2), .B(n1681), .Y(n27) );
  OR2X2 U1208 ( .A(n2), .B(n1672), .Y(n9) );
  OR2X2 U1209 ( .A(n2), .B(n1680), .Y(n25) );
  OR2X2 U1210 ( .A(n2), .B(n1678), .Y(n21) );
  OR2X2 U1211 ( .A(n2), .B(n1676), .Y(n17) );
  OR2X2 U1212 ( .A(n2), .B(n1674), .Y(n13) );
  OR2X2 U1213 ( .A(n2), .B(n1670), .Y(n5) );
  INVX8 U1214 ( .A(n1), .Y(n2) );
  INVX1 U1215 ( .A(n3), .Y(\data_out<0> ) );
  INVX1 U1216 ( .A(n5), .Y(\data_out<1> ) );
  INVX1 U1217 ( .A(n7), .Y(\data_out<2> ) );
  INVX1 U1218 ( .A(n9), .Y(\data_out<3> ) );
  INVX1 U1219 ( .A(n11), .Y(\data_out<4> ) );
  INVX1 U1220 ( .A(n13), .Y(\data_out<5> ) );
  INVX1 U1221 ( .A(n15), .Y(\data_out<6> ) );
  INVX1 U1222 ( .A(n17), .Y(\data_out<7> ) );
  INVX1 U1223 ( .A(n19), .Y(\data_out<8> ) );
  INVX1 U1224 ( .A(n21), .Y(\data_out<9> ) );
  INVX1 U1225 ( .A(n23), .Y(\data_out<10> ) );
  INVX1 U1226 ( .A(n25), .Y(\data_out<11> ) );
  INVX1 U1227 ( .A(n27), .Y(\data_out<12> ) );
  INVX1 U1228 ( .A(n29), .Y(\data_out<13> ) );
  INVX1 U1229 ( .A(n31), .Y(\data_out<14> ) );
  INVX1 U1230 ( .A(n33), .Y(\data_out<15> ) );
  INVX1 U1231 ( .A(n1849), .Y(n1848) );
  INVX1 U1232 ( .A(n1847), .Y(n1846) );
  BUFX2 U1233 ( .A(n2368), .Y(n35) );
  INVX1 U1234 ( .A(n35), .Y(n1852) );
  BUFX2 U1235 ( .A(n2497), .Y(n36) );
  INVX1 U1236 ( .A(n36), .Y(n1855) );
  BUFX2 U1237 ( .A(n2626), .Y(n37) );
  INVX1 U1238 ( .A(n37), .Y(n1853) );
  BUFX2 U1239 ( .A(n2756), .Y(n38) );
  INVX1 U1240 ( .A(n38), .Y(n1854) );
  AND2X1 U1241 ( .A(n1852), .B(n2757), .Y(n40) );
  AND2X1 U1242 ( .A(\data_in<14> ), .B(n1822), .Y(n41) );
  AND2X1 U1243 ( .A(\data_in<12> ), .B(n1821), .Y(n43) );
  AND2X1 U1244 ( .A(\data_in<10> ), .B(n1823), .Y(n45) );
  AND2X1 U1245 ( .A(\data_in<8> ), .B(n1822), .Y(n48) );
  AND2X1 U1246 ( .A(\data_in<1> ), .B(n1823), .Y(n62) );
  AND2X1 U1247 ( .A(n1852), .B(n2774), .Y(n66) );
  AND2X1 U1248 ( .A(n1852), .B(n2791), .Y(n68) );
  AND2X1 U1249 ( .A(n1852), .B(n2808), .Y(n70) );
  AND2X1 U1250 ( .A(n1852), .B(n2825), .Y(n72) );
  AND2X1 U1251 ( .A(n1852), .B(n2842), .Y(n74) );
  AND2X1 U1252 ( .A(n1852), .B(n2859), .Y(n76) );
  AND2X1 U1253 ( .A(n1852), .B(n2876), .Y(n80) );
  AND2X1 U1254 ( .A(n1855), .B(n2757), .Y(n82) );
  AND2X1 U1255 ( .A(n1855), .B(n2774), .Y(n99) );
  AND2X1 U1256 ( .A(n1855), .B(n2791), .Y(n101) );
  AND2X1 U1257 ( .A(n1855), .B(n2808), .Y(n118) );
  AND2X1 U1258 ( .A(n1855), .B(n2825), .Y(n120) );
  AND2X1 U1259 ( .A(n1855), .B(n2842), .Y(n137) );
  AND2X1 U1260 ( .A(n1855), .B(n2859), .Y(n139) );
  AND2X1 U1261 ( .A(n1855), .B(n2876), .Y(n156) );
  AND2X1 U1262 ( .A(n1853), .B(n2757), .Y(n158) );
  AND2X1 U1263 ( .A(n1853), .B(n2774), .Y(n175) );
  AND2X1 U1264 ( .A(n1853), .B(n2791), .Y(n177) );
  AND2X1 U1265 ( .A(n1853), .B(n2808), .Y(n194) );
  AND2X1 U1266 ( .A(n1853), .B(n2825), .Y(n196) );
  AND2X1 U1267 ( .A(n1853), .B(n2842), .Y(n215) );
  AND2X1 U1268 ( .A(n1853), .B(n2859), .Y(n217) );
  AND2X1 U1269 ( .A(n1853), .B(n2876), .Y(n233) );
  AND2X1 U1270 ( .A(n2757), .B(n1854), .Y(n235) );
  AND2X1 U1271 ( .A(n2774), .B(n1854), .Y(n251) );
  AND2X1 U1272 ( .A(n2791), .B(n1854), .Y(n253) );
  AND2X1 U1273 ( .A(n2808), .B(n1854), .Y(n269) );
  AND2X1 U1274 ( .A(n2825), .B(n1854), .Y(n271) );
  AND2X1 U1275 ( .A(n2842), .B(n1854), .Y(n287) );
  AND2X1 U1276 ( .A(n2859), .B(n1854), .Y(n289) );
  AND2X1 U1277 ( .A(n2876), .B(n1854), .Y(n305) );
  AND2X1 U1278 ( .A(n40), .B(n1823), .Y(n307) );
  INVX1 U1279 ( .A(n307), .Y(n323) );
  AND2X1 U1280 ( .A(n66), .B(n1823), .Y(n325) );
  INVX1 U1281 ( .A(n325), .Y(n341) );
  AND2X1 U1282 ( .A(n68), .B(n1823), .Y(n343) );
  INVX1 U1283 ( .A(n343), .Y(n360) );
  AND2X1 U1284 ( .A(n70), .B(n1823), .Y(n362) );
  INVX1 U1285 ( .A(n362), .Y(n378) );
  AND2X1 U1286 ( .A(n72), .B(n1823), .Y(n380) );
  INVX1 U1287 ( .A(n380), .Y(n396) );
  AND2X1 U1288 ( .A(n74), .B(n1823), .Y(n398) );
  INVX1 U1289 ( .A(n398), .Y(n414) );
  AND2X1 U1290 ( .A(n76), .B(n1822), .Y(n416) );
  INVX1 U1291 ( .A(n416), .Y(n432) );
  AND2X1 U1292 ( .A(n80), .B(n1822), .Y(n434) );
  INVX1 U1293 ( .A(n434), .Y(n450) );
  AND2X1 U1294 ( .A(n82), .B(n1822), .Y(n452) );
  INVX1 U1295 ( .A(n452), .Y(n468) );
  AND2X1 U1296 ( .A(n99), .B(n1822), .Y(n470) );
  INVX1 U1297 ( .A(n470), .Y(n486) );
  AND2X1 U1298 ( .A(n101), .B(n1822), .Y(n488) );
  INVX1 U1299 ( .A(n488), .Y(n505) );
  AND2X1 U1300 ( .A(n118), .B(n1822), .Y(n507) );
  INVX1 U1301 ( .A(n507), .Y(n523) );
  AND2X1 U1302 ( .A(n120), .B(n1822), .Y(n525) );
  INVX1 U1303 ( .A(n525), .Y(n541) );
  AND2X1 U1304 ( .A(n137), .B(n1822), .Y(n543) );
  INVX1 U1305 ( .A(n543), .Y(n559) );
  AND2X1 U1306 ( .A(n139), .B(n1822), .Y(n561) );
  INVX1 U1307 ( .A(n561), .Y(n577) );
  AND2X1 U1308 ( .A(n156), .B(n1822), .Y(n579) );
  INVX1 U1309 ( .A(n579), .Y(n595) );
  AND2X1 U1310 ( .A(n158), .B(n1822), .Y(n597) );
  INVX1 U1311 ( .A(n597), .Y(n613) );
  AND2X1 U1312 ( .A(n175), .B(n1822), .Y(n615) );
  INVX1 U1313 ( .A(n615), .Y(n631) );
  AND2X1 U1314 ( .A(n177), .B(n1822), .Y(n633) );
  INVX1 U1315 ( .A(n633), .Y(n650) );
  AND2X1 U1316 ( .A(n194), .B(n1821), .Y(n1163) );
  INVX1 U1317 ( .A(n1163), .Y(n1164) );
  AND2X1 U1318 ( .A(n196), .B(n1821), .Y(n1165) );
  INVX1 U1319 ( .A(n1165), .Y(n1166) );
  AND2X1 U1320 ( .A(n215), .B(n1821), .Y(n1167) );
  INVX1 U1321 ( .A(n1167), .Y(n1168) );
  AND2X1 U1322 ( .A(n217), .B(n1821), .Y(n1169) );
  INVX1 U1323 ( .A(n1169), .Y(n1170) );
  AND2X1 U1324 ( .A(n233), .B(n1821), .Y(n1171) );
  INVX1 U1325 ( .A(n1171), .Y(n1172) );
  AND2X1 U1326 ( .A(n235), .B(n1821), .Y(n1173) );
  INVX1 U1327 ( .A(n1173), .Y(n1174) );
  AND2X1 U1328 ( .A(n251), .B(n1821), .Y(n1175) );
  INVX1 U1329 ( .A(n1175), .Y(n1176) );
  AND2X1 U1330 ( .A(n253), .B(n1821), .Y(n1177) );
  INVX1 U1331 ( .A(n1177), .Y(n1178) );
  AND2X1 U1332 ( .A(n269), .B(n1821), .Y(n1179) );
  INVX1 U1333 ( .A(n1179), .Y(n1180) );
  AND2X1 U1334 ( .A(n271), .B(n1821), .Y(n1181) );
  INVX1 U1335 ( .A(n1181), .Y(n1182) );
  AND2X1 U1336 ( .A(n287), .B(n1821), .Y(n1183) );
  INVX1 U1337 ( .A(n1183), .Y(n1184) );
  AND2X1 U1338 ( .A(n289), .B(n1821), .Y(n1185) );
  INVX1 U1339 ( .A(n1185), .Y(n1186) );
  AND2X1 U1340 ( .A(n305), .B(n1821), .Y(n1187) );
  INVX1 U1341 ( .A(n1187), .Y(n1188) );
  MUX2X1 U1342 ( .B(n1190), .A(n1191), .S(n1696), .Y(n1189) );
  MUX2X1 U1343 ( .B(n1193), .A(n1194), .S(n1696), .Y(n1192) );
  MUX2X1 U1344 ( .B(n1196), .A(n1197), .S(n1696), .Y(n1195) );
  MUX2X1 U1345 ( .B(n1199), .A(n1200), .S(n1696), .Y(n1198) );
  MUX2X1 U1346 ( .B(n1202), .A(n1203), .S(n1687), .Y(n1201) );
  MUX2X1 U1347 ( .B(n1205), .A(n1206), .S(n1696), .Y(n1204) );
  MUX2X1 U1348 ( .B(n1208), .A(n1209), .S(n1696), .Y(n1207) );
  MUX2X1 U1349 ( .B(n1211), .A(n1212), .S(n1696), .Y(n1210) );
  MUX2X1 U1350 ( .B(n1214), .A(n1215), .S(n1696), .Y(n1213) );
  MUX2X1 U1351 ( .B(n1217), .A(n1218), .S(n1687), .Y(n1216) );
  MUX2X1 U1352 ( .B(n1220), .A(n1221), .S(n1697), .Y(n1219) );
  MUX2X1 U1353 ( .B(n1223), .A(n1224), .S(n1697), .Y(n1222) );
  MUX2X1 U1354 ( .B(n1226), .A(n1227), .S(n1697), .Y(n1225) );
  MUX2X1 U1355 ( .B(n1229), .A(n1230), .S(n1697), .Y(n1228) );
  MUX2X1 U1356 ( .B(n1232), .A(n1233), .S(n1687), .Y(n1231) );
  MUX2X1 U1357 ( .B(n1235), .A(n1236), .S(n1697), .Y(n1234) );
  MUX2X1 U1358 ( .B(n1238), .A(n1239), .S(n1697), .Y(n1237) );
  MUX2X1 U1359 ( .B(n1241), .A(n1242), .S(n1697), .Y(n1240) );
  MUX2X1 U1360 ( .B(n1244), .A(n1245), .S(n1697), .Y(n1243) );
  MUX2X1 U1361 ( .B(n1247), .A(n1248), .S(n1687), .Y(n1246) );
  MUX2X1 U1362 ( .B(n1250), .A(n1251), .S(n1697), .Y(n1249) );
  MUX2X1 U1363 ( .B(n1253), .A(n1254), .S(n1697), .Y(n1252) );
  MUX2X1 U1364 ( .B(n1256), .A(n1257), .S(n1697), .Y(n1255) );
  MUX2X1 U1365 ( .B(n1259), .A(n1260), .S(n1697), .Y(n1258) );
  MUX2X1 U1366 ( .B(n1262), .A(n1263), .S(n1687), .Y(n1261) );
  MUX2X1 U1367 ( .B(n1265), .A(n1266), .S(n1697), .Y(n1264) );
  MUX2X1 U1368 ( .B(n1268), .A(n1269), .S(n1696), .Y(n1267) );
  MUX2X1 U1369 ( .B(n1271), .A(n1272), .S(n1697), .Y(n1270) );
  MUX2X1 U1370 ( .B(n1274), .A(n1275), .S(n1696), .Y(n1273) );
  MUX2X1 U1371 ( .B(n1277), .A(n1278), .S(n1687), .Y(n1276) );
  MUX2X1 U1372 ( .B(n1280), .A(n1281), .S(n1696), .Y(n1279) );
  MUX2X1 U1373 ( .B(n1283), .A(n1284), .S(n1696), .Y(n1282) );
  MUX2X1 U1374 ( .B(n1286), .A(n1287), .S(n1697), .Y(n1285) );
  MUX2X1 U1375 ( .B(n1289), .A(n1290), .S(n1696), .Y(n1288) );
  MUX2X1 U1376 ( .B(n1292), .A(n1293), .S(n1687), .Y(n1291) );
  MUX2X1 U1377 ( .B(n1295), .A(n1296), .S(n1697), .Y(n1294) );
  MUX2X1 U1378 ( .B(n1298), .A(n1299), .S(n1697), .Y(n1297) );
  MUX2X1 U1379 ( .B(n1301), .A(n1302), .S(n1697), .Y(n1300) );
  MUX2X1 U1380 ( .B(n1304), .A(n1305), .S(n1697), .Y(n1303) );
  MUX2X1 U1381 ( .B(n1307), .A(n1308), .S(n1687), .Y(n1306) );
  MUX2X1 U1382 ( .B(n1310), .A(n1311), .S(n1698), .Y(n1309) );
  MUX2X1 U1383 ( .B(n1313), .A(n1314), .S(n1698), .Y(n1312) );
  MUX2X1 U1384 ( .B(n1316), .A(n1317), .S(n1698), .Y(n1315) );
  MUX2X1 U1385 ( .B(n1319), .A(n1320), .S(n1698), .Y(n1318) );
  MUX2X1 U1386 ( .B(n1322), .A(n1323), .S(n1687), .Y(n1321) );
  MUX2X1 U1387 ( .B(n1325), .A(n1326), .S(n1698), .Y(n1324) );
  MUX2X1 U1388 ( .B(n1328), .A(n1329), .S(n1698), .Y(n1327) );
  MUX2X1 U1389 ( .B(n1331), .A(n1332), .S(n1698), .Y(n1330) );
  MUX2X1 U1390 ( .B(n1334), .A(n1335), .S(n1698), .Y(n1333) );
  MUX2X1 U1391 ( .B(n1337), .A(n1338), .S(n1687), .Y(n1336) );
  MUX2X1 U1392 ( .B(n1340), .A(n1341), .S(n1698), .Y(n1339) );
  MUX2X1 U1393 ( .B(n1343), .A(n1344), .S(n1698), .Y(n1342) );
  MUX2X1 U1394 ( .B(n1346), .A(n1347), .S(n1698), .Y(n1345) );
  MUX2X1 U1395 ( .B(n1349), .A(n1350), .S(n1698), .Y(n1348) );
  MUX2X1 U1396 ( .B(n1352), .A(n1353), .S(n1687), .Y(n1351) );
  MUX2X1 U1397 ( .B(n1355), .A(n1356), .S(n1699), .Y(n1354) );
  MUX2X1 U1398 ( .B(n1358), .A(n1359), .S(n1699), .Y(n1357) );
  MUX2X1 U1399 ( .B(n1361), .A(n1362), .S(n1699), .Y(n1360) );
  MUX2X1 U1400 ( .B(n1364), .A(n1365), .S(n1699), .Y(n1363) );
  MUX2X1 U1401 ( .B(n1367), .A(n1368), .S(n1687), .Y(n1366) );
  MUX2X1 U1402 ( .B(n1370), .A(n1371), .S(n1699), .Y(n1369) );
  MUX2X1 U1403 ( .B(n1373), .A(n1374), .S(n1699), .Y(n1372) );
  MUX2X1 U1404 ( .B(n1376), .A(n1377), .S(n1699), .Y(n1375) );
  MUX2X1 U1405 ( .B(n1379), .A(n1380), .S(n1699), .Y(n1378) );
  MUX2X1 U1406 ( .B(n1382), .A(n1383), .S(n1686), .Y(n1381) );
  MUX2X1 U1407 ( .B(n1385), .A(n1386), .S(n1699), .Y(n1384) );
  MUX2X1 U1408 ( .B(n1388), .A(n1389), .S(n1699), .Y(n1387) );
  MUX2X1 U1409 ( .B(n1391), .A(n1392), .S(n1699), .Y(n1390) );
  MUX2X1 U1410 ( .B(n1394), .A(n1395), .S(n1699), .Y(n1393) );
  MUX2X1 U1411 ( .B(n1397), .A(n1398), .S(n1686), .Y(n1396) );
  MUX2X1 U1412 ( .B(n1400), .A(n1401), .S(n1700), .Y(n1399) );
  MUX2X1 U1413 ( .B(n1403), .A(n1404), .S(n1700), .Y(n1402) );
  MUX2X1 U1414 ( .B(n1406), .A(n1407), .S(n1700), .Y(n1405) );
  MUX2X1 U1415 ( .B(n1409), .A(n1410), .S(n1700), .Y(n1408) );
  MUX2X1 U1416 ( .B(n1412), .A(n1413), .S(n1686), .Y(n1411) );
  MUX2X1 U1417 ( .B(n1415), .A(n1416), .S(n1700), .Y(n1414) );
  MUX2X1 U1418 ( .B(n1418), .A(n1419), .S(n1700), .Y(n1417) );
  MUX2X1 U1419 ( .B(n1421), .A(n1422), .S(n1700), .Y(n1420) );
  MUX2X1 U1420 ( .B(n1424), .A(n1425), .S(n1700), .Y(n1423) );
  MUX2X1 U1421 ( .B(n1427), .A(n1428), .S(n1686), .Y(n1426) );
  MUX2X1 U1422 ( .B(n1430), .A(n1431), .S(n1700), .Y(n1429) );
  MUX2X1 U1423 ( .B(n1433), .A(n1434), .S(n1700), .Y(n1432) );
  MUX2X1 U1424 ( .B(n1436), .A(n1437), .S(n1700), .Y(n1435) );
  MUX2X1 U1425 ( .B(n1439), .A(n1440), .S(n1700), .Y(n1438) );
  MUX2X1 U1426 ( .B(n1442), .A(n1443), .S(n1686), .Y(n1441) );
  MUX2X1 U1427 ( .B(n1445), .A(n1446), .S(n1701), .Y(n1444) );
  MUX2X1 U1428 ( .B(n1448), .A(n1449), .S(n1701), .Y(n1447) );
  MUX2X1 U1429 ( .B(n1451), .A(n1452), .S(n1701), .Y(n1450) );
  MUX2X1 U1430 ( .B(n1454), .A(n1455), .S(n1701), .Y(n1453) );
  MUX2X1 U1431 ( .B(n1457), .A(n1458), .S(n1686), .Y(n1456) );
  MUX2X1 U1432 ( .B(n1460), .A(n1461), .S(n1701), .Y(n1459) );
  MUX2X1 U1433 ( .B(n1463), .A(n1464), .S(n1701), .Y(n1462) );
  MUX2X1 U1434 ( .B(n1466), .A(n1467), .S(n1701), .Y(n1465) );
  MUX2X1 U1435 ( .B(n1469), .A(n1470), .S(n1701), .Y(n1468) );
  MUX2X1 U1436 ( .B(n1472), .A(n1473), .S(n1686), .Y(n1471) );
  MUX2X1 U1437 ( .B(n1475), .A(n1476), .S(n1701), .Y(n1474) );
  MUX2X1 U1438 ( .B(n1478), .A(n1479), .S(n1701), .Y(n1477) );
  MUX2X1 U1439 ( .B(n1481), .A(n1482), .S(n1701), .Y(n1480) );
  MUX2X1 U1440 ( .B(n1484), .A(n1485), .S(n1701), .Y(n1483) );
  MUX2X1 U1441 ( .B(n1487), .A(n1488), .S(n1686), .Y(n1486) );
  MUX2X1 U1442 ( .B(n1490), .A(n1491), .S(n1702), .Y(n1489) );
  MUX2X1 U1443 ( .B(n1493), .A(n1494), .S(n1702), .Y(n1492) );
  MUX2X1 U1444 ( .B(n1496), .A(n1497), .S(n1702), .Y(n1495) );
  MUX2X1 U1445 ( .B(n1499), .A(n1500), .S(n1702), .Y(n1498) );
  MUX2X1 U1446 ( .B(n1502), .A(n1503), .S(n1686), .Y(n1501) );
  MUX2X1 U1447 ( .B(n1505), .A(n1506), .S(n1702), .Y(n1504) );
  MUX2X1 U1448 ( .B(n1508), .A(n1509), .S(n1702), .Y(n1507) );
  MUX2X1 U1449 ( .B(n1511), .A(n1512), .S(n1702), .Y(n1510) );
  MUX2X1 U1450 ( .B(n1514), .A(n1515), .S(n1702), .Y(n1513) );
  MUX2X1 U1451 ( .B(n1517), .A(n1518), .S(n1686), .Y(n1516) );
  MUX2X1 U1452 ( .B(n1520), .A(n1521), .S(n1702), .Y(n1519) );
  MUX2X1 U1453 ( .B(n1523), .A(n1524), .S(n1702), .Y(n1522) );
  MUX2X1 U1454 ( .B(n1526), .A(n1527), .S(n1702), .Y(n1525) );
  MUX2X1 U1455 ( .B(n1529), .A(n1530), .S(n1702), .Y(n1528) );
  MUX2X1 U1456 ( .B(n1532), .A(n1533), .S(n1686), .Y(n1531) );
  MUX2X1 U1457 ( .B(n1535), .A(n1536), .S(n1703), .Y(n1534) );
  MUX2X1 U1458 ( .B(n1538), .A(n1539), .S(n1703), .Y(n1537) );
  MUX2X1 U1459 ( .B(n1541), .A(n1542), .S(n1703), .Y(n1540) );
  MUX2X1 U1460 ( .B(n1544), .A(n1545), .S(n1703), .Y(n1543) );
  MUX2X1 U1461 ( .B(n1547), .A(n1548), .S(n1686), .Y(n1546) );
  MUX2X1 U1462 ( .B(n1550), .A(n1551), .S(n1703), .Y(n1549) );
  MUX2X1 U1463 ( .B(n1553), .A(n1554), .S(n1703), .Y(n1552) );
  MUX2X1 U1464 ( .B(n1556), .A(n1557), .S(n1703), .Y(n1555) );
  MUX2X1 U1465 ( .B(n1559), .A(n1560), .S(n1703), .Y(n1558) );
  MUX2X1 U1466 ( .B(n1562), .A(n1563), .S(n1686), .Y(n1561) );
  MUX2X1 U1467 ( .B(n1565), .A(n1566), .S(n1703), .Y(n1564) );
  MUX2X1 U1468 ( .B(n1568), .A(n1569), .S(n1703), .Y(n1567) );
  MUX2X1 U1469 ( .B(n1571), .A(n1572), .S(n1703), .Y(n1570) );
  MUX2X1 U1470 ( .B(n1574), .A(n1575), .S(n1703), .Y(n1573) );
  MUX2X1 U1471 ( .B(n1577), .A(n1578), .S(n1687), .Y(n1576) );
  MUX2X1 U1472 ( .B(n1580), .A(n1581), .S(n1704), .Y(n1579) );
  MUX2X1 U1473 ( .B(n1583), .A(n1584), .S(n1704), .Y(n1582) );
  MUX2X1 U1474 ( .B(n1586), .A(n1587), .S(n1704), .Y(n1585) );
  MUX2X1 U1475 ( .B(n1589), .A(n1590), .S(n1704), .Y(n1588) );
  MUX2X1 U1476 ( .B(n1592), .A(n1593), .S(n1686), .Y(n1591) );
  MUX2X1 U1477 ( .B(n1595), .A(n1596), .S(n1704), .Y(n1594) );
  MUX2X1 U1478 ( .B(n1598), .A(n1599), .S(n1704), .Y(n1597) );
  MUX2X1 U1479 ( .B(n1601), .A(n1602), .S(n1704), .Y(n1600) );
  MUX2X1 U1480 ( .B(n1604), .A(n1605), .S(n1704), .Y(n1603) );
  MUX2X1 U1481 ( .B(n1607), .A(n1608), .S(n1686), .Y(n1606) );
  MUX2X1 U1482 ( .B(n1610), .A(n1611), .S(n1704), .Y(n1609) );
  MUX2X1 U1483 ( .B(n1613), .A(n1614), .S(n1704), .Y(n1612) );
  MUX2X1 U1484 ( .B(n1616), .A(n1617), .S(n1704), .Y(n1615) );
  MUX2X1 U1485 ( .B(n1619), .A(n1620), .S(n1704), .Y(n1618) );
  MUX2X1 U1486 ( .B(n1622), .A(n1623), .S(n1687), .Y(n1621) );
  MUX2X1 U1487 ( .B(n1625), .A(n1626), .S(n1705), .Y(n1624) );
  MUX2X1 U1488 ( .B(n1628), .A(n1629), .S(n1705), .Y(n1627) );
  MUX2X1 U1489 ( .B(n1631), .A(n1632), .S(n1705), .Y(n1630) );
  MUX2X1 U1490 ( .B(n1634), .A(n1635), .S(n1705), .Y(n1633) );
  MUX2X1 U1491 ( .B(n1637), .A(n1638), .S(n1686), .Y(n1636) );
  MUX2X1 U1492 ( .B(n1640), .A(n1641), .S(n1705), .Y(n1639) );
  MUX2X1 U1493 ( .B(n1643), .A(n1644), .S(n1705), .Y(n1642) );
  MUX2X1 U1494 ( .B(n1646), .A(n1647), .S(n1705), .Y(n1645) );
  MUX2X1 U1495 ( .B(n1649), .A(n1650), .S(n1705), .Y(n1648) );
  MUX2X1 U1496 ( .B(n1652), .A(n1653), .S(n1687), .Y(n1651) );
  MUX2X1 U1497 ( .B(n1655), .A(n1656), .S(n1705), .Y(n1654) );
  MUX2X1 U1498 ( .B(n1658), .A(n1659), .S(n1705), .Y(n1657) );
  MUX2X1 U1499 ( .B(n1661), .A(n1662), .S(n1705), .Y(n1660) );
  MUX2X1 U1500 ( .B(n1664), .A(n1665), .S(n1705), .Y(n1663) );
  MUX2X1 U1501 ( .B(n1667), .A(n1668), .S(n1687), .Y(n1666) );
  MUX2X1 U1502 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1711), .Y(n1191) );
  MUX2X1 U1503 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1714), .Y(n1190) );
  MUX2X1 U1504 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1716), .Y(n1194) );
  MUX2X1 U1505 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1722), .Y(n1193) );
  MUX2X1 U1506 ( .B(n1192), .A(n1189), .S(n1693), .Y(n1203) );
  MUX2X1 U1507 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1713), .Y(n1197) );
  MUX2X1 U1508 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1709), .Y(n1196) );
  MUX2X1 U1509 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1715), .Y(n1200) );
  MUX2X1 U1510 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1721), .Y(n1199) );
  MUX2X1 U1511 ( .B(n1198), .A(n1195), .S(n1693), .Y(n1202) );
  MUX2X1 U1512 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1723), .Y(n1206) );
  MUX2X1 U1513 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1717), .Y(n1205) );
  MUX2X1 U1514 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1722), .Y(n1209) );
  MUX2X1 U1515 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1721), .Y(n1208) );
  MUX2X1 U1516 ( .B(n1207), .A(n1204), .S(n1693), .Y(n1218) );
  MUX2X1 U1517 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1716), .Y(n1212) );
  MUX2X1 U1518 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1724), .Y(n1211) );
  MUX2X1 U1519 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1723), .Y(n1215) );
  MUX2X1 U1520 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1717), .Y(n1214) );
  MUX2X1 U1521 ( .B(n1213), .A(n1210), .S(n1693), .Y(n1217) );
  MUX2X1 U1522 ( .B(n1216), .A(n1201), .S(n1685), .Y(n1669) );
  MUX2X1 U1523 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1721), .Y(n1221) );
  MUX2X1 U1524 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1709), .Y(n1220) );
  MUX2X1 U1525 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1716), .Y(n1224) );
  MUX2X1 U1526 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1720), .Y(n1223) );
  MUX2X1 U1527 ( .B(n1222), .A(n1219), .S(n1693), .Y(n1233) );
  MUX2X1 U1528 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1723), .Y(n1227) );
  MUX2X1 U1529 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1720), .Y(n1226) );
  MUX2X1 U1530 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1722), .Y(n1230) );
  MUX2X1 U1531 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1709), .Y(n1229) );
  MUX2X1 U1532 ( .B(n1228), .A(n1225), .S(n1693), .Y(n1232) );
  MUX2X1 U1533 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1709), .Y(n1236) );
  MUX2X1 U1534 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1715), .Y(n1235) );
  MUX2X1 U1535 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1709), .Y(n1239) );
  MUX2X1 U1536 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1709), .Y(n1238) );
  MUX2X1 U1537 ( .B(n1237), .A(n1234), .S(n1693), .Y(n1248) );
  MUX2X1 U1538 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1709), .Y(n1242) );
  MUX2X1 U1539 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1709), .Y(n1241) );
  MUX2X1 U1540 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1709), .Y(n1245) );
  MUX2X1 U1541 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1709), .Y(n1244) );
  MUX2X1 U1542 ( .B(n1243), .A(n1240), .S(n1693), .Y(n1247) );
  MUX2X1 U1543 ( .B(n1246), .A(n1231), .S(n1685), .Y(n1670) );
  MUX2X1 U1544 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1709), .Y(n1251) );
  MUX2X1 U1545 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1709), .Y(n1250) );
  MUX2X1 U1546 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1709), .Y(n1254) );
  MUX2X1 U1547 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1709), .Y(n1253) );
  MUX2X1 U1548 ( .B(n1252), .A(n1249), .S(n1693), .Y(n1263) );
  MUX2X1 U1549 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1709), .Y(n1257) );
  MUX2X1 U1550 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1709), .Y(n1256) );
  MUX2X1 U1551 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1709), .Y(n1260) );
  MUX2X1 U1552 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1709), .Y(n1259) );
  MUX2X1 U1553 ( .B(n1258), .A(n1255), .S(n1693), .Y(n1262) );
  MUX2X1 U1554 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1710), .Y(n1266) );
  MUX2X1 U1555 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1710), .Y(n1265) );
  MUX2X1 U1556 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1710), .Y(n1269) );
  MUX2X1 U1557 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1710), .Y(n1268) );
  MUX2X1 U1558 ( .B(n1267), .A(n1264), .S(n1693), .Y(n1278) );
  MUX2X1 U1559 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1710), .Y(n1272) );
  MUX2X1 U1560 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1710), .Y(n1271) );
  MUX2X1 U1561 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1710), .Y(n1275) );
  MUX2X1 U1562 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1710), .Y(n1274) );
  MUX2X1 U1563 ( .B(n1273), .A(n1270), .S(n1693), .Y(n1277) );
  MUX2X1 U1564 ( .B(n1276), .A(n1261), .S(n1685), .Y(n1671) );
  MUX2X1 U1565 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1710), .Y(n1281) );
  MUX2X1 U1566 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1710), .Y(n1280) );
  MUX2X1 U1567 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1710), .Y(n1284) );
  MUX2X1 U1568 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1710), .Y(n1283) );
  MUX2X1 U1569 ( .B(n1282), .A(n1279), .S(n1692), .Y(n1293) );
  MUX2X1 U1570 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1711), .Y(n1287) );
  MUX2X1 U1571 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1711), .Y(n1286) );
  MUX2X1 U1572 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1711), .Y(n1290) );
  MUX2X1 U1573 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1711), .Y(n1289) );
  MUX2X1 U1574 ( .B(n1288), .A(n1285), .S(n1692), .Y(n1292) );
  MUX2X1 U1575 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1711), .Y(n1296) );
  MUX2X1 U1576 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1711), .Y(n1295) );
  MUX2X1 U1577 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1711), .Y(n1299) );
  MUX2X1 U1578 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1711), .Y(n1298) );
  MUX2X1 U1579 ( .B(n1297), .A(n1294), .S(n1692), .Y(n1308) );
  MUX2X1 U1580 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1711), .Y(n1302) );
  MUX2X1 U1581 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1711), .Y(n1301) );
  MUX2X1 U1582 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1711), .Y(n1305) );
  MUX2X1 U1583 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1711), .Y(n1304) );
  MUX2X1 U1584 ( .B(n1303), .A(n1300), .S(n1692), .Y(n1307) );
  MUX2X1 U1585 ( .B(n1306), .A(n1291), .S(n1685), .Y(n1672) );
  MUX2X1 U1586 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1712), .Y(n1311) );
  MUX2X1 U1587 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1712), .Y(n1310) );
  MUX2X1 U1588 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1712), .Y(n1314) );
  MUX2X1 U1589 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1712), .Y(n1313) );
  MUX2X1 U1590 ( .B(n1312), .A(n1309), .S(n1692), .Y(n1323) );
  MUX2X1 U1591 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1712), .Y(n1317) );
  MUX2X1 U1592 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1712), .Y(n1316) );
  MUX2X1 U1593 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1712), .Y(n1320) );
  MUX2X1 U1594 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1712), .Y(n1319) );
  MUX2X1 U1595 ( .B(n1318), .A(n1315), .S(n1692), .Y(n1322) );
  MUX2X1 U1596 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1712), .Y(n1326) );
  MUX2X1 U1597 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1712), .Y(n1325) );
  MUX2X1 U1598 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1712), .Y(n1329) );
  MUX2X1 U1599 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1712), .Y(n1328) );
  MUX2X1 U1600 ( .B(n1327), .A(n1324), .S(n1692), .Y(n1338) );
  MUX2X1 U1601 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1713), .Y(n1332) );
  MUX2X1 U1602 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1713), .Y(n1331) );
  MUX2X1 U1603 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1713), .Y(n1335) );
  MUX2X1 U1604 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1713), .Y(n1334) );
  MUX2X1 U1605 ( .B(n1333), .A(n1330), .S(n1692), .Y(n1337) );
  MUX2X1 U1606 ( .B(n1336), .A(n1321), .S(n1685), .Y(n1673) );
  MUX2X1 U1607 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1713), .Y(n1341) );
  MUX2X1 U1608 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1713), .Y(n1340) );
  MUX2X1 U1609 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1713), .Y(n1344) );
  MUX2X1 U1610 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1713), .Y(n1343) );
  MUX2X1 U1611 ( .B(n1342), .A(n1339), .S(n1692), .Y(n1353) );
  MUX2X1 U1612 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1713), .Y(n1347) );
  MUX2X1 U1613 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1713), .Y(n1346) );
  MUX2X1 U1614 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1713), .Y(n1350) );
  MUX2X1 U1615 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1713), .Y(n1349) );
  MUX2X1 U1616 ( .B(n1348), .A(n1345), .S(n1692), .Y(n1352) );
  MUX2X1 U1617 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1714), .Y(n1356) );
  MUX2X1 U1618 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1714), .Y(n1355) );
  MUX2X1 U1619 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1714), .Y(n1359) );
  MUX2X1 U1620 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1714), .Y(n1358) );
  MUX2X1 U1621 ( .B(n1357), .A(n1354), .S(n1692), .Y(n1368) );
  MUX2X1 U1622 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1714), .Y(n1362) );
  MUX2X1 U1623 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1714), .Y(n1361) );
  MUX2X1 U1624 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1714), .Y(n1365) );
  MUX2X1 U1625 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1714), .Y(n1364) );
  MUX2X1 U1626 ( .B(n1363), .A(n1360), .S(n1692), .Y(n1367) );
  MUX2X1 U1627 ( .B(n1366), .A(n1351), .S(n1685), .Y(n1674) );
  MUX2X1 U1628 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1714), .Y(n1371) );
  MUX2X1 U1629 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1714), .Y(n1370) );
  MUX2X1 U1630 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1714), .Y(n1374) );
  MUX2X1 U1631 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1714), .Y(n1373) );
  MUX2X1 U1632 ( .B(n1372), .A(n1369), .S(n1691), .Y(n1383) );
  MUX2X1 U1633 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1715), .Y(n1377) );
  MUX2X1 U1634 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1715), .Y(n1376) );
  MUX2X1 U1635 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1715), .Y(n1380) );
  MUX2X1 U1636 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1715), .Y(n1379) );
  MUX2X1 U1637 ( .B(n1378), .A(n1375), .S(n1691), .Y(n1382) );
  MUX2X1 U1638 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1715), .Y(n1386) );
  MUX2X1 U1639 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1715), .Y(n1385) );
  MUX2X1 U1640 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1715), .Y(n1389) );
  MUX2X1 U1641 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1715), .Y(n1388) );
  MUX2X1 U1642 ( .B(n1387), .A(n1384), .S(n1691), .Y(n1398) );
  MUX2X1 U1643 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1715), .Y(n1392) );
  MUX2X1 U1644 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1715), .Y(n1391) );
  MUX2X1 U1645 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1715), .Y(n1395) );
  MUX2X1 U1646 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1715), .Y(n1394) );
  MUX2X1 U1647 ( .B(n1393), .A(n1390), .S(n1691), .Y(n1397) );
  MUX2X1 U1648 ( .B(n1396), .A(n1381), .S(n1685), .Y(n1675) );
  MUX2X1 U1649 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1716), .Y(n1401) );
  MUX2X1 U1650 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1716), .Y(n1400) );
  MUX2X1 U1651 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1716), .Y(n1404) );
  MUX2X1 U1652 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1716), .Y(n1403) );
  MUX2X1 U1653 ( .B(n1402), .A(n1399), .S(n1691), .Y(n1413) );
  MUX2X1 U1654 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1716), .Y(n1407) );
  MUX2X1 U1655 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1716), .Y(n1406) );
  MUX2X1 U1656 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1716), .Y(n1410) );
  MUX2X1 U1657 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1716), .Y(n1409) );
  MUX2X1 U1658 ( .B(n1408), .A(n1405), .S(n1691), .Y(n1412) );
  MUX2X1 U1659 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1716), .Y(n1416) );
  MUX2X1 U1660 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1716), .Y(n1415) );
  MUX2X1 U1661 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1716), .Y(n1419) );
  MUX2X1 U1662 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1716), .Y(n1418) );
  MUX2X1 U1663 ( .B(n1417), .A(n1414), .S(n1691), .Y(n1428) );
  MUX2X1 U1664 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1717), .Y(n1422) );
  MUX2X1 U1665 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1717), .Y(n1421) );
  MUX2X1 U1666 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1717), .Y(n1425) );
  MUX2X1 U1667 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1717), .Y(n1424) );
  MUX2X1 U1668 ( .B(n1423), .A(n1420), .S(n1691), .Y(n1427) );
  MUX2X1 U1669 ( .B(n1426), .A(n1411), .S(n1685), .Y(n1676) );
  MUX2X1 U1670 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1717), .Y(n1431) );
  MUX2X1 U1671 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1717), .Y(n1430) );
  MUX2X1 U1672 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1717), .Y(n1434) );
  MUX2X1 U1673 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1717), .Y(n1433) );
  MUX2X1 U1674 ( .B(n1432), .A(n1429), .S(n1691), .Y(n1443) );
  MUX2X1 U1675 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1717), .Y(n1437) );
  MUX2X1 U1676 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1717), .Y(n1436) );
  MUX2X1 U1677 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1717), .Y(n1440) );
  MUX2X1 U1678 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1717), .Y(n1439) );
  MUX2X1 U1679 ( .B(n1438), .A(n1435), .S(n1691), .Y(n1442) );
  MUX2X1 U1680 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1718), .Y(n1446) );
  MUX2X1 U1681 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1718), .Y(n1445) );
  MUX2X1 U1682 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1718), .Y(n1449) );
  MUX2X1 U1683 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1718), .Y(n1448) );
  MUX2X1 U1684 ( .B(n1447), .A(n1444), .S(n1691), .Y(n1458) );
  MUX2X1 U1685 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1718), .Y(n1452) );
  MUX2X1 U1686 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1718), .Y(n1451) );
  MUX2X1 U1687 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1718), .Y(n1455) );
  MUX2X1 U1688 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1718), .Y(n1454) );
  MUX2X1 U1689 ( .B(n1453), .A(n1450), .S(n1691), .Y(n1457) );
  MUX2X1 U1690 ( .B(n1456), .A(n1441), .S(n1685), .Y(n1677) );
  MUX2X1 U1691 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1718), .Y(n1461) );
  MUX2X1 U1692 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1718), .Y(n1460) );
  MUX2X1 U1693 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1718), .Y(n1464) );
  MUX2X1 U1694 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1718), .Y(n1463) );
  MUX2X1 U1695 ( .B(n1462), .A(n1459), .S(n1690), .Y(n1473) );
  MUX2X1 U1696 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1718), .Y(n1467) );
  MUX2X1 U1697 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1719), .Y(n1466) );
  MUX2X1 U1698 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1715), .Y(n1470) );
  MUX2X1 U1699 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1715), .Y(n1469) );
  MUX2X1 U1700 ( .B(n1468), .A(n1465), .S(n1690), .Y(n1472) );
  MUX2X1 U1701 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1717), .Y(n1476) );
  MUX2X1 U1702 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1716), .Y(n1475) );
  MUX2X1 U1703 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1715), .Y(n1479) );
  MUX2X1 U1704 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1718), .Y(n1478) );
  MUX2X1 U1705 ( .B(n1477), .A(n1474), .S(n1690), .Y(n1488) );
  MUX2X1 U1706 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1716), .Y(n1482) );
  MUX2X1 U1707 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1720), .Y(n1481) );
  MUX2X1 U1708 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1717), .Y(n1485) );
  MUX2X1 U1709 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1719), .Y(n1484) );
  MUX2X1 U1710 ( .B(n1483), .A(n1480), .S(n1690), .Y(n1487) );
  MUX2X1 U1711 ( .B(n1486), .A(n1471), .S(n1685), .Y(n1678) );
  MUX2X1 U1712 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1719), .Y(n1491) );
  MUX2X1 U1713 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1719), .Y(n1490) );
  MUX2X1 U1714 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1719), .Y(n1494) );
  MUX2X1 U1715 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1719), .Y(n1493) );
  MUX2X1 U1716 ( .B(n1492), .A(n1489), .S(n1690), .Y(n1503) );
  MUX2X1 U1717 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1719), .Y(n1497) );
  MUX2X1 U1718 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1719), .Y(n1496) );
  MUX2X1 U1719 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1719), .Y(n1500) );
  MUX2X1 U1720 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1719), .Y(n1499) );
  MUX2X1 U1721 ( .B(n1498), .A(n1495), .S(n1690), .Y(n1502) );
  MUX2X1 U1722 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1719), .Y(n1506) );
  MUX2X1 U1723 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1719), .Y(n1505) );
  MUX2X1 U1724 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1719), .Y(n1509) );
  MUX2X1 U1725 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1719), .Y(n1508) );
  MUX2X1 U1726 ( .B(n1507), .A(n1504), .S(n1690), .Y(n1518) );
  MUX2X1 U1727 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1720), .Y(n1512) );
  MUX2X1 U1728 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1720), .Y(n1511) );
  MUX2X1 U1729 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1720), .Y(n1515) );
  MUX2X1 U1730 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1720), .Y(n1514) );
  MUX2X1 U1731 ( .B(n1513), .A(n1510), .S(n1690), .Y(n1517) );
  MUX2X1 U1732 ( .B(n1516), .A(n1501), .S(n1685), .Y(n1679) );
  MUX2X1 U1733 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1720), .Y(n1521) );
  MUX2X1 U1734 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1720), .Y(n1520) );
  MUX2X1 U1735 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1720), .Y(n1524) );
  MUX2X1 U1736 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1720), .Y(n1523) );
  MUX2X1 U1737 ( .B(n1522), .A(n1519), .S(n1690), .Y(n1533) );
  MUX2X1 U1738 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1720), .Y(n1527) );
  MUX2X1 U1739 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1720), .Y(n1526) );
  MUX2X1 U1740 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1720), .Y(n1530) );
  MUX2X1 U1741 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1720), .Y(n1529) );
  MUX2X1 U1742 ( .B(n1528), .A(n1525), .S(n1690), .Y(n1532) );
  MUX2X1 U1743 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1721), .Y(n1536) );
  MUX2X1 U1744 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1715), .Y(n1535) );
  MUX2X1 U1745 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1716), .Y(n1539) );
  MUX2X1 U1746 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1722), .Y(n1538) );
  MUX2X1 U1747 ( .B(n1537), .A(n1534), .S(n1690), .Y(n1548) );
  MUX2X1 U1748 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1722), .Y(n1542) );
  MUX2X1 U1749 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1723), .Y(n1541) );
  MUX2X1 U1750 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1717), .Y(n1545) );
  MUX2X1 U1751 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1717), .Y(n1544) );
  MUX2X1 U1752 ( .B(n1543), .A(n1540), .S(n1690), .Y(n1547) );
  MUX2X1 U1753 ( .B(n1546), .A(n1531), .S(n1685), .Y(n1680) );
  MUX2X1 U1754 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1717), .Y(n1551) );
  MUX2X1 U1755 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1721), .Y(n1550) );
  MUX2X1 U1756 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1715), .Y(n1554) );
  MUX2X1 U1757 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1723), .Y(n1553) );
  MUX2X1 U1758 ( .B(n1552), .A(n1549), .S(n1689), .Y(n1563) );
  MUX2X1 U1759 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1710), .Y(n1557) );
  MUX2X1 U1760 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1711), .Y(n1556) );
  MUX2X1 U1761 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1711), .Y(n1560) );
  MUX2X1 U1762 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1710), .Y(n1559) );
  MUX2X1 U1763 ( .B(n1558), .A(n1555), .S(n1689), .Y(n1562) );
  MUX2X1 U1764 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1710), .Y(n1566) );
  MUX2X1 U1765 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1711), .Y(n1565) );
  MUX2X1 U1766 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1711), .Y(n1569) );
  MUX2X1 U1767 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1710), .Y(n1568) );
  MUX2X1 U1768 ( .B(n1567), .A(n1564), .S(n1689), .Y(n1578) );
  MUX2X1 U1769 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1710), .Y(n1572) );
  MUX2X1 U1770 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1711), .Y(n1571) );
  MUX2X1 U1771 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1710), .Y(n1575) );
  MUX2X1 U1772 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1710), .Y(n1574) );
  MUX2X1 U1773 ( .B(n1573), .A(n1570), .S(n1689), .Y(n1577) );
  MUX2X1 U1774 ( .B(n1576), .A(n1561), .S(n1685), .Y(n1681) );
  MUX2X1 U1775 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1721), .Y(n1581) );
  MUX2X1 U1776 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1721), .Y(n1580) );
  MUX2X1 U1777 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1721), .Y(n1584) );
  MUX2X1 U1778 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1721), .Y(n1583) );
  MUX2X1 U1779 ( .B(n1582), .A(n1579), .S(n1689), .Y(n1593) );
  MUX2X1 U1780 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1721), .Y(n1587) );
  MUX2X1 U1781 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1721), .Y(n1586) );
  MUX2X1 U1782 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1721), .Y(n1590) );
  MUX2X1 U1783 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1721), .Y(n1589) );
  MUX2X1 U1784 ( .B(n1588), .A(n1585), .S(n1689), .Y(n1592) );
  MUX2X1 U1785 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1721), .Y(n1596) );
  MUX2X1 U1786 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1721), .Y(n1595) );
  MUX2X1 U1787 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1721), .Y(n1599) );
  MUX2X1 U1788 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1721), .Y(n1598) );
  MUX2X1 U1789 ( .B(n1597), .A(n1594), .S(n1689), .Y(n1608) );
  MUX2X1 U1790 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1722), .Y(n1602) );
  MUX2X1 U1791 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1722), .Y(n1601) );
  MUX2X1 U1792 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1722), .Y(n1605) );
  MUX2X1 U1793 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1722), .Y(n1604) );
  MUX2X1 U1794 ( .B(n1603), .A(n1600), .S(n1689), .Y(n1607) );
  MUX2X1 U1795 ( .B(n1606), .A(n1591), .S(n1685), .Y(n1682) );
  MUX2X1 U1796 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1722), .Y(n1611) );
  MUX2X1 U1797 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1722), .Y(n1610) );
  MUX2X1 U1798 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1722), .Y(n1614) );
  MUX2X1 U1799 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1722), .Y(n1613) );
  MUX2X1 U1800 ( .B(n1612), .A(n1609), .S(n1689), .Y(n1623) );
  MUX2X1 U1801 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1722), .Y(n1617) );
  MUX2X1 U1802 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1722), .Y(n1616) );
  MUX2X1 U1803 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1722), .Y(n1620) );
  MUX2X1 U1804 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1722), .Y(n1619) );
  MUX2X1 U1805 ( .B(n1618), .A(n1615), .S(n1689), .Y(n1622) );
  MUX2X1 U1806 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1723), .Y(n1626) );
  MUX2X1 U1807 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1723), .Y(n1625) );
  MUX2X1 U1808 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1723), .Y(n1629) );
  MUX2X1 U1809 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1723), .Y(n1628) );
  MUX2X1 U1810 ( .B(n1627), .A(n1624), .S(n1689), .Y(n1638) );
  MUX2X1 U1811 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1723), .Y(n1632) );
  MUX2X1 U1812 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1723), .Y(n1631) );
  MUX2X1 U1813 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1723), .Y(n1635) );
  MUX2X1 U1814 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1723), .Y(n1634) );
  MUX2X1 U1815 ( .B(n1633), .A(n1630), .S(n1689), .Y(n1637) );
  MUX2X1 U1816 ( .B(n1636), .A(n1621), .S(n1685), .Y(n1683) );
  MUX2X1 U1817 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1723), .Y(n1641) );
  MUX2X1 U1818 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1723), .Y(n1640) );
  MUX2X1 U1819 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1723), .Y(n1644) );
  MUX2X1 U1820 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1723), .Y(n1643) );
  MUX2X1 U1821 ( .B(n1642), .A(n1639), .S(n1688), .Y(n1653) );
  MUX2X1 U1822 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1714), .Y(n1647) );
  MUX2X1 U1823 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1709), .Y(n1646) );
  MUX2X1 U1824 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1722), .Y(n1650) );
  MUX2X1 U1825 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1721), .Y(n1649) );
  MUX2X1 U1826 ( .B(n1648), .A(n1645), .S(n1688), .Y(n1652) );
  MUX2X1 U1827 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1716), .Y(n1656) );
  MUX2X1 U1828 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1717), .Y(n1655) );
  MUX2X1 U1829 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1722), .Y(n1659) );
  MUX2X1 U1830 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1723), .Y(n1658) );
  MUX2X1 U1831 ( .B(n1657), .A(n1654), .S(n1688), .Y(n1668) );
  MUX2X1 U1832 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1723), .Y(n1662) );
  MUX2X1 U1833 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1724), .Y(n1661) );
  MUX2X1 U1834 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1716), .Y(n1665) );
  MUX2X1 U1835 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1721), .Y(n1664) );
  MUX2X1 U1836 ( .B(n1663), .A(n1660), .S(n1688), .Y(n1667) );
  MUX2X1 U1837 ( .B(n1666), .A(n1651), .S(n1685), .Y(n1684) );
  INVX8 U1838 ( .A(n1845), .Y(n1689) );
  INVX8 U1839 ( .A(n1707), .Y(n1712) );
  INVX8 U1840 ( .A(n1707), .Y(n1713) );
  INVX8 U1841 ( .A(n1707), .Y(n1714) );
  INVX1 U1842 ( .A(N11), .Y(n1844) );
  INVX1 U1843 ( .A(N10), .Y(n1842) );
  INVX8 U1844 ( .A(n1824), .Y(n1821) );
  INVX8 U1845 ( .A(n1824), .Y(n1822) );
  INVX8 U1846 ( .A(n1824), .Y(n1823) );
  INVX8 U1847 ( .A(n2877), .Y(n1824) );
  INVX8 U1848 ( .A(n39), .Y(n1825) );
  INVX8 U1849 ( .A(n42), .Y(n1827) );
  INVX8 U1850 ( .A(n44), .Y(n1829) );
  INVX8 U1851 ( .A(n47), .Y(n1831) );
  INVX8 U1852 ( .A(n50), .Y(n1833) );
  INVX8 U1853 ( .A(n54), .Y(n1835) );
  INVX8 U1854 ( .A(n58), .Y(n1837) );
  INVX8 U1855 ( .A(n62), .Y(n1839) );
  OR2X2 U1856 ( .A(write), .B(rst), .Y(n1851) );
endmodule


module memc_Size16_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1847), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1848), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1849), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1850), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1851), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1852), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1853), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1854), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1855), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1856), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1857), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1858), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1859), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1860), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1861), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1862), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1863), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1864), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1865), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1866), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1867), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1868), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1869), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1870), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1871), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1872), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1873), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1874), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1875), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1876), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1877), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1878), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1879), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1880), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1881), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1882), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1883), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1884), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1885), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1886), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1887), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1888), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1889), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1890), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1891), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1892), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1893), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1894), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1895), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1896), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1897), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1898), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1899), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1900), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1901), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1902), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1903), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1904), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1905), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1906), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1907), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1908), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1909), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1910), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1911), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1912), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1913), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1914), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1915), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1916), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1917), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1918), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1919), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1920), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1921), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1922), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1923), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1924), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1925), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1926), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1927), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1928), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1929), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1930), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1931), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1932), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1933), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1934), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1935), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1936), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1937), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1938), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1939), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1940), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1941), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1942), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1943), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1944), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1945), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1946), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1947), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1948), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1949), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1950), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1951), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1952), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1953), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1954), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1955), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1956), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1957), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1958), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1959), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1960), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1961), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1962), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1963), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1964), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1965), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1966), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1967), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1968), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1969), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1970), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1971), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1972), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1973), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1974), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1975), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1976), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1977), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1978), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1979), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1980), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1981), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1982), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1983), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1984), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1985), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1986), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1987), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1988), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1989), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1990), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1991), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1992), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1993), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1994), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1995), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1996), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1997), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1998), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1999), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2000), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2001), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2002), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2003), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2004), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2005), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2006), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2007), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2008), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2009), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2010), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2011), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2012), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2013), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2014), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2015), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2016), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2017), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2018), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2019), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2020), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2021), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2022), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2023), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2024), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2025), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2026), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2027), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2028), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2029), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2030), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2031), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2032), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2033), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2034), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2035), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2036), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2037), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2038), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2039), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2040), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2041), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2042), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2043), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2044), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2045), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2046), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2047), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2048), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2049), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2050), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2051), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2052), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2053), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2054), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2055), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2056), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2057), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2058), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2059), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2060), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2061), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2062), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2063), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2064), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2065), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2066), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2067), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2068), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2069), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2070), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2071), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2072), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2073), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2074), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2075), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2076), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2077), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2078), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2079), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2080), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2081), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2082), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2083), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2084), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2085), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2086), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2087), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2088), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2089), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2090), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2091), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2092), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2093), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2094), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2095), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2096), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2097), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2098), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2099), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2100), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2101), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2102), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2103), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2104), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2105), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2106), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2107), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2108), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2109), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2110), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2111), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2112), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2113), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2114), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2115), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2116), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2117), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2118), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2119), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2120), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2121), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2122), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2123), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2124), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2125), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2126), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2127), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2128), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2129), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2130), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2131), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2132), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2133), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2134), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2135), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2136), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2137), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2138), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2139), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2140), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2141), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2142), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2143), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2144), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2145), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2146), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2147), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2148), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2149), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2150), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2151), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2152), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2153), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2154), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2155), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2156), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2157), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2158), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2159), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2160), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2161), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2162), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2163), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2164), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2165), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2166), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2167), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2168), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2169), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2170), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2171), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2172), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2173), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2174), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2175), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2176), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2177), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2178), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2179), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2180), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2181), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2182), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2183), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2184), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2185), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2186), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2187), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2188), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2189), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2190), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2191), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2192), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2193), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2194), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2195), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2196), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2197), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2198), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2199), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2200), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2201), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2202), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2203), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2204), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2205), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2206), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2207), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2208), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2209), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2210), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2211), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2212), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2213), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2214), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2215), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2216), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2217), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2218), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2219), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2220), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2221), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2222), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2223), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2224), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2225), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2226), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2227), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2228), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2229), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2230), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2231), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2232), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2233), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2234), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2235), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2236), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2237), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2238), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2239), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2240), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2241), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2242), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2243), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2244), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2245), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2246), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2247), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2248), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2249), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2250), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2251), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2252), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2253), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2254), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2255), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2256), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2257), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2258), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2259), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2260), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2261), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2262), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2263), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2264), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2265), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2266), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2267), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2268), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2269), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2270), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2271), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2272), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2273), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2274), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2275), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2276), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2277), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2278), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2279), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2280), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2281), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2282), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2283), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2284), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2285), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2286), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2287), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2288), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2289), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2290), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2291), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2292), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2293), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2294), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2295), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2296), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2297), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2298), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2299), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2300), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2301), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2302), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2303), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2304), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2305), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2306), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2307), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2308), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2309), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2310), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2311), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2312), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2313), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2314), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2315), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2316), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2317), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2318), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2319), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2320), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2321), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2322), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2323), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2324), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2325), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2326), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2327), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2328), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2329), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2330), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2331), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2332), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2333), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2334), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2335), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2336), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2337), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2338), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2339), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2340), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2341), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2342), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2343), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2344), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2345), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2346), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2347), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2348), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2349), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2350), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2351), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2352), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2353), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2354), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2355), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2356), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2357), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2358), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2359) );
  INVX1 U2 ( .A(n1309), .Y(n1200) );
  INVX1 U3 ( .A(n1190), .Y(n1197) );
  INVX1 U4 ( .A(n1309), .Y(n1198) );
  INVX1 U5 ( .A(n1309), .Y(n1199) );
  INVX1 U6 ( .A(n1188), .Y(n1201) );
  INVX2 U7 ( .A(n1188), .Y(n1202) );
  INVX2 U8 ( .A(n1188), .Y(n1203) );
  INVX1 U9 ( .A(N10), .Y(n1188) );
  INVX1 U10 ( .A(n1207), .Y(n1190) );
  INVX1 U11 ( .A(n1314), .Y(n1168) );
  INVX1 U12 ( .A(n1314), .Y(n1170) );
  INVX1 U13 ( .A(n1314), .Y(n1169) );
  INVX1 U14 ( .A(n1309), .Y(n1207) );
  INVX1 U15 ( .A(n1190), .Y(n1191) );
  INVX1 U16 ( .A(n1176), .Y(n1177) );
  INVX1 U17 ( .A(n1176), .Y(n1178) );
  INVX2 U18 ( .A(n1207), .Y(n1189) );
  INVX1 U19 ( .A(n1175), .Y(n1180) );
  INVX1 U20 ( .A(n1175), .Y(n1181) );
  INVX1 U21 ( .A(n1176), .Y(n1185) );
  INVX1 U22 ( .A(n1175), .Y(n1186) );
  INVX1 U23 ( .A(n1176), .Y(n1179) );
  INVX1 U24 ( .A(n1175), .Y(n1182) );
  INVX1 U25 ( .A(n639), .Y(N32) );
  INVX1 U26 ( .A(n640), .Y(N31) );
  INVX1 U27 ( .A(n641), .Y(N30) );
  INVX1 U28 ( .A(n643), .Y(N28) );
  INVX1 U29 ( .A(n644), .Y(N27) );
  INVX1 U30 ( .A(n645), .Y(N26) );
  INVX1 U31 ( .A(n647), .Y(N24) );
  INVX1 U32 ( .A(n648), .Y(N23) );
  INVX1 U33 ( .A(n649), .Y(N22) );
  INVX1 U34 ( .A(n1163), .Y(N20) );
  INVX1 U35 ( .A(n1164), .Y(N19) );
  INVX1 U36 ( .A(n1165), .Y(N18) );
  INVX1 U37 ( .A(n1166), .Y(N17) );
  INVX1 U38 ( .A(n642), .Y(N29) );
  INVX1 U39 ( .A(n646), .Y(N25) );
  INVX1 U40 ( .A(n650), .Y(N21) );
  BUFX2 U41 ( .A(n41), .Y(n1209) );
  BUFX2 U42 ( .A(n39), .Y(n1208) );
  BUFX2 U43 ( .A(n41), .Y(n1210) );
  BUFX2 U44 ( .A(n45), .Y(n1211) );
  BUFX2 U45 ( .A(n45), .Y(n1212) );
  BUFX2 U46 ( .A(n49), .Y(n1214) );
  BUFX2 U47 ( .A(n47), .Y(n1213) );
  BUFX2 U48 ( .A(n49), .Y(n1215) );
  BUFX2 U49 ( .A(n53), .Y(n1217) );
  BUFX2 U50 ( .A(n51), .Y(n1216) );
  BUFX2 U51 ( .A(n53), .Y(n1218) );
  BUFX2 U52 ( .A(n57), .Y(n1219) );
  BUFX2 U53 ( .A(n57), .Y(n1220) );
  BUFX2 U54 ( .A(n61), .Y(n1221) );
  BUFX2 U55 ( .A(n61), .Y(n1222) );
  BUFX2 U56 ( .A(n65), .Y(n1223) );
  BUFX2 U57 ( .A(n65), .Y(n1224) );
  BUFX2 U58 ( .A(n67), .Y(n1225) );
  BUFX2 U59 ( .A(n67), .Y(n1226) );
  BUFX2 U60 ( .A(n71), .Y(n1229) );
  BUFX2 U61 ( .A(n69), .Y(n1227) );
  BUFX2 U62 ( .A(n71), .Y(n1230) );
  BUFX2 U63 ( .A(n75), .Y(n1231) );
  BUFX2 U64 ( .A(n75), .Y(n1232) );
  BUFX2 U65 ( .A(n79), .Y(n1234) );
  BUFX2 U66 ( .A(n77), .Y(n1233) );
  BUFX2 U67 ( .A(n79), .Y(n1235) );
  BUFX2 U68 ( .A(n83), .Y(n1237) );
  BUFX2 U69 ( .A(n81), .Y(n1236) );
  BUFX2 U70 ( .A(n83), .Y(n1238) );
  BUFX2 U71 ( .A(n87), .Y(n1239) );
  BUFX2 U72 ( .A(n87), .Y(n1240) );
  BUFX2 U73 ( .A(n91), .Y(n1241) );
  BUFX2 U74 ( .A(n91), .Y(n1242) );
  BUFX2 U75 ( .A(n95), .Y(n1243) );
  BUFX2 U76 ( .A(n95), .Y(n1244) );
  BUFX2 U77 ( .A(n97), .Y(n1246) );
  BUFX2 U78 ( .A(n97), .Y(n1247) );
  BUFX2 U79 ( .A(n101), .Y(n1250) );
  BUFX2 U80 ( .A(n99), .Y(n1248) );
  BUFX2 U81 ( .A(n101), .Y(n1251) );
  BUFX2 U82 ( .A(n105), .Y(n1252) );
  BUFX2 U83 ( .A(n105), .Y(n1253) );
  BUFX2 U84 ( .A(n109), .Y(n1255) );
  BUFX2 U85 ( .A(n107), .Y(n1254) );
  BUFX2 U86 ( .A(n109), .Y(n1256) );
  BUFX2 U87 ( .A(n113), .Y(n1258) );
  BUFX2 U88 ( .A(n111), .Y(n1257) );
  BUFX2 U89 ( .A(n113), .Y(n1259) );
  BUFX2 U90 ( .A(n117), .Y(n1260) );
  BUFX2 U91 ( .A(n117), .Y(n1261) );
  BUFX2 U92 ( .A(n121), .Y(n1262) );
  BUFX2 U93 ( .A(n121), .Y(n1263) );
  BUFX2 U94 ( .A(n125), .Y(n1264) );
  BUFX2 U95 ( .A(n125), .Y(n1265) );
  BUFX2 U96 ( .A(n127), .Y(n1266) );
  BUFX2 U97 ( .A(n127), .Y(n1267) );
  BUFX2 U98 ( .A(n131), .Y(n1270) );
  BUFX2 U99 ( .A(n129), .Y(n1268) );
  BUFX2 U100 ( .A(n131), .Y(n1271) );
  BUFX2 U101 ( .A(n135), .Y(n1272) );
  BUFX2 U102 ( .A(n135), .Y(n1273) );
  BUFX2 U103 ( .A(n139), .Y(n1275) );
  BUFX2 U104 ( .A(n137), .Y(n1274) );
  BUFX2 U105 ( .A(n139), .Y(n1276) );
  BUFX2 U106 ( .A(n143), .Y(n1278) );
  BUFX2 U107 ( .A(n141), .Y(n1277) );
  BUFX2 U108 ( .A(n143), .Y(n1279) );
  BUFX2 U109 ( .A(n147), .Y(n1280) );
  BUFX2 U110 ( .A(n147), .Y(n1281) );
  BUFX2 U111 ( .A(n151), .Y(n1282) );
  BUFX2 U112 ( .A(n151), .Y(n1283) );
  BUFX2 U113 ( .A(n155), .Y(n1284) );
  BUFX2 U114 ( .A(n155), .Y(n1285) );
  BUFX2 U115 ( .A(n157), .Y(n1286) );
  BUFX2 U116 ( .A(n157), .Y(n1287) );
  INVX2 U117 ( .A(n1187), .Y(n1183) );
  INVX1 U118 ( .A(n1187), .Y(n1184) );
  INVX2 U119 ( .A(n1171), .Y(n1172) );
  INVX2 U120 ( .A(n1188), .Y(n1204) );
  INVX2 U121 ( .A(n1190), .Y(n1206) );
  INVX1 U122 ( .A(n1312), .Y(n1173) );
  INVX1 U123 ( .A(n1312), .Y(n1174) );
  INVX1 U124 ( .A(n1310), .Y(n1187) );
  INVX1 U125 ( .A(N12), .Y(n1312) );
  INVX1 U126 ( .A(n1310), .Y(n1175) );
  INVX1 U127 ( .A(n1310), .Y(n1176) );
  INVX1 U128 ( .A(N13), .Y(n1314) );
  INVX1 U129 ( .A(N14), .Y(n1316) );
  INVX1 U130 ( .A(N12), .Y(n1171) );
  INVX1 U131 ( .A(n1316), .Y(n1167) );
  INVX1 U132 ( .A(rst), .Y(n1317) );
  BUFX2 U133 ( .A(n69), .Y(n1228) );
  BUFX2 U134 ( .A(n99), .Y(n1249) );
  BUFX2 U135 ( .A(n129), .Y(n1269) );
  INVX1 U136 ( .A(n33), .Y(n1245) );
  AND2X2 U137 ( .A(\data_in<11> ), .B(n1289), .Y(n1) );
  AND2X2 U138 ( .A(\data_in<12> ), .B(n1289), .Y(n2) );
  AND2X2 U139 ( .A(\data_in<13> ), .B(n1289), .Y(n3) );
  AND2X2 U140 ( .A(\data_in<14> ), .B(n1289), .Y(n4) );
  AND2X2 U141 ( .A(\data_in<15> ), .B(n1289), .Y(n5) );
  INVX1 U142 ( .A(n1309), .Y(n1308) );
  INVX1 U143 ( .A(n1314), .Y(n1313) );
  AND2X1 U144 ( .A(n1173), .B(n1310), .Y(n6) );
  INVX1 U145 ( .A(n1311), .Y(n1310) );
  AND2X1 U146 ( .A(n2359), .B(n1315), .Y(n7) );
  INVX1 U147 ( .A(n1316), .Y(n1315) );
  BUFX2 U148 ( .A(n1352), .Y(n8) );
  INVX1 U149 ( .A(n8), .Y(n1744) );
  BUFX2 U150 ( .A(n1369), .Y(n9) );
  INVX1 U151 ( .A(n9), .Y(n1761) );
  BUFX2 U152 ( .A(n1386), .Y(n10) );
  INVX1 U153 ( .A(n10), .Y(n1778) );
  BUFX2 U154 ( .A(n1403), .Y(n11) );
  INVX1 U155 ( .A(n11), .Y(n1795) );
  BUFX2 U156 ( .A(n1420), .Y(n12) );
  INVX1 U157 ( .A(n12), .Y(n1812) );
  BUFX2 U158 ( .A(n1581), .Y(n13) );
  INVX1 U159 ( .A(n13), .Y(n1694) );
  BUFX2 U160 ( .A(n1711), .Y(n14) );
  INVX1 U161 ( .A(n14), .Y(n1829) );
  AND2X1 U162 ( .A(n1308), .B(n6), .Y(n15) );
  AND2X1 U163 ( .A(n1313), .B(n7), .Y(n16) );
  AND2X2 U164 ( .A(write), .B(n1317), .Y(n17) );
  AND2X1 U165 ( .A(n1309), .B(n6), .Y(n18) );
  AND2X1 U166 ( .A(n1314), .B(n7), .Y(n19) );
  AND2X2 U167 ( .A(\data_in<0> ), .B(n1290), .Y(n20) );
  AND2X2 U168 ( .A(\data_in<1> ), .B(n1290), .Y(n21) );
  AND2X2 U169 ( .A(\data_in<2> ), .B(n1290), .Y(n22) );
  AND2X2 U170 ( .A(\data_in<3> ), .B(n1290), .Y(n23) );
  AND2X2 U171 ( .A(\data_in<4> ), .B(n1290), .Y(n24) );
  AND2X2 U172 ( .A(\data_in<5> ), .B(n1290), .Y(n25) );
  AND2X2 U173 ( .A(\data_in<6> ), .B(n1290), .Y(n26) );
  AND2X2 U174 ( .A(\data_in<7> ), .B(n1290), .Y(n27) );
  AND2X2 U175 ( .A(\data_in<8> ), .B(n1290), .Y(n28) );
  AND2X2 U176 ( .A(\data_in<9> ), .B(n1290), .Y(n29) );
  AND2X2 U177 ( .A(\data_in<10> ), .B(n1290), .Y(n30) );
  AND2X1 U178 ( .A(n16), .B(n1830), .Y(n31) );
  INVX1 U179 ( .A(n31), .Y(n32) );
  AND2X1 U180 ( .A(n1830), .B(n19), .Y(n33) );
  AND2X1 U181 ( .A(n1830), .B(n1694), .Y(n34) );
  INVX1 U182 ( .A(n34), .Y(n35) );
  AND2X1 U183 ( .A(n1830), .B(n1829), .Y(n36) );
  INVX1 U184 ( .A(n36), .Y(n37) );
  AND2X1 U185 ( .A(n15), .B(n16), .Y(n38) );
  INVX1 U186 ( .A(n38), .Y(n39) );
  AND2X1 U187 ( .A(n1290), .B(n38), .Y(n40) );
  INVX1 U188 ( .A(n40), .Y(n41) );
  AND2X1 U189 ( .A(n16), .B(n18), .Y(n42) );
  INVX1 U190 ( .A(n42), .Y(n43) );
  AND2X1 U191 ( .A(n1290), .B(n42), .Y(n44) );
  INVX1 U192 ( .A(n44), .Y(n45) );
  AND2X1 U193 ( .A(n16), .B(n1744), .Y(n46) );
  INVX1 U194 ( .A(n46), .Y(n47) );
  AND2X1 U195 ( .A(n1288), .B(n46), .Y(n48) );
  INVX1 U196 ( .A(n48), .Y(n49) );
  AND2X1 U197 ( .A(n16), .B(n1761), .Y(n50) );
  INVX1 U198 ( .A(n50), .Y(n51) );
  AND2X1 U199 ( .A(n1289), .B(n50), .Y(n52) );
  INVX1 U200 ( .A(n52), .Y(n53) );
  AND2X1 U201 ( .A(n16), .B(n1778), .Y(n54) );
  INVX1 U202 ( .A(n54), .Y(n55) );
  AND2X1 U203 ( .A(n1290), .B(n54), .Y(n56) );
  INVX1 U204 ( .A(n56), .Y(n57) );
  AND2X1 U205 ( .A(n16), .B(n1795), .Y(n58) );
  INVX1 U206 ( .A(n58), .Y(n59) );
  AND2X1 U207 ( .A(n1289), .B(n58), .Y(n60) );
  INVX1 U208 ( .A(n60), .Y(n61) );
  AND2X1 U209 ( .A(n16), .B(n1812), .Y(n62) );
  INVX1 U210 ( .A(n62), .Y(n63) );
  AND2X1 U211 ( .A(n1288), .B(n62), .Y(n64) );
  INVX1 U212 ( .A(n64), .Y(n65) );
  AND2X1 U213 ( .A(n1290), .B(n31), .Y(n66) );
  INVX1 U214 ( .A(n66), .Y(n67) );
  AND2X1 U215 ( .A(n15), .B(n19), .Y(n68) );
  INVX1 U216 ( .A(n68), .Y(n69) );
  AND2X1 U217 ( .A(n1290), .B(n68), .Y(n70) );
  INVX1 U218 ( .A(n70), .Y(n71) );
  AND2X1 U219 ( .A(n18), .B(n19), .Y(n72) );
  INVX1 U220 ( .A(n72), .Y(n73) );
  AND2X1 U221 ( .A(n1289), .B(n72), .Y(n74) );
  INVX1 U222 ( .A(n74), .Y(n75) );
  AND2X1 U223 ( .A(n1744), .B(n19), .Y(n76) );
  INVX1 U224 ( .A(n76), .Y(n77) );
  AND2X1 U225 ( .A(n1288), .B(n76), .Y(n78) );
  INVX1 U226 ( .A(n78), .Y(n79) );
  AND2X1 U227 ( .A(n1761), .B(n19), .Y(n80) );
  INVX1 U228 ( .A(n80), .Y(n81) );
  AND2X1 U229 ( .A(n1290), .B(n80), .Y(n82) );
  INVX1 U230 ( .A(n82), .Y(n83) );
  AND2X1 U231 ( .A(n1778), .B(n19), .Y(n84) );
  INVX1 U232 ( .A(n84), .Y(n85) );
  AND2X1 U233 ( .A(n1288), .B(n84), .Y(n86) );
  INVX1 U234 ( .A(n86), .Y(n87) );
  AND2X1 U235 ( .A(n1795), .B(n19), .Y(n88) );
  INVX1 U236 ( .A(n88), .Y(n89) );
  AND2X1 U237 ( .A(n1288), .B(n88), .Y(n90) );
  INVX1 U238 ( .A(n90), .Y(n91) );
  AND2X1 U239 ( .A(n1812), .B(n19), .Y(n92) );
  INVX1 U240 ( .A(n92), .Y(n93) );
  AND2X1 U241 ( .A(n1288), .B(n92), .Y(n94) );
  INVX1 U242 ( .A(n94), .Y(n95) );
  AND2X1 U243 ( .A(n1288), .B(n33), .Y(n96) );
  INVX1 U244 ( .A(n96), .Y(n97) );
  AND2X1 U245 ( .A(n15), .B(n1694), .Y(n98) );
  INVX1 U246 ( .A(n98), .Y(n99) );
  AND2X1 U247 ( .A(n1288), .B(n98), .Y(n100) );
  INVX1 U248 ( .A(n100), .Y(n101) );
  AND2X1 U249 ( .A(n18), .B(n1694), .Y(n102) );
  INVX1 U250 ( .A(n102), .Y(n103) );
  AND2X1 U251 ( .A(n1288), .B(n102), .Y(n104) );
  INVX1 U252 ( .A(n104), .Y(n105) );
  AND2X1 U253 ( .A(n1744), .B(n1694), .Y(n106) );
  INVX1 U254 ( .A(n106), .Y(n107) );
  AND2X1 U255 ( .A(n1288), .B(n106), .Y(n108) );
  INVX1 U256 ( .A(n108), .Y(n109) );
  AND2X1 U257 ( .A(n1761), .B(n1694), .Y(n110) );
  INVX1 U258 ( .A(n110), .Y(n111) );
  AND2X1 U259 ( .A(n1288), .B(n110), .Y(n112) );
  INVX1 U260 ( .A(n112), .Y(n113) );
  AND2X1 U261 ( .A(n1778), .B(n1694), .Y(n114) );
  INVX1 U262 ( .A(n114), .Y(n115) );
  AND2X1 U263 ( .A(n1288), .B(n114), .Y(n116) );
  INVX1 U264 ( .A(n116), .Y(n117) );
  AND2X1 U265 ( .A(n1795), .B(n1694), .Y(n118) );
  INVX1 U266 ( .A(n118), .Y(n119) );
  AND2X1 U267 ( .A(n1288), .B(n118), .Y(n120) );
  INVX1 U268 ( .A(n120), .Y(n121) );
  AND2X1 U269 ( .A(n1812), .B(n1694), .Y(n122) );
  INVX1 U270 ( .A(n122), .Y(n123) );
  AND2X1 U271 ( .A(n1288), .B(n122), .Y(n124) );
  INVX1 U272 ( .A(n124), .Y(n125) );
  AND2X1 U273 ( .A(n1289), .B(n34), .Y(n126) );
  INVX1 U274 ( .A(n126), .Y(n127) );
  AND2X1 U275 ( .A(n15), .B(n1829), .Y(n128) );
  INVX1 U276 ( .A(n128), .Y(n129) );
  AND2X1 U277 ( .A(n1289), .B(n128), .Y(n130) );
  INVX1 U278 ( .A(n130), .Y(n131) );
  AND2X1 U279 ( .A(n18), .B(n1829), .Y(n132) );
  INVX1 U280 ( .A(n132), .Y(n133) );
  AND2X1 U281 ( .A(n1289), .B(n132), .Y(n134) );
  INVX1 U282 ( .A(n134), .Y(n135) );
  AND2X1 U283 ( .A(n1744), .B(n1829), .Y(n136) );
  INVX1 U284 ( .A(n136), .Y(n137) );
  AND2X1 U285 ( .A(n1289), .B(n136), .Y(n138) );
  INVX1 U286 ( .A(n138), .Y(n139) );
  AND2X1 U287 ( .A(n1761), .B(n1829), .Y(n140) );
  INVX1 U288 ( .A(n140), .Y(n141) );
  AND2X1 U289 ( .A(n1289), .B(n140), .Y(n142) );
  INVX1 U290 ( .A(n142), .Y(n143) );
  AND2X1 U291 ( .A(n1778), .B(n1829), .Y(n144) );
  INVX1 U292 ( .A(n144), .Y(n145) );
  AND2X1 U293 ( .A(n1289), .B(n144), .Y(n146) );
  INVX1 U294 ( .A(n146), .Y(n147) );
  AND2X1 U295 ( .A(n1795), .B(n1829), .Y(n148) );
  INVX1 U296 ( .A(n148), .Y(n149) );
  AND2X1 U297 ( .A(n1289), .B(n148), .Y(n150) );
  INVX1 U298 ( .A(n150), .Y(n151) );
  AND2X1 U299 ( .A(n1812), .B(n1829), .Y(n152) );
  INVX1 U300 ( .A(n152), .Y(n153) );
  AND2X1 U301 ( .A(n1289), .B(n152), .Y(n154) );
  INVX1 U302 ( .A(n154), .Y(n155) );
  AND2X1 U303 ( .A(n1288), .B(n36), .Y(n156) );
  INVX1 U304 ( .A(n156), .Y(n157) );
  MUX2X1 U305 ( .B(n159), .A(n160), .S(n1177), .Y(n158) );
  MUX2X1 U306 ( .B(n162), .A(n163), .S(n1177), .Y(n161) );
  MUX2X1 U307 ( .B(n165), .A(n166), .S(n1177), .Y(n164) );
  MUX2X1 U308 ( .B(n168), .A(n169), .S(n1177), .Y(n167) );
  MUX2X1 U309 ( .B(n171), .A(n172), .S(n1170), .Y(n170) );
  MUX2X1 U310 ( .B(n174), .A(n175), .S(n1177), .Y(n173) );
  MUX2X1 U311 ( .B(n177), .A(n178), .S(n1177), .Y(n176) );
  MUX2X1 U312 ( .B(n180), .A(n181), .S(n1177), .Y(n179) );
  MUX2X1 U313 ( .B(n183), .A(n184), .S(n1177), .Y(n182) );
  MUX2X1 U314 ( .B(n186), .A(n187), .S(n1170), .Y(n185) );
  MUX2X1 U315 ( .B(n189), .A(n190), .S(n1178), .Y(n188) );
  MUX2X1 U316 ( .B(n192), .A(n193), .S(n1178), .Y(n191) );
  MUX2X1 U317 ( .B(n195), .A(n196), .S(n1178), .Y(n194) );
  MUX2X1 U318 ( .B(n198), .A(n199), .S(n1178), .Y(n197) );
  MUX2X1 U319 ( .B(n201), .A(n202), .S(n1170), .Y(n200) );
  MUX2X1 U320 ( .B(n204), .A(n205), .S(n1178), .Y(n203) );
  MUX2X1 U321 ( .B(n207), .A(n208), .S(n1178), .Y(n206) );
  MUX2X1 U322 ( .B(n210), .A(n211), .S(n1178), .Y(n209) );
  MUX2X1 U323 ( .B(n213), .A(n215), .S(n1178), .Y(n212) );
  MUX2X1 U324 ( .B(n217), .A(n218), .S(n1170), .Y(n216) );
  MUX2X1 U325 ( .B(n220), .A(n221), .S(n1178), .Y(n219) );
  MUX2X1 U326 ( .B(n223), .A(n224), .S(n1178), .Y(n222) );
  MUX2X1 U327 ( .B(n226), .A(n227), .S(n1178), .Y(n225) );
  MUX2X1 U328 ( .B(n229), .A(n230), .S(n1178), .Y(n228) );
  MUX2X1 U329 ( .B(n232), .A(n233), .S(n1170), .Y(n231) );
  MUX2X1 U330 ( .B(n235), .A(n236), .S(n1179), .Y(n234) );
  MUX2X1 U331 ( .B(n238), .A(n239), .S(n1179), .Y(n237) );
  MUX2X1 U332 ( .B(n241), .A(n242), .S(n1179), .Y(n240) );
  MUX2X1 U333 ( .B(n244), .A(n245), .S(n1179), .Y(n243) );
  MUX2X1 U334 ( .B(n247), .A(n248), .S(n1170), .Y(n246) );
  MUX2X1 U335 ( .B(n250), .A(n251), .S(n1179), .Y(n249) );
  MUX2X1 U336 ( .B(n253), .A(n254), .S(n1179), .Y(n252) );
  MUX2X1 U337 ( .B(n256), .A(n257), .S(n1179), .Y(n255) );
  MUX2X1 U338 ( .B(n259), .A(n260), .S(n1179), .Y(n258) );
  MUX2X1 U339 ( .B(n262), .A(n263), .S(n1170), .Y(n261) );
  MUX2X1 U340 ( .B(n265), .A(n266), .S(n1179), .Y(n264) );
  MUX2X1 U341 ( .B(n268), .A(n269), .S(n1179), .Y(n267) );
  MUX2X1 U342 ( .B(n271), .A(n272), .S(n1179), .Y(n270) );
  MUX2X1 U343 ( .B(n274), .A(n275), .S(n1179), .Y(n273) );
  MUX2X1 U344 ( .B(n277), .A(n278), .S(n1170), .Y(n276) );
  MUX2X1 U345 ( .B(n280), .A(n281), .S(n1180), .Y(n279) );
  MUX2X1 U346 ( .B(n283), .A(n284), .S(n1180), .Y(n282) );
  MUX2X1 U347 ( .B(n286), .A(n287), .S(n1180), .Y(n285) );
  MUX2X1 U348 ( .B(n289), .A(n290), .S(n1180), .Y(n288) );
  MUX2X1 U349 ( .B(n292), .A(n293), .S(n1170), .Y(n291) );
  MUX2X1 U350 ( .B(n295), .A(n296), .S(n1180), .Y(n294) );
  MUX2X1 U351 ( .B(n298), .A(n299), .S(n1180), .Y(n297) );
  MUX2X1 U352 ( .B(n301), .A(n302), .S(n1180), .Y(n300) );
  MUX2X1 U353 ( .B(n304), .A(n305), .S(n1180), .Y(n303) );
  MUX2X1 U354 ( .B(n307), .A(n308), .S(n1170), .Y(n306) );
  MUX2X1 U355 ( .B(n310), .A(n311), .S(n1180), .Y(n309) );
  MUX2X1 U356 ( .B(n313), .A(n314), .S(n1180), .Y(n312) );
  MUX2X1 U357 ( .B(n316), .A(n317), .S(n1180), .Y(n315) );
  MUX2X1 U358 ( .B(n319), .A(n320), .S(n1180), .Y(n318) );
  MUX2X1 U359 ( .B(n322), .A(n323), .S(n1170), .Y(n321) );
  MUX2X1 U360 ( .B(n325), .A(n326), .S(n1181), .Y(n324) );
  MUX2X1 U361 ( .B(n328), .A(n329), .S(n1181), .Y(n327) );
  MUX2X1 U362 ( .B(n331), .A(n332), .S(n1181), .Y(n330) );
  MUX2X1 U363 ( .B(n334), .A(n335), .S(n1181), .Y(n333) );
  MUX2X1 U364 ( .B(n337), .A(n338), .S(n1170), .Y(n336) );
  MUX2X1 U365 ( .B(n340), .A(n341), .S(n1181), .Y(n339) );
  MUX2X1 U366 ( .B(n343), .A(n344), .S(n1181), .Y(n342) );
  MUX2X1 U367 ( .B(n346), .A(n347), .S(n1181), .Y(n345) );
  MUX2X1 U368 ( .B(n349), .A(n350), .S(n1181), .Y(n348) );
  MUX2X1 U369 ( .B(n352), .A(n353), .S(n1169), .Y(n351) );
  MUX2X1 U370 ( .B(n355), .A(n356), .S(n1181), .Y(n354) );
  MUX2X1 U371 ( .B(n358), .A(n359), .S(n1181), .Y(n357) );
  MUX2X1 U372 ( .B(n361), .A(n362), .S(n1181), .Y(n360) );
  MUX2X1 U373 ( .B(n364), .A(n365), .S(n1181), .Y(n363) );
  MUX2X1 U374 ( .B(n367), .A(n368), .S(n1169), .Y(n366) );
  MUX2X1 U375 ( .B(n370), .A(n371), .S(n1182), .Y(n369) );
  MUX2X1 U376 ( .B(n373), .A(n374), .S(n1182), .Y(n372) );
  MUX2X1 U377 ( .B(n376), .A(n377), .S(n1182), .Y(n375) );
  MUX2X1 U378 ( .B(n379), .A(n380), .S(n1182), .Y(n378) );
  MUX2X1 U379 ( .B(n382), .A(n383), .S(n1169), .Y(n381) );
  MUX2X1 U380 ( .B(n385), .A(n386), .S(n1182), .Y(n384) );
  MUX2X1 U381 ( .B(n388), .A(n389), .S(n1182), .Y(n387) );
  MUX2X1 U382 ( .B(n391), .A(n392), .S(n1182), .Y(n390) );
  MUX2X1 U383 ( .B(n394), .A(n395), .S(n1182), .Y(n393) );
  MUX2X1 U384 ( .B(n397), .A(n398), .S(n1169), .Y(n396) );
  MUX2X1 U385 ( .B(n400), .A(n401), .S(n1182), .Y(n399) );
  MUX2X1 U386 ( .B(n403), .A(n404), .S(n1182), .Y(n402) );
  MUX2X1 U387 ( .B(n406), .A(n407), .S(n1182), .Y(n405) );
  MUX2X1 U388 ( .B(n409), .A(n410), .S(n1182), .Y(n408) );
  MUX2X1 U389 ( .B(n412), .A(n413), .S(n1169), .Y(n411) );
  MUX2X1 U390 ( .B(n415), .A(n416), .S(n1183), .Y(n414) );
  MUX2X1 U391 ( .B(n418), .A(n419), .S(n1183), .Y(n417) );
  MUX2X1 U392 ( .B(n421), .A(n422), .S(n1183), .Y(n420) );
  MUX2X1 U393 ( .B(n424), .A(n425), .S(n1183), .Y(n423) );
  MUX2X1 U394 ( .B(n427), .A(n428), .S(n1169), .Y(n426) );
  MUX2X1 U395 ( .B(n430), .A(n431), .S(n1183), .Y(n429) );
  MUX2X1 U396 ( .B(n433), .A(n434), .S(n1183), .Y(n432) );
  MUX2X1 U397 ( .B(n436), .A(n437), .S(n1183), .Y(n435) );
  MUX2X1 U398 ( .B(n439), .A(n440), .S(n1183), .Y(n438) );
  MUX2X1 U399 ( .B(n442), .A(n443), .S(n1169), .Y(n441) );
  MUX2X1 U400 ( .B(n445), .A(n446), .S(n1183), .Y(n444) );
  MUX2X1 U401 ( .B(n448), .A(n449), .S(n1183), .Y(n447) );
  MUX2X1 U402 ( .B(n451), .A(n452), .S(n1183), .Y(n450) );
  MUX2X1 U403 ( .B(n454), .A(n455), .S(n1183), .Y(n453) );
  MUX2X1 U404 ( .B(n457), .A(n458), .S(n1169), .Y(n456) );
  MUX2X1 U405 ( .B(n460), .A(n461), .S(n1183), .Y(n459) );
  MUX2X1 U406 ( .B(n463), .A(n464), .S(n1183), .Y(n462) );
  MUX2X1 U407 ( .B(n466), .A(n467), .S(n1183), .Y(n465) );
  MUX2X1 U408 ( .B(n469), .A(n470), .S(n1183), .Y(n468) );
  MUX2X1 U409 ( .B(n472), .A(n473), .S(n1169), .Y(n471) );
  MUX2X1 U410 ( .B(n475), .A(n476), .S(n1183), .Y(n474) );
  MUX2X1 U411 ( .B(n478), .A(n479), .S(n1183), .Y(n477) );
  MUX2X1 U412 ( .B(n481), .A(n482), .S(n1184), .Y(n480) );
  MUX2X1 U413 ( .B(n484), .A(n485), .S(n1183), .Y(n483) );
  MUX2X1 U414 ( .B(n487), .A(n488), .S(n1169), .Y(n486) );
  MUX2X1 U415 ( .B(n490), .A(n491), .S(n1184), .Y(n489) );
  MUX2X1 U416 ( .B(n493), .A(n494), .S(n1184), .Y(n492) );
  MUX2X1 U417 ( .B(n496), .A(n497), .S(n1184), .Y(n495) );
  MUX2X1 U418 ( .B(n499), .A(n500), .S(n1183), .Y(n498) );
  MUX2X1 U419 ( .B(n502), .A(n503), .S(n1169), .Y(n501) );
  MUX2X1 U420 ( .B(n505), .A(n506), .S(n1184), .Y(n504) );
  MUX2X1 U421 ( .B(n508), .A(n509), .S(n1184), .Y(n507) );
  MUX2X1 U422 ( .B(n511), .A(n512), .S(n1184), .Y(n510) );
  MUX2X1 U423 ( .B(n514), .A(n515), .S(n1184), .Y(n513) );
  MUX2X1 U424 ( .B(n517), .A(n518), .S(n1169), .Y(n516) );
  MUX2X1 U425 ( .B(n520), .A(n521), .S(n1184), .Y(n519) );
  MUX2X1 U426 ( .B(n523), .A(n524), .S(n1184), .Y(n522) );
  MUX2X1 U427 ( .B(n526), .A(n527), .S(n1184), .Y(n525) );
  MUX2X1 U428 ( .B(n529), .A(n530), .S(n1184), .Y(n528) );
  MUX2X1 U429 ( .B(n532), .A(n533), .S(n1168), .Y(n531) );
  MUX2X1 U430 ( .B(n535), .A(n536), .S(n1184), .Y(n534) );
  MUX2X1 U431 ( .B(n538), .A(n539), .S(n1184), .Y(n537) );
  MUX2X1 U432 ( .B(n541), .A(n542), .S(n1184), .Y(n540) );
  MUX2X1 U433 ( .B(n544), .A(n545), .S(n1184), .Y(n543) );
  MUX2X1 U434 ( .B(n547), .A(n548), .S(n1168), .Y(n546) );
  MUX2X1 U435 ( .B(n550), .A(n551), .S(n1185), .Y(n549) );
  MUX2X1 U436 ( .B(n553), .A(n554), .S(n1185), .Y(n552) );
  MUX2X1 U437 ( .B(n556), .A(n557), .S(n1185), .Y(n555) );
  MUX2X1 U438 ( .B(n559), .A(n560), .S(n1185), .Y(n558) );
  MUX2X1 U439 ( .B(n562), .A(n563), .S(n1168), .Y(n561) );
  MUX2X1 U440 ( .B(n565), .A(n566), .S(n1185), .Y(n564) );
  MUX2X1 U441 ( .B(n568), .A(n569), .S(n1185), .Y(n567) );
  MUX2X1 U442 ( .B(n571), .A(n572), .S(n1185), .Y(n570) );
  MUX2X1 U443 ( .B(n574), .A(n575), .S(n1185), .Y(n573) );
  MUX2X1 U444 ( .B(n577), .A(n578), .S(n1168), .Y(n576) );
  MUX2X1 U445 ( .B(n580), .A(n581), .S(n1185), .Y(n579) );
  MUX2X1 U446 ( .B(n583), .A(n584), .S(n1185), .Y(n582) );
  MUX2X1 U447 ( .B(n586), .A(n587), .S(n1185), .Y(n585) );
  MUX2X1 U448 ( .B(n589), .A(n590), .S(n1185), .Y(n588) );
  MUX2X1 U449 ( .B(n592), .A(n593), .S(n1168), .Y(n591) );
  MUX2X1 U450 ( .B(n595), .A(n596), .S(n1186), .Y(n594) );
  MUX2X1 U451 ( .B(n598), .A(n599), .S(n1186), .Y(n597) );
  MUX2X1 U452 ( .B(n601), .A(n602), .S(n1186), .Y(n600) );
  MUX2X1 U453 ( .B(n604), .A(n605), .S(n1186), .Y(n603) );
  MUX2X1 U454 ( .B(n607), .A(n608), .S(n1168), .Y(n606) );
  MUX2X1 U455 ( .B(n610), .A(n611), .S(n1186), .Y(n609) );
  MUX2X1 U456 ( .B(n613), .A(n614), .S(n1186), .Y(n612) );
  MUX2X1 U457 ( .B(n616), .A(n617), .S(n1186), .Y(n615) );
  MUX2X1 U458 ( .B(n619), .A(n620), .S(n1186), .Y(n618) );
  MUX2X1 U459 ( .B(n622), .A(n623), .S(n1168), .Y(n621) );
  MUX2X1 U460 ( .B(n625), .A(n626), .S(n1186), .Y(n624) );
  MUX2X1 U461 ( .B(n628), .A(n629), .S(n1186), .Y(n627) );
  MUX2X1 U462 ( .B(n631), .A(n632), .S(n1186), .Y(n630) );
  MUX2X1 U463 ( .B(n634), .A(n635), .S(n1186), .Y(n633) );
  MUX2X1 U464 ( .B(n637), .A(n638), .S(n1168), .Y(n636) );
  MUX2X1 U465 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1191), .Y(n160) );
  MUX2X1 U466 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1191), .Y(n159) );
  MUX2X1 U467 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1191), .Y(n163) );
  MUX2X1 U468 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1191), .Y(n162) );
  MUX2X1 U469 ( .B(n161), .A(n158), .S(n1174), .Y(n172) );
  MUX2X1 U470 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1197), .Y(n166) );
  MUX2X1 U471 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1191), .Y(n165) );
  MUX2X1 U472 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1204), .Y(n169) );
  MUX2X1 U473 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1204), .Y(n168) );
  MUX2X1 U474 ( .B(n167), .A(n164), .S(n1174), .Y(n171) );
  MUX2X1 U475 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1202), .Y(n175) );
  MUX2X1 U476 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1200), .Y(n174) );
  MUX2X1 U477 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1191), .Y(n178) );
  MUX2X1 U478 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1191), .Y(n177) );
  MUX2X1 U479 ( .B(n176), .A(n173), .S(n1174), .Y(n187) );
  MUX2X1 U480 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1202), .Y(n181) );
  MUX2X1 U481 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1202), .Y(n180) );
  MUX2X1 U482 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1191), .Y(n184) );
  MUX2X1 U483 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1200), .Y(n183) );
  MUX2X1 U484 ( .B(n182), .A(n179), .S(n1174), .Y(n186) );
  MUX2X1 U485 ( .B(n185), .A(n170), .S(n1167), .Y(n639) );
  MUX2X1 U486 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1199), .Y(n190) );
  MUX2X1 U487 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1199), .Y(n189) );
  MUX2X1 U488 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1308), .Y(n193) );
  MUX2X1 U489 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1198), .Y(n192) );
  MUX2X1 U490 ( .B(n191), .A(n188), .S(n1174), .Y(n202) );
  MUX2X1 U491 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1198), .Y(n196) );
  MUX2X1 U492 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1308), .Y(n195) );
  MUX2X1 U493 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1199), .Y(n199) );
  MUX2X1 U494 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1308), .Y(n198) );
  MUX2X1 U495 ( .B(n197), .A(n194), .S(n1174), .Y(n201) );
  MUX2X1 U496 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1308), .Y(n205) );
  MUX2X1 U497 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1198), .Y(n204) );
  MUX2X1 U498 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1308), .Y(n208) );
  MUX2X1 U499 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1308), .Y(n207) );
  MUX2X1 U500 ( .B(n206), .A(n203), .S(n1174), .Y(n218) );
  MUX2X1 U501 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1192), .Y(n211) );
  MUX2X1 U502 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1192), .Y(n210) );
  MUX2X1 U503 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1192), .Y(n215) );
  MUX2X1 U504 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1192), .Y(n213) );
  MUX2X1 U505 ( .B(n212), .A(n209), .S(n1174), .Y(n217) );
  MUX2X1 U506 ( .B(n216), .A(n200), .S(n1167), .Y(n640) );
  MUX2X1 U507 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1192), .Y(n221) );
  MUX2X1 U508 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1192), .Y(n220) );
  MUX2X1 U509 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1192), .Y(n224) );
  MUX2X1 U510 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1192), .Y(n223) );
  MUX2X1 U511 ( .B(n222), .A(n219), .S(n1174), .Y(n233) );
  MUX2X1 U512 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1192), .Y(n227) );
  MUX2X1 U513 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1192), .Y(n226) );
  MUX2X1 U514 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1192), .Y(n230) );
  MUX2X1 U515 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1192), .Y(n229) );
  MUX2X1 U516 ( .B(n228), .A(n225), .S(n1174), .Y(n232) );
  MUX2X1 U517 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1193), .Y(n236) );
  MUX2X1 U518 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1193), .Y(n235) );
  MUX2X1 U519 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1193), .Y(n239) );
  MUX2X1 U520 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1193), .Y(n238) );
  MUX2X1 U521 ( .B(n237), .A(n234), .S(n1174), .Y(n248) );
  MUX2X1 U522 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1193), .Y(n242) );
  MUX2X1 U523 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1193), .Y(n241) );
  MUX2X1 U524 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1193), .Y(n245) );
  MUX2X1 U525 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1193), .Y(n244) );
  MUX2X1 U526 ( .B(n243), .A(n240), .S(n1174), .Y(n247) );
  MUX2X1 U527 ( .B(n246), .A(n231), .S(n1167), .Y(n641) );
  MUX2X1 U528 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1193), .Y(n251) );
  MUX2X1 U529 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1193), .Y(n250) );
  MUX2X1 U530 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1193), .Y(n254) );
  MUX2X1 U531 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1193), .Y(n253) );
  MUX2X1 U532 ( .B(n252), .A(n249), .S(n1173), .Y(n263) );
  MUX2X1 U533 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1194), .Y(n257) );
  MUX2X1 U534 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1194), .Y(n256) );
  MUX2X1 U535 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1194), .Y(n260) );
  MUX2X1 U536 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1194), .Y(n259) );
  MUX2X1 U537 ( .B(n258), .A(n255), .S(n1173), .Y(n262) );
  MUX2X1 U538 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1194), .Y(n266) );
  MUX2X1 U539 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1194), .Y(n265) );
  MUX2X1 U540 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1194), .Y(n269) );
  MUX2X1 U541 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1194), .Y(n268) );
  MUX2X1 U542 ( .B(n267), .A(n264), .S(n1173), .Y(n278) );
  MUX2X1 U543 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1194), .Y(n272) );
  MUX2X1 U544 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1194), .Y(n271) );
  MUX2X1 U545 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1194), .Y(n275) );
  MUX2X1 U546 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1194), .Y(n274) );
  MUX2X1 U547 ( .B(n273), .A(n270), .S(n1173), .Y(n277) );
  MUX2X1 U548 ( .B(n276), .A(n261), .S(n1167), .Y(n642) );
  MUX2X1 U549 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1195), .Y(n281) );
  MUX2X1 U550 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1195), .Y(n280) );
  MUX2X1 U551 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1195), .Y(n284) );
  MUX2X1 U552 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1195), .Y(n283) );
  MUX2X1 U553 ( .B(n282), .A(n279), .S(n1173), .Y(n293) );
  MUX2X1 U554 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1195), .Y(n287) );
  MUX2X1 U555 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1195), .Y(n286) );
  MUX2X1 U556 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1195), .Y(n290) );
  MUX2X1 U557 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1195), .Y(n289) );
  MUX2X1 U558 ( .B(n288), .A(n285), .S(n1173), .Y(n292) );
  MUX2X1 U559 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1195), .Y(n296) );
  MUX2X1 U560 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1195), .Y(n295) );
  MUX2X1 U561 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1195), .Y(n299) );
  MUX2X1 U562 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1195), .Y(n298) );
  MUX2X1 U563 ( .B(n297), .A(n294), .S(n1173), .Y(n308) );
  MUX2X1 U564 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1196), .Y(n302) );
  MUX2X1 U565 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1196), .Y(n301) );
  MUX2X1 U566 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1196), .Y(n305) );
  MUX2X1 U567 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1196), .Y(n304) );
  MUX2X1 U568 ( .B(n303), .A(n300), .S(n1173), .Y(n307) );
  MUX2X1 U569 ( .B(n306), .A(n291), .S(n1167), .Y(n643) );
  MUX2X1 U570 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1196), .Y(n311) );
  MUX2X1 U571 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1196), .Y(n310) );
  MUX2X1 U572 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1196), .Y(n314) );
  MUX2X1 U573 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1196), .Y(n313) );
  MUX2X1 U574 ( .B(n312), .A(n309), .S(n1173), .Y(n323) );
  MUX2X1 U575 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1196), .Y(n317) );
  MUX2X1 U576 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1196), .Y(n316) );
  MUX2X1 U577 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1196), .Y(n320) );
  MUX2X1 U578 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1196), .Y(n319) );
  MUX2X1 U579 ( .B(n318), .A(n315), .S(n1173), .Y(n322) );
  MUX2X1 U580 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1197), .Y(n326) );
  MUX2X1 U581 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1197), .Y(n325) );
  MUX2X1 U582 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1197), .Y(n329) );
  MUX2X1 U583 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1197), .Y(n328) );
  MUX2X1 U584 ( .B(n327), .A(n324), .S(n1173), .Y(n338) );
  MUX2X1 U585 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1197), .Y(n332) );
  MUX2X1 U586 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1197), .Y(n331) );
  MUX2X1 U587 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1197), .Y(n335) );
  MUX2X1 U588 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1197), .Y(n334) );
  MUX2X1 U589 ( .B(n333), .A(n330), .S(n1173), .Y(n337) );
  MUX2X1 U590 ( .B(n336), .A(n321), .S(n1167), .Y(n644) );
  MUX2X1 U591 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1197), .Y(n341) );
  MUX2X1 U592 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1197), .Y(n340) );
  MUX2X1 U593 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1197), .Y(n344) );
  MUX2X1 U594 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1197), .Y(n343) );
  MUX2X1 U595 ( .B(n342), .A(n339), .S(n1173), .Y(n353) );
  MUX2X1 U596 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1198), .Y(n347) );
  MUX2X1 U597 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1198), .Y(n346) );
  MUX2X1 U598 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1198), .Y(n350) );
  MUX2X1 U599 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1198), .Y(n349) );
  MUX2X1 U600 ( .B(n348), .A(n345), .S(n1174), .Y(n352) );
  MUX2X1 U601 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1198), .Y(n356) );
  MUX2X1 U602 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1198), .Y(n355) );
  MUX2X1 U603 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1198), .Y(n359) );
  MUX2X1 U604 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1198), .Y(n358) );
  MUX2X1 U605 ( .B(n357), .A(n354), .S(n1173), .Y(n368) );
  MUX2X1 U606 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1198), .Y(n362) );
  MUX2X1 U607 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1198), .Y(n361) );
  MUX2X1 U608 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1198), .Y(n365) );
  MUX2X1 U609 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1198), .Y(n364) );
  MUX2X1 U610 ( .B(n363), .A(n360), .S(n1173), .Y(n367) );
  MUX2X1 U611 ( .B(n366), .A(n351), .S(n1167), .Y(n645) );
  MUX2X1 U612 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1199), .Y(n371) );
  MUX2X1 U613 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1199), .Y(n370) );
  MUX2X1 U614 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1199), .Y(n374) );
  MUX2X1 U615 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1199), .Y(n373) );
  MUX2X1 U616 ( .B(n372), .A(n369), .S(n1173), .Y(n383) );
  MUX2X1 U617 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1199), .Y(n377) );
  MUX2X1 U618 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1199), .Y(n376) );
  MUX2X1 U619 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1199), .Y(n380) );
  MUX2X1 U620 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1199), .Y(n379) );
  MUX2X1 U621 ( .B(n378), .A(n375), .S(n1173), .Y(n382) );
  MUX2X1 U622 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1199), .Y(n386) );
  MUX2X1 U623 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1199), .Y(n385) );
  MUX2X1 U624 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1199), .Y(n389) );
  MUX2X1 U625 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1199), .Y(n388) );
  MUX2X1 U626 ( .B(n387), .A(n384), .S(n1174), .Y(n398) );
  MUX2X1 U627 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1200), .Y(n392) );
  MUX2X1 U628 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1200), .Y(n391) );
  MUX2X1 U629 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1200), .Y(n395) );
  MUX2X1 U630 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1200), .Y(n394) );
  MUX2X1 U631 ( .B(n393), .A(n390), .S(n1174), .Y(n397) );
  MUX2X1 U632 ( .B(n396), .A(n381), .S(n1167), .Y(n646) );
  MUX2X1 U633 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1200), .Y(n401) );
  MUX2X1 U634 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1200), .Y(n400) );
  MUX2X1 U635 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1200), .Y(n404) );
  MUX2X1 U636 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1200), .Y(n403) );
  MUX2X1 U637 ( .B(n402), .A(n399), .S(n1174), .Y(n413) );
  MUX2X1 U638 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1200), .Y(n407) );
  MUX2X1 U639 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1200), .Y(n406) );
  MUX2X1 U640 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1200), .Y(n410) );
  MUX2X1 U641 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1200), .Y(n409) );
  MUX2X1 U642 ( .B(n408), .A(n405), .S(n1173), .Y(n412) );
  MUX2X1 U643 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1201), .Y(n416) );
  MUX2X1 U644 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1201), .Y(n415) );
  MUX2X1 U645 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1201), .Y(n419) );
  MUX2X1 U646 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1201), .Y(n418) );
  MUX2X1 U647 ( .B(n417), .A(n414), .S(n1174), .Y(n428) );
  MUX2X1 U648 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1201), .Y(n422) );
  MUX2X1 U649 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1201), .Y(n421) );
  MUX2X1 U650 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1201), .Y(n425) );
  MUX2X1 U651 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1201), .Y(n424) );
  MUX2X1 U652 ( .B(n423), .A(n420), .S(n1174), .Y(n427) );
  MUX2X1 U653 ( .B(n426), .A(n411), .S(n1167), .Y(n647) );
  MUX2X1 U654 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1201), .Y(n431) );
  MUX2X1 U655 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1201), .Y(n430) );
  MUX2X1 U656 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1201), .Y(n434) );
  MUX2X1 U657 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1201), .Y(n433) );
  MUX2X1 U658 ( .B(n432), .A(n429), .S(n1172), .Y(n443) );
  MUX2X1 U659 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1202), .Y(n437) );
  MUX2X1 U660 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1202), .Y(n436) );
  MUX2X1 U661 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1202), .Y(n440) );
  MUX2X1 U662 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1202), .Y(n439) );
  MUX2X1 U663 ( .B(n438), .A(n435), .S(n1172), .Y(n442) );
  MUX2X1 U664 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1202), .Y(n446) );
  MUX2X1 U665 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1202), .Y(n445) );
  MUX2X1 U666 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1202), .Y(n449) );
  MUX2X1 U667 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1202), .Y(n448) );
  MUX2X1 U668 ( .B(n447), .A(n444), .S(n1172), .Y(n458) );
  MUX2X1 U669 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1202), .Y(n452) );
  MUX2X1 U670 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1202), .Y(n451) );
  MUX2X1 U671 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1202), .Y(n455) );
  MUX2X1 U672 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1202), .Y(n454) );
  MUX2X1 U673 ( .B(n453), .A(n450), .S(n1172), .Y(n457) );
  MUX2X1 U674 ( .B(n456), .A(n441), .S(n1167), .Y(n648) );
  MUX2X1 U675 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1205), .Y(n461) );
  MUX2X1 U676 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1205), .Y(n460) );
  MUX2X1 U677 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1205), .Y(n464) );
  MUX2X1 U678 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1205), .Y(n463) );
  MUX2X1 U679 ( .B(n462), .A(n459), .S(n1172), .Y(n473) );
  MUX2X1 U680 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1205), .Y(n467) );
  MUX2X1 U681 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1205), .Y(n466) );
  MUX2X1 U682 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1205), .Y(n470) );
  MUX2X1 U683 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1205), .Y(n469) );
  MUX2X1 U684 ( .B(n468), .A(n465), .S(n1172), .Y(n472) );
  MUX2X1 U685 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1205), .Y(n476) );
  MUX2X1 U686 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1205), .Y(n475) );
  MUX2X1 U687 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1205), .Y(n479) );
  MUX2X1 U688 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1205), .Y(n478) );
  MUX2X1 U689 ( .B(n477), .A(n474), .S(n1172), .Y(n488) );
  MUX2X1 U690 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1203), .Y(n482) );
  MUX2X1 U691 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1203), .Y(n481) );
  MUX2X1 U692 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1203), .Y(n485) );
  MUX2X1 U693 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1203), .Y(n484) );
  MUX2X1 U694 ( .B(n483), .A(n480), .S(n1172), .Y(n487) );
  MUX2X1 U695 ( .B(n486), .A(n471), .S(n1167), .Y(n649) );
  MUX2X1 U696 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1203), .Y(n491) );
  MUX2X1 U697 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1203), .Y(n490) );
  MUX2X1 U698 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1203), .Y(n494) );
  MUX2X1 U699 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1203), .Y(n493) );
  MUX2X1 U700 ( .B(n492), .A(n489), .S(n1172), .Y(n503) );
  MUX2X1 U701 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1203), .Y(n497) );
  MUX2X1 U702 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1203), .Y(n496) );
  MUX2X1 U703 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1203), .Y(n500) );
  MUX2X1 U704 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1203), .Y(n499) );
  MUX2X1 U705 ( .B(n498), .A(n495), .S(n1172), .Y(n502) );
  MUX2X1 U706 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1206), .Y(n506) );
  MUX2X1 U707 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1206), .Y(n505) );
  MUX2X1 U708 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1204), .Y(n509) );
  MUX2X1 U709 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1204), .Y(n508) );
  MUX2X1 U710 ( .B(n507), .A(n504), .S(n1172), .Y(n518) );
  MUX2X1 U711 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1204), .Y(n512) );
  MUX2X1 U712 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1202), .Y(n511) );
  MUX2X1 U713 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1205), .Y(n515) );
  MUX2X1 U714 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1206), .Y(n514) );
  MUX2X1 U715 ( .B(n513), .A(n510), .S(n1172), .Y(n517) );
  MUX2X1 U716 ( .B(n516), .A(n501), .S(n1167), .Y(n650) );
  MUX2X1 U717 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1204), .Y(n521) );
  MUX2X1 U718 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1202), .Y(n520) );
  MUX2X1 U719 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1204), .Y(n524) );
  MUX2X1 U720 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1206), .Y(n523) );
  MUX2X1 U721 ( .B(n522), .A(n519), .S(n1172), .Y(n533) );
  MUX2X1 U722 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1203), .Y(n527) );
  MUX2X1 U723 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1202), .Y(n526) );
  MUX2X1 U724 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1204), .Y(n530) );
  MUX2X1 U725 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1203), .Y(n529) );
  MUX2X1 U726 ( .B(n528), .A(n525), .S(n1172), .Y(n532) );
  MUX2X1 U727 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1202), .Y(n536) );
  MUX2X1 U728 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1204), .Y(n535) );
  MUX2X1 U729 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1203), .Y(n539) );
  MUX2X1 U730 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1203), .Y(n538) );
  MUX2X1 U731 ( .B(n537), .A(n534), .S(n1172), .Y(n548) );
  MUX2X1 U732 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1203), .Y(n542) );
  MUX2X1 U733 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1203), .Y(n541) );
  MUX2X1 U734 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1203), .Y(n545) );
  MUX2X1 U735 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1203), .Y(n544) );
  MUX2X1 U736 ( .B(n543), .A(n540), .S(n1172), .Y(n547) );
  MUX2X1 U737 ( .B(n546), .A(n531), .S(n1167), .Y(n1163) );
  MUX2X1 U738 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1202), .Y(n551) );
  MUX2X1 U739 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1203), .Y(n550) );
  MUX2X1 U740 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1205), .Y(n554) );
  MUX2X1 U741 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1203), .Y(n553) );
  MUX2X1 U742 ( .B(n552), .A(n549), .S(n1172), .Y(n563) );
  MUX2X1 U743 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1202), .Y(n557) );
  MUX2X1 U744 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1201), .Y(n556) );
  MUX2X1 U745 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1205), .Y(n560) );
  MUX2X1 U746 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1202), .Y(n559) );
  MUX2X1 U747 ( .B(n558), .A(n555), .S(n1172), .Y(n562) );
  MUX2X1 U748 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1205), .Y(n566) );
  MUX2X1 U749 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1205), .Y(n565) );
  MUX2X1 U750 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1205), .Y(n569) );
  MUX2X1 U751 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1205), .Y(n568) );
  MUX2X1 U752 ( .B(n567), .A(n564), .S(n1172), .Y(n578) );
  MUX2X1 U753 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1204), .Y(n572) );
  MUX2X1 U754 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1204), .Y(n571) );
  MUX2X1 U755 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1204), .Y(n575) );
  MUX2X1 U756 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1204), .Y(n574) );
  MUX2X1 U757 ( .B(n573), .A(n570), .S(n1172), .Y(n577) );
  MUX2X1 U758 ( .B(n576), .A(n561), .S(n1167), .Y(n1164) );
  MUX2X1 U759 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1204), .Y(n581) );
  MUX2X1 U760 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1204), .Y(n580) );
  MUX2X1 U761 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1204), .Y(n584) );
  MUX2X1 U762 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1204), .Y(n583) );
  MUX2X1 U763 ( .B(n582), .A(n579), .S(n1172), .Y(n593) );
  MUX2X1 U764 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1204), .Y(n587) );
  MUX2X1 U765 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1204), .Y(n586) );
  MUX2X1 U766 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1204), .Y(n590) );
  MUX2X1 U767 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1204), .Y(n589) );
  MUX2X1 U768 ( .B(n588), .A(n585), .S(n1172), .Y(n592) );
  MUX2X1 U769 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1205), .Y(n596) );
  MUX2X1 U770 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1205), .Y(n595) );
  MUX2X1 U771 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1205), .Y(n599) );
  MUX2X1 U772 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1205), .Y(n598) );
  MUX2X1 U773 ( .B(n597), .A(n594), .S(n1172), .Y(n608) );
  MUX2X1 U774 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1205), .Y(n602) );
  MUX2X1 U775 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1205), .Y(n601) );
  MUX2X1 U776 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1205), .Y(n605) );
  MUX2X1 U777 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1205), .Y(n604) );
  MUX2X1 U778 ( .B(n603), .A(n600), .S(n1172), .Y(n607) );
  MUX2X1 U779 ( .B(n606), .A(n591), .S(n1167), .Y(n1165) );
  MUX2X1 U780 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1205), .Y(n611) );
  MUX2X1 U781 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1205), .Y(n610) );
  MUX2X1 U782 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1205), .Y(n614) );
  MUX2X1 U783 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1205), .Y(n613) );
  MUX2X1 U784 ( .B(n612), .A(n609), .S(n1172), .Y(n623) );
  MUX2X1 U785 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1206), .Y(n617) );
  MUX2X1 U786 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1206), .Y(n616) );
  MUX2X1 U787 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1206), .Y(n620) );
  MUX2X1 U788 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1206), .Y(n619) );
  MUX2X1 U789 ( .B(n618), .A(n615), .S(n1172), .Y(n622) );
  MUX2X1 U790 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1206), .Y(n626) );
  MUX2X1 U791 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1206), .Y(n625) );
  MUX2X1 U792 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1206), .Y(n629) );
  MUX2X1 U793 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1206), .Y(n628) );
  MUX2X1 U794 ( .B(n627), .A(n624), .S(n1172), .Y(n638) );
  MUX2X1 U795 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1206), .Y(n632) );
  MUX2X1 U796 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1206), .Y(n631) );
  MUX2X1 U797 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1206), .Y(n635) );
  MUX2X1 U798 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1206), .Y(n634) );
  MUX2X1 U799 ( .B(n633), .A(n630), .S(n1172), .Y(n637) );
  MUX2X1 U800 ( .B(n636), .A(n621), .S(n1167), .Y(n1166) );
  INVX8 U801 ( .A(n1189), .Y(n1192) );
  INVX8 U802 ( .A(n1189), .Y(n1193) );
  INVX8 U803 ( .A(n1189), .Y(n1194) );
  INVX8 U804 ( .A(n1189), .Y(n1195) );
  INVX8 U805 ( .A(n1189), .Y(n1196) );
  INVX8 U806 ( .A(n1189), .Y(n1205) );
  INVX1 U807 ( .A(N11), .Y(n1311) );
  INVX1 U808 ( .A(N10), .Y(n1309) );
  INVX4 U809 ( .A(n1318), .Y(n1319) );
  INVX8 U810 ( .A(n1291), .Y(n1288) );
  INVX8 U811 ( .A(n1291), .Y(n1289) );
  INVX8 U812 ( .A(n1291), .Y(n1290) );
  INVX8 U813 ( .A(n17), .Y(n1291) );
  INVX8 U814 ( .A(n20), .Y(n1292) );
  INVX8 U815 ( .A(n21), .Y(n1293) );
  INVX8 U816 ( .A(n22), .Y(n1294) );
  INVX8 U817 ( .A(n23), .Y(n1295) );
  INVX8 U818 ( .A(n24), .Y(n1296) );
  INVX8 U819 ( .A(n25), .Y(n1297) );
  INVX8 U820 ( .A(n26), .Y(n1298) );
  INVX8 U821 ( .A(n27), .Y(n1299) );
  INVX8 U822 ( .A(n28), .Y(n1300) );
  INVX8 U823 ( .A(n29), .Y(n1301) );
  INVX8 U824 ( .A(n30), .Y(n1302) );
  INVX8 U825 ( .A(n1), .Y(n1303) );
  INVX8 U826 ( .A(n2), .Y(n1304) );
  INVX8 U827 ( .A(n3), .Y(n1305) );
  INVX8 U828 ( .A(n4), .Y(n1306) );
  INVX8 U829 ( .A(n5), .Y(n1307) );
  OR2X2 U830 ( .A(write), .B(rst), .Y(n1318) );
  AND2X2 U831 ( .A(N32), .B(n1319), .Y(\data_out<0> ) );
  AND2X2 U832 ( .A(N31), .B(n1319), .Y(\data_out<1> ) );
  AND2X2 U833 ( .A(N30), .B(n1319), .Y(\data_out<2> ) );
  AND2X2 U834 ( .A(N29), .B(n1319), .Y(\data_out<3> ) );
  AND2X2 U835 ( .A(N28), .B(n1319), .Y(\data_out<4> ) );
  AND2X2 U836 ( .A(N27), .B(n1319), .Y(\data_out<5> ) );
  AND2X2 U837 ( .A(N26), .B(n1319), .Y(\data_out<6> ) );
  AND2X2 U838 ( .A(N25), .B(n1319), .Y(\data_out<7> ) );
  AND2X2 U839 ( .A(N24), .B(n1319), .Y(\data_out<8> ) );
  AND2X2 U840 ( .A(N23), .B(n1319), .Y(\data_out<9> ) );
  AND2X2 U841 ( .A(N22), .B(n1319), .Y(\data_out<10> ) );
  AND2X2 U842 ( .A(N21), .B(n1319), .Y(\data_out<11> ) );
  AND2X2 U843 ( .A(N20), .B(n1319), .Y(\data_out<12> ) );
  AND2X2 U844 ( .A(N19), .B(n1319), .Y(\data_out<13> ) );
  AND2X2 U845 ( .A(N18), .B(n1319), .Y(\data_out<14> ) );
  AND2X2 U846 ( .A(N17), .B(n1319), .Y(\data_out<15> ) );
  NAND2X1 U847 ( .A(\mem<31><0> ), .B(n1209), .Y(n1320) );
  OAI21X1 U848 ( .A(n1208), .B(n1292), .C(n1320), .Y(n2358) );
  NAND2X1 U849 ( .A(\mem<31><1> ), .B(n1209), .Y(n1321) );
  OAI21X1 U850 ( .A(n1293), .B(n1208), .C(n1321), .Y(n2357) );
  NAND2X1 U851 ( .A(\mem<31><2> ), .B(n1209), .Y(n1322) );
  OAI21X1 U852 ( .A(n1294), .B(n1208), .C(n1322), .Y(n2356) );
  NAND2X1 U853 ( .A(\mem<31><3> ), .B(n1209), .Y(n1323) );
  OAI21X1 U854 ( .A(n1295), .B(n1208), .C(n1323), .Y(n2355) );
  NAND2X1 U855 ( .A(\mem<31><4> ), .B(n1209), .Y(n1324) );
  OAI21X1 U856 ( .A(n1296), .B(n1208), .C(n1324), .Y(n2354) );
  NAND2X1 U857 ( .A(\mem<31><5> ), .B(n1209), .Y(n1325) );
  OAI21X1 U858 ( .A(n1297), .B(n1208), .C(n1325), .Y(n2353) );
  NAND2X1 U859 ( .A(\mem<31><6> ), .B(n1209), .Y(n1326) );
  OAI21X1 U860 ( .A(n1298), .B(n1208), .C(n1326), .Y(n2352) );
  NAND2X1 U861 ( .A(\mem<31><7> ), .B(n1209), .Y(n1327) );
  OAI21X1 U862 ( .A(n1299), .B(n1208), .C(n1327), .Y(n2351) );
  NAND2X1 U863 ( .A(\mem<31><8> ), .B(n1210), .Y(n1328) );
  OAI21X1 U864 ( .A(n1300), .B(n1208), .C(n1328), .Y(n2350) );
  NAND2X1 U865 ( .A(\mem<31><9> ), .B(n1210), .Y(n1329) );
  OAI21X1 U866 ( .A(n1301), .B(n39), .C(n1329), .Y(n2349) );
  NAND2X1 U867 ( .A(\mem<31><10> ), .B(n1210), .Y(n1330) );
  OAI21X1 U868 ( .A(n1302), .B(n39), .C(n1330), .Y(n2348) );
  NAND2X1 U869 ( .A(\mem<31><11> ), .B(n1210), .Y(n1331) );
  OAI21X1 U870 ( .A(n1303), .B(n39), .C(n1331), .Y(n2347) );
  NAND2X1 U871 ( .A(\mem<31><12> ), .B(n1210), .Y(n1332) );
  OAI21X1 U872 ( .A(n1304), .B(n39), .C(n1332), .Y(n2346) );
  NAND2X1 U873 ( .A(\mem<31><13> ), .B(n1210), .Y(n1333) );
  OAI21X1 U874 ( .A(n1305), .B(n39), .C(n1333), .Y(n2345) );
  NAND2X1 U875 ( .A(\mem<31><14> ), .B(n1210), .Y(n1334) );
  OAI21X1 U876 ( .A(n1306), .B(n39), .C(n1334), .Y(n2344) );
  NAND2X1 U877 ( .A(\mem<31><15> ), .B(n1210), .Y(n1335) );
  OAI21X1 U878 ( .A(n1307), .B(n39), .C(n1335), .Y(n2343) );
  NAND2X1 U879 ( .A(\mem<30><0> ), .B(n1211), .Y(n1336) );
  OAI21X1 U880 ( .A(n43), .B(n1292), .C(n1336), .Y(n2342) );
  NAND2X1 U881 ( .A(\mem<30><1> ), .B(n1211), .Y(n1337) );
  OAI21X1 U882 ( .A(n43), .B(n1293), .C(n1337), .Y(n2341) );
  NAND2X1 U883 ( .A(\mem<30><2> ), .B(n1211), .Y(n1338) );
  OAI21X1 U884 ( .A(n43), .B(n1294), .C(n1338), .Y(n2340) );
  NAND2X1 U885 ( .A(\mem<30><3> ), .B(n1211), .Y(n1339) );
  OAI21X1 U886 ( .A(n43), .B(n1295), .C(n1339), .Y(n2339) );
  NAND2X1 U887 ( .A(\mem<30><4> ), .B(n1211), .Y(n1340) );
  OAI21X1 U888 ( .A(n43), .B(n1296), .C(n1340), .Y(n2338) );
  NAND2X1 U889 ( .A(\mem<30><5> ), .B(n1211), .Y(n1341) );
  OAI21X1 U890 ( .A(n43), .B(n1297), .C(n1341), .Y(n2337) );
  NAND2X1 U891 ( .A(\mem<30><6> ), .B(n1211), .Y(n1342) );
  OAI21X1 U892 ( .A(n43), .B(n1298), .C(n1342), .Y(n2336) );
  NAND2X1 U893 ( .A(\mem<30><7> ), .B(n1211), .Y(n1343) );
  OAI21X1 U894 ( .A(n43), .B(n1299), .C(n1343), .Y(n2335) );
  NAND2X1 U895 ( .A(\mem<30><8> ), .B(n1212), .Y(n1344) );
  OAI21X1 U896 ( .A(n43), .B(n1300), .C(n1344), .Y(n2334) );
  NAND2X1 U897 ( .A(\mem<30><9> ), .B(n1212), .Y(n1345) );
  OAI21X1 U898 ( .A(n43), .B(n1301), .C(n1345), .Y(n2333) );
  NAND2X1 U899 ( .A(\mem<30><10> ), .B(n1212), .Y(n1346) );
  OAI21X1 U900 ( .A(n43), .B(n1302), .C(n1346), .Y(n2332) );
  NAND2X1 U901 ( .A(\mem<30><11> ), .B(n1212), .Y(n1347) );
  OAI21X1 U902 ( .A(n43), .B(n1303), .C(n1347), .Y(n2331) );
  NAND2X1 U903 ( .A(\mem<30><12> ), .B(n1212), .Y(n1348) );
  OAI21X1 U904 ( .A(n43), .B(n1304), .C(n1348), .Y(n2330) );
  NAND2X1 U905 ( .A(\mem<30><13> ), .B(n1212), .Y(n1349) );
  OAI21X1 U906 ( .A(n43), .B(n1305), .C(n1349), .Y(n2329) );
  NAND2X1 U907 ( .A(\mem<30><14> ), .B(n1212), .Y(n1350) );
  OAI21X1 U908 ( .A(n43), .B(n1306), .C(n1350), .Y(n2328) );
  NAND2X1 U909 ( .A(\mem<30><15> ), .B(n1212), .Y(n1351) );
  OAI21X1 U910 ( .A(n43), .B(n1307), .C(n1351), .Y(n2327) );
  NAND3X1 U911 ( .A(n1308), .B(N12), .C(n1311), .Y(n1352) );
  NAND2X1 U912 ( .A(\mem<29><0> ), .B(n1214), .Y(n1353) );
  OAI21X1 U913 ( .A(n1213), .B(n1292), .C(n1353), .Y(n2326) );
  NAND2X1 U914 ( .A(\mem<29><1> ), .B(n1214), .Y(n1354) );
  OAI21X1 U915 ( .A(n1213), .B(n1293), .C(n1354), .Y(n2325) );
  NAND2X1 U916 ( .A(\mem<29><2> ), .B(n1214), .Y(n1355) );
  OAI21X1 U917 ( .A(n1213), .B(n1294), .C(n1355), .Y(n2324) );
  NAND2X1 U918 ( .A(\mem<29><3> ), .B(n1214), .Y(n1356) );
  OAI21X1 U919 ( .A(n1213), .B(n1295), .C(n1356), .Y(n2323) );
  NAND2X1 U920 ( .A(\mem<29><4> ), .B(n1214), .Y(n1357) );
  OAI21X1 U921 ( .A(n1213), .B(n1296), .C(n1357), .Y(n2322) );
  NAND2X1 U922 ( .A(\mem<29><5> ), .B(n1214), .Y(n1358) );
  OAI21X1 U923 ( .A(n1213), .B(n1297), .C(n1358), .Y(n2321) );
  NAND2X1 U924 ( .A(\mem<29><6> ), .B(n1214), .Y(n1359) );
  OAI21X1 U925 ( .A(n1213), .B(n1298), .C(n1359), .Y(n2320) );
  NAND2X1 U926 ( .A(\mem<29><7> ), .B(n1214), .Y(n1360) );
  OAI21X1 U927 ( .A(n1213), .B(n1299), .C(n1360), .Y(n2319) );
  NAND2X1 U928 ( .A(\mem<29><8> ), .B(n1215), .Y(n1361) );
  OAI21X1 U929 ( .A(n47), .B(n1300), .C(n1361), .Y(n2318) );
  NAND2X1 U930 ( .A(\mem<29><9> ), .B(n1215), .Y(n1362) );
  OAI21X1 U931 ( .A(n47), .B(n1301), .C(n1362), .Y(n2317) );
  NAND2X1 U932 ( .A(\mem<29><10> ), .B(n1215), .Y(n1363) );
  OAI21X1 U933 ( .A(n47), .B(n1302), .C(n1363), .Y(n2316) );
  NAND2X1 U934 ( .A(\mem<29><11> ), .B(n1215), .Y(n1364) );
  OAI21X1 U935 ( .A(n47), .B(n1303), .C(n1364), .Y(n2315) );
  NAND2X1 U936 ( .A(\mem<29><12> ), .B(n1215), .Y(n1365) );
  OAI21X1 U937 ( .A(n47), .B(n1304), .C(n1365), .Y(n2314) );
  NAND2X1 U938 ( .A(\mem<29><13> ), .B(n1215), .Y(n1366) );
  OAI21X1 U939 ( .A(n47), .B(n1305), .C(n1366), .Y(n2313) );
  NAND2X1 U940 ( .A(\mem<29><14> ), .B(n1215), .Y(n1367) );
  OAI21X1 U941 ( .A(n1213), .B(n1306), .C(n1367), .Y(n2312) );
  NAND2X1 U942 ( .A(\mem<29><15> ), .B(n1215), .Y(n1368) );
  OAI21X1 U943 ( .A(n1213), .B(n1307), .C(n1368), .Y(n2311) );
  NAND3X1 U944 ( .A(N12), .B(n1311), .C(n1309), .Y(n1369) );
  NAND2X1 U945 ( .A(\mem<28><0> ), .B(n1217), .Y(n1370) );
  OAI21X1 U946 ( .A(n1216), .B(n1292), .C(n1370), .Y(n2310) );
  NAND2X1 U947 ( .A(\mem<28><1> ), .B(n1217), .Y(n1371) );
  OAI21X1 U948 ( .A(n1216), .B(n1293), .C(n1371), .Y(n2309) );
  NAND2X1 U949 ( .A(\mem<28><2> ), .B(n1217), .Y(n1372) );
  OAI21X1 U950 ( .A(n1216), .B(n1294), .C(n1372), .Y(n2308) );
  NAND2X1 U951 ( .A(\mem<28><3> ), .B(n1217), .Y(n1373) );
  OAI21X1 U952 ( .A(n1216), .B(n1295), .C(n1373), .Y(n2307) );
  NAND2X1 U953 ( .A(\mem<28><4> ), .B(n1217), .Y(n1374) );
  OAI21X1 U954 ( .A(n1216), .B(n1296), .C(n1374), .Y(n2306) );
  NAND2X1 U955 ( .A(\mem<28><5> ), .B(n1217), .Y(n1375) );
  OAI21X1 U956 ( .A(n1216), .B(n1297), .C(n1375), .Y(n2305) );
  NAND2X1 U957 ( .A(\mem<28><6> ), .B(n1217), .Y(n1376) );
  OAI21X1 U958 ( .A(n1216), .B(n1298), .C(n1376), .Y(n2304) );
  NAND2X1 U959 ( .A(\mem<28><7> ), .B(n1217), .Y(n1377) );
  OAI21X1 U960 ( .A(n1216), .B(n1299), .C(n1377), .Y(n2303) );
  NAND2X1 U961 ( .A(\mem<28><8> ), .B(n1218), .Y(n1378) );
  OAI21X1 U962 ( .A(n51), .B(n1300), .C(n1378), .Y(n2302) );
  NAND2X1 U963 ( .A(\mem<28><9> ), .B(n1218), .Y(n1379) );
  OAI21X1 U964 ( .A(n51), .B(n1301), .C(n1379), .Y(n2301) );
  NAND2X1 U965 ( .A(\mem<28><10> ), .B(n1218), .Y(n1380) );
  OAI21X1 U966 ( .A(n51), .B(n1302), .C(n1380), .Y(n2300) );
  NAND2X1 U967 ( .A(\mem<28><11> ), .B(n1218), .Y(n1381) );
  OAI21X1 U968 ( .A(n51), .B(n1303), .C(n1381), .Y(n2299) );
  NAND2X1 U969 ( .A(\mem<28><12> ), .B(n1218), .Y(n1382) );
  OAI21X1 U970 ( .A(n51), .B(n1304), .C(n1382), .Y(n2298) );
  NAND2X1 U971 ( .A(\mem<28><13> ), .B(n1218), .Y(n1383) );
  OAI21X1 U972 ( .A(n51), .B(n1305), .C(n1383), .Y(n2297) );
  NAND2X1 U973 ( .A(\mem<28><14> ), .B(n1218), .Y(n1384) );
  OAI21X1 U974 ( .A(n1216), .B(n1306), .C(n1384), .Y(n2296) );
  NAND2X1 U975 ( .A(\mem<28><15> ), .B(n1218), .Y(n1385) );
  OAI21X1 U976 ( .A(n1216), .B(n1307), .C(n1385), .Y(n2295) );
  NAND3X1 U977 ( .A(n1308), .B(n1310), .C(n1312), .Y(n1386) );
  NAND2X1 U978 ( .A(\mem<27><0> ), .B(n1219), .Y(n1387) );
  OAI21X1 U979 ( .A(n55), .B(n1292), .C(n1387), .Y(n2294) );
  NAND2X1 U980 ( .A(\mem<27><1> ), .B(n1219), .Y(n1388) );
  OAI21X1 U981 ( .A(n55), .B(n1293), .C(n1388), .Y(n2293) );
  NAND2X1 U982 ( .A(\mem<27><2> ), .B(n1219), .Y(n1389) );
  OAI21X1 U983 ( .A(n55), .B(n1294), .C(n1389), .Y(n2292) );
  NAND2X1 U984 ( .A(\mem<27><3> ), .B(n1219), .Y(n1390) );
  OAI21X1 U985 ( .A(n55), .B(n1295), .C(n1390), .Y(n2291) );
  NAND2X1 U986 ( .A(\mem<27><4> ), .B(n1219), .Y(n1391) );
  OAI21X1 U987 ( .A(n55), .B(n1296), .C(n1391), .Y(n2290) );
  NAND2X1 U988 ( .A(\mem<27><5> ), .B(n1219), .Y(n1392) );
  OAI21X1 U989 ( .A(n55), .B(n1297), .C(n1392), .Y(n2289) );
  NAND2X1 U990 ( .A(\mem<27><6> ), .B(n1219), .Y(n1393) );
  OAI21X1 U991 ( .A(n55), .B(n1298), .C(n1393), .Y(n2288) );
  NAND2X1 U992 ( .A(\mem<27><7> ), .B(n1219), .Y(n1394) );
  OAI21X1 U993 ( .A(n55), .B(n1299), .C(n1394), .Y(n2287) );
  NAND2X1 U994 ( .A(\mem<27><8> ), .B(n1220), .Y(n1395) );
  OAI21X1 U995 ( .A(n55), .B(n1300), .C(n1395), .Y(n2286) );
  NAND2X1 U996 ( .A(\mem<27><9> ), .B(n1220), .Y(n1396) );
  OAI21X1 U997 ( .A(n55), .B(n1301), .C(n1396), .Y(n2285) );
  NAND2X1 U998 ( .A(\mem<27><10> ), .B(n1220), .Y(n1397) );
  OAI21X1 U999 ( .A(n55), .B(n1302), .C(n1397), .Y(n2284) );
  NAND2X1 U1000 ( .A(\mem<27><11> ), .B(n1220), .Y(n1398) );
  OAI21X1 U1001 ( .A(n55), .B(n1303), .C(n1398), .Y(n2283) );
  NAND2X1 U1002 ( .A(\mem<27><12> ), .B(n1220), .Y(n1399) );
  OAI21X1 U1003 ( .A(n55), .B(n1304), .C(n1399), .Y(n2282) );
  NAND2X1 U1004 ( .A(\mem<27><13> ), .B(n1220), .Y(n1400) );
  OAI21X1 U1005 ( .A(n55), .B(n1305), .C(n1400), .Y(n2281) );
  NAND2X1 U1006 ( .A(\mem<27><14> ), .B(n1220), .Y(n1401) );
  OAI21X1 U1007 ( .A(n55), .B(n1306), .C(n1401), .Y(n2280) );
  NAND2X1 U1008 ( .A(\mem<27><15> ), .B(n1220), .Y(n1402) );
  OAI21X1 U1009 ( .A(n55), .B(n1307), .C(n1402), .Y(n2279) );
  NAND3X1 U1010 ( .A(n1312), .B(n1310), .C(n1309), .Y(n1403) );
  NAND2X1 U1011 ( .A(\mem<26><0> ), .B(n1221), .Y(n1404) );
  OAI21X1 U1012 ( .A(n59), .B(n1292), .C(n1404), .Y(n2278) );
  NAND2X1 U1013 ( .A(\mem<26><1> ), .B(n1221), .Y(n1405) );
  OAI21X1 U1014 ( .A(n59), .B(n1293), .C(n1405), .Y(n2277) );
  NAND2X1 U1015 ( .A(\mem<26><2> ), .B(n1221), .Y(n1406) );
  OAI21X1 U1016 ( .A(n59), .B(n1294), .C(n1406), .Y(n2276) );
  NAND2X1 U1017 ( .A(\mem<26><3> ), .B(n1221), .Y(n1407) );
  OAI21X1 U1018 ( .A(n59), .B(n1295), .C(n1407), .Y(n2275) );
  NAND2X1 U1019 ( .A(\mem<26><4> ), .B(n1221), .Y(n1408) );
  OAI21X1 U1020 ( .A(n59), .B(n1296), .C(n1408), .Y(n2274) );
  NAND2X1 U1021 ( .A(\mem<26><5> ), .B(n1221), .Y(n1409) );
  OAI21X1 U1022 ( .A(n59), .B(n1297), .C(n1409), .Y(n2273) );
  NAND2X1 U1023 ( .A(\mem<26><6> ), .B(n1221), .Y(n1410) );
  OAI21X1 U1024 ( .A(n59), .B(n1298), .C(n1410), .Y(n2272) );
  NAND2X1 U1025 ( .A(\mem<26><7> ), .B(n1221), .Y(n1411) );
  OAI21X1 U1026 ( .A(n59), .B(n1299), .C(n1411), .Y(n2271) );
  NAND2X1 U1027 ( .A(\mem<26><8> ), .B(n1222), .Y(n1412) );
  OAI21X1 U1028 ( .A(n59), .B(n1300), .C(n1412), .Y(n2270) );
  NAND2X1 U1029 ( .A(\mem<26><9> ), .B(n1222), .Y(n1413) );
  OAI21X1 U1030 ( .A(n59), .B(n1301), .C(n1413), .Y(n2269) );
  NAND2X1 U1031 ( .A(\mem<26><10> ), .B(n1222), .Y(n1414) );
  OAI21X1 U1032 ( .A(n59), .B(n1302), .C(n1414), .Y(n2268) );
  NAND2X1 U1033 ( .A(\mem<26><11> ), .B(n1222), .Y(n1415) );
  OAI21X1 U1034 ( .A(n59), .B(n1303), .C(n1415), .Y(n2267) );
  NAND2X1 U1035 ( .A(\mem<26><12> ), .B(n1222), .Y(n1416) );
  OAI21X1 U1036 ( .A(n59), .B(n1304), .C(n1416), .Y(n2266) );
  NAND2X1 U1037 ( .A(\mem<26><13> ), .B(n1222), .Y(n1417) );
  OAI21X1 U1038 ( .A(n59), .B(n1305), .C(n1417), .Y(n2265) );
  NAND2X1 U1039 ( .A(\mem<26><14> ), .B(n1222), .Y(n1418) );
  OAI21X1 U1040 ( .A(n59), .B(n1306), .C(n1418), .Y(n2264) );
  NAND2X1 U1041 ( .A(\mem<26><15> ), .B(n1222), .Y(n1419) );
  OAI21X1 U1042 ( .A(n59), .B(n1307), .C(n1419), .Y(n2263) );
  NAND3X1 U1043 ( .A(n1308), .B(n1312), .C(n1311), .Y(n1420) );
  NAND2X1 U1044 ( .A(\mem<25><0> ), .B(n1223), .Y(n1421) );
  OAI21X1 U1045 ( .A(n63), .B(n1292), .C(n1421), .Y(n2262) );
  NAND2X1 U1046 ( .A(\mem<25><1> ), .B(n1223), .Y(n1422) );
  OAI21X1 U1047 ( .A(n63), .B(n1293), .C(n1422), .Y(n2261) );
  NAND2X1 U1048 ( .A(\mem<25><2> ), .B(n1223), .Y(n1423) );
  OAI21X1 U1049 ( .A(n63), .B(n1294), .C(n1423), .Y(n2260) );
  NAND2X1 U1050 ( .A(\mem<25><3> ), .B(n1223), .Y(n1424) );
  OAI21X1 U1051 ( .A(n63), .B(n1295), .C(n1424), .Y(n2259) );
  NAND2X1 U1052 ( .A(\mem<25><4> ), .B(n1223), .Y(n1425) );
  OAI21X1 U1053 ( .A(n63), .B(n1296), .C(n1425), .Y(n2258) );
  NAND2X1 U1054 ( .A(\mem<25><5> ), .B(n1223), .Y(n1426) );
  OAI21X1 U1055 ( .A(n63), .B(n1297), .C(n1426), .Y(n2257) );
  NAND2X1 U1056 ( .A(\mem<25><6> ), .B(n1223), .Y(n1427) );
  OAI21X1 U1057 ( .A(n63), .B(n1298), .C(n1427), .Y(n2256) );
  NAND2X1 U1058 ( .A(\mem<25><7> ), .B(n1223), .Y(n1428) );
  OAI21X1 U1059 ( .A(n63), .B(n1299), .C(n1428), .Y(n2255) );
  NAND2X1 U1060 ( .A(\mem<25><8> ), .B(n1224), .Y(n1429) );
  OAI21X1 U1061 ( .A(n63), .B(n1300), .C(n1429), .Y(n2254) );
  NAND2X1 U1062 ( .A(\mem<25><9> ), .B(n1224), .Y(n1430) );
  OAI21X1 U1063 ( .A(n63), .B(n1301), .C(n1430), .Y(n2253) );
  NAND2X1 U1064 ( .A(\mem<25><10> ), .B(n1224), .Y(n1431) );
  OAI21X1 U1065 ( .A(n63), .B(n1302), .C(n1431), .Y(n2252) );
  NAND2X1 U1066 ( .A(\mem<25><11> ), .B(n1224), .Y(n1432) );
  OAI21X1 U1067 ( .A(n63), .B(n1303), .C(n1432), .Y(n2251) );
  NAND2X1 U1068 ( .A(\mem<25><12> ), .B(n1224), .Y(n1433) );
  OAI21X1 U1069 ( .A(n63), .B(n1304), .C(n1433), .Y(n2250) );
  NAND2X1 U1070 ( .A(\mem<25><13> ), .B(n1224), .Y(n1434) );
  OAI21X1 U1071 ( .A(n63), .B(n1305), .C(n1434), .Y(n2249) );
  NAND2X1 U1072 ( .A(\mem<25><14> ), .B(n1224), .Y(n1435) );
  OAI21X1 U1073 ( .A(n63), .B(n1306), .C(n1435), .Y(n2248) );
  NAND2X1 U1074 ( .A(\mem<25><15> ), .B(n1224), .Y(n1436) );
  OAI21X1 U1075 ( .A(n63), .B(n1307), .C(n1436), .Y(n2247) );
  NOR3X1 U1076 ( .A(n1308), .B(n1310), .C(n1174), .Y(n1830) );
  NAND2X1 U1077 ( .A(\mem<24><0> ), .B(n1225), .Y(n1437) );
  OAI21X1 U1078 ( .A(n32), .B(n1292), .C(n1437), .Y(n2246) );
  NAND2X1 U1079 ( .A(\mem<24><1> ), .B(n1225), .Y(n1438) );
  OAI21X1 U1080 ( .A(n32), .B(n1293), .C(n1438), .Y(n2245) );
  NAND2X1 U1081 ( .A(\mem<24><2> ), .B(n1225), .Y(n1439) );
  OAI21X1 U1082 ( .A(n32), .B(n1294), .C(n1439), .Y(n2244) );
  NAND2X1 U1083 ( .A(\mem<24><3> ), .B(n1225), .Y(n1440) );
  OAI21X1 U1084 ( .A(n32), .B(n1295), .C(n1440), .Y(n2243) );
  NAND2X1 U1085 ( .A(\mem<24><4> ), .B(n1225), .Y(n1441) );
  OAI21X1 U1086 ( .A(n32), .B(n1296), .C(n1441), .Y(n2242) );
  NAND2X1 U1087 ( .A(\mem<24><5> ), .B(n1225), .Y(n1442) );
  OAI21X1 U1088 ( .A(n32), .B(n1297), .C(n1442), .Y(n2241) );
  NAND2X1 U1089 ( .A(\mem<24><6> ), .B(n1225), .Y(n1443) );
  OAI21X1 U1090 ( .A(n32), .B(n1298), .C(n1443), .Y(n2240) );
  NAND2X1 U1091 ( .A(\mem<24><7> ), .B(n1225), .Y(n1444) );
  OAI21X1 U1092 ( .A(n32), .B(n1299), .C(n1444), .Y(n2239) );
  NAND2X1 U1093 ( .A(\mem<24><8> ), .B(n1226), .Y(n1445) );
  OAI21X1 U1094 ( .A(n32), .B(n1300), .C(n1445), .Y(n2238) );
  NAND2X1 U1095 ( .A(\mem<24><9> ), .B(n1226), .Y(n1446) );
  OAI21X1 U1096 ( .A(n32), .B(n1301), .C(n1446), .Y(n2237) );
  NAND2X1 U1097 ( .A(\mem<24><10> ), .B(n1226), .Y(n1447) );
  OAI21X1 U1098 ( .A(n32), .B(n1302), .C(n1447), .Y(n2236) );
  NAND2X1 U1099 ( .A(\mem<24><11> ), .B(n1226), .Y(n1448) );
  OAI21X1 U1100 ( .A(n32), .B(n1303), .C(n1448), .Y(n2235) );
  NAND2X1 U1101 ( .A(\mem<24><12> ), .B(n1226), .Y(n1449) );
  OAI21X1 U1102 ( .A(n32), .B(n1304), .C(n1449), .Y(n2234) );
  NAND2X1 U1103 ( .A(\mem<24><13> ), .B(n1226), .Y(n1450) );
  OAI21X1 U1104 ( .A(n32), .B(n1305), .C(n1450), .Y(n2233) );
  NAND2X1 U1105 ( .A(\mem<24><14> ), .B(n1226), .Y(n1451) );
  OAI21X1 U1106 ( .A(n32), .B(n1306), .C(n1451), .Y(n2232) );
  NAND2X1 U1107 ( .A(\mem<24><15> ), .B(n1226), .Y(n1452) );
  OAI21X1 U1108 ( .A(n32), .B(n1307), .C(n1452), .Y(n2231) );
  NAND2X1 U1109 ( .A(\mem<23><0> ), .B(n1229), .Y(n1453) );
  OAI21X1 U1110 ( .A(n1227), .B(n1292), .C(n1453), .Y(n2230) );
  NAND2X1 U1111 ( .A(\mem<23><1> ), .B(n1229), .Y(n1454) );
  OAI21X1 U1112 ( .A(n1227), .B(n1293), .C(n1454), .Y(n2229) );
  NAND2X1 U1113 ( .A(\mem<23><2> ), .B(n1229), .Y(n1455) );
  OAI21X1 U1114 ( .A(n1227), .B(n1294), .C(n1455), .Y(n2228) );
  NAND2X1 U1115 ( .A(\mem<23><3> ), .B(n1229), .Y(n1456) );
  OAI21X1 U1116 ( .A(n1227), .B(n1295), .C(n1456), .Y(n2227) );
  NAND2X1 U1117 ( .A(\mem<23><4> ), .B(n1229), .Y(n1457) );
  OAI21X1 U1118 ( .A(n1227), .B(n1296), .C(n1457), .Y(n2226) );
  NAND2X1 U1119 ( .A(\mem<23><5> ), .B(n1229), .Y(n1458) );
  OAI21X1 U1120 ( .A(n1227), .B(n1297), .C(n1458), .Y(n2225) );
  NAND2X1 U1121 ( .A(\mem<23><6> ), .B(n1229), .Y(n1459) );
  OAI21X1 U1122 ( .A(n1227), .B(n1298), .C(n1459), .Y(n2224) );
  NAND2X1 U1123 ( .A(\mem<23><7> ), .B(n1229), .Y(n1460) );
  OAI21X1 U1124 ( .A(n1227), .B(n1299), .C(n1460), .Y(n2223) );
  NAND2X1 U1125 ( .A(\mem<23><8> ), .B(n1230), .Y(n1461) );
  OAI21X1 U1126 ( .A(n1228), .B(n1300), .C(n1461), .Y(n2222) );
  NAND2X1 U1127 ( .A(\mem<23><9> ), .B(n1230), .Y(n1462) );
  OAI21X1 U1128 ( .A(n1228), .B(n1301), .C(n1462), .Y(n2221) );
  NAND2X1 U1129 ( .A(\mem<23><10> ), .B(n1230), .Y(n1463) );
  OAI21X1 U1130 ( .A(n1228), .B(n1302), .C(n1463), .Y(n2220) );
  NAND2X1 U1131 ( .A(\mem<23><11> ), .B(n1230), .Y(n1464) );
  OAI21X1 U1132 ( .A(n1228), .B(n1303), .C(n1464), .Y(n2219) );
  NAND2X1 U1133 ( .A(\mem<23><12> ), .B(n1230), .Y(n1465) );
  OAI21X1 U1134 ( .A(n1228), .B(n1304), .C(n1465), .Y(n2218) );
  NAND2X1 U1135 ( .A(\mem<23><13> ), .B(n1230), .Y(n1466) );
  OAI21X1 U1136 ( .A(n1228), .B(n1305), .C(n1466), .Y(n2217) );
  NAND2X1 U1137 ( .A(\mem<23><14> ), .B(n1230), .Y(n1467) );
  OAI21X1 U1138 ( .A(n1228), .B(n1306), .C(n1467), .Y(n2216) );
  NAND2X1 U1139 ( .A(\mem<23><15> ), .B(n1230), .Y(n1468) );
  OAI21X1 U1140 ( .A(n1228), .B(n1307), .C(n1468), .Y(n2215) );
  NAND2X1 U1141 ( .A(\mem<22><0> ), .B(n1231), .Y(n1469) );
  OAI21X1 U1142 ( .A(n73), .B(n1292), .C(n1469), .Y(n2214) );
  NAND2X1 U1143 ( .A(\mem<22><1> ), .B(n1231), .Y(n1470) );
  OAI21X1 U1144 ( .A(n73), .B(n1293), .C(n1470), .Y(n2213) );
  NAND2X1 U1145 ( .A(\mem<22><2> ), .B(n1231), .Y(n1471) );
  OAI21X1 U1146 ( .A(n73), .B(n1294), .C(n1471), .Y(n2212) );
  NAND2X1 U1147 ( .A(\mem<22><3> ), .B(n1231), .Y(n1472) );
  OAI21X1 U1148 ( .A(n73), .B(n1295), .C(n1472), .Y(n2211) );
  NAND2X1 U1149 ( .A(\mem<22><4> ), .B(n1231), .Y(n1473) );
  OAI21X1 U1150 ( .A(n73), .B(n1296), .C(n1473), .Y(n2210) );
  NAND2X1 U1151 ( .A(\mem<22><5> ), .B(n1231), .Y(n1474) );
  OAI21X1 U1152 ( .A(n73), .B(n1297), .C(n1474), .Y(n2209) );
  NAND2X1 U1153 ( .A(\mem<22><6> ), .B(n1231), .Y(n1475) );
  OAI21X1 U1154 ( .A(n73), .B(n1298), .C(n1475), .Y(n2208) );
  NAND2X1 U1155 ( .A(\mem<22><7> ), .B(n1231), .Y(n1476) );
  OAI21X1 U1156 ( .A(n73), .B(n1299), .C(n1476), .Y(n2207) );
  NAND2X1 U1157 ( .A(\mem<22><8> ), .B(n1232), .Y(n1477) );
  OAI21X1 U1158 ( .A(n73), .B(n1300), .C(n1477), .Y(n2206) );
  NAND2X1 U1159 ( .A(\mem<22><9> ), .B(n1232), .Y(n1478) );
  OAI21X1 U1160 ( .A(n73), .B(n1301), .C(n1478), .Y(n2205) );
  NAND2X1 U1161 ( .A(\mem<22><10> ), .B(n1232), .Y(n1479) );
  OAI21X1 U1162 ( .A(n73), .B(n1302), .C(n1479), .Y(n2204) );
  NAND2X1 U1163 ( .A(\mem<22><11> ), .B(n1232), .Y(n1480) );
  OAI21X1 U1164 ( .A(n73), .B(n1303), .C(n1480), .Y(n2203) );
  NAND2X1 U1165 ( .A(\mem<22><12> ), .B(n1232), .Y(n1481) );
  OAI21X1 U1166 ( .A(n73), .B(n1304), .C(n1481), .Y(n2202) );
  NAND2X1 U1167 ( .A(\mem<22><13> ), .B(n1232), .Y(n1482) );
  OAI21X1 U1168 ( .A(n73), .B(n1305), .C(n1482), .Y(n2201) );
  NAND2X1 U1169 ( .A(\mem<22><14> ), .B(n1232), .Y(n1483) );
  OAI21X1 U1170 ( .A(n73), .B(n1306), .C(n1483), .Y(n2200) );
  NAND2X1 U1171 ( .A(\mem<22><15> ), .B(n1232), .Y(n1484) );
  OAI21X1 U1172 ( .A(n73), .B(n1307), .C(n1484), .Y(n2199) );
  NAND2X1 U1173 ( .A(\mem<21><0> ), .B(n1234), .Y(n1485) );
  OAI21X1 U1174 ( .A(n1233), .B(n1292), .C(n1485), .Y(n2198) );
  NAND2X1 U1175 ( .A(\mem<21><1> ), .B(n1234), .Y(n1486) );
  OAI21X1 U1177 ( .A(n1233), .B(n1293), .C(n1486), .Y(n2197) );
  NAND2X1 U1178 ( .A(\mem<21><2> ), .B(n1234), .Y(n1487) );
  OAI21X1 U1179 ( .A(n1233), .B(n1294), .C(n1487), .Y(n2196) );
  NAND2X1 U1180 ( .A(\mem<21><3> ), .B(n1234), .Y(n1488) );
  OAI21X1 U1181 ( .A(n1233), .B(n1295), .C(n1488), .Y(n2195) );
  NAND2X1 U1182 ( .A(\mem<21><4> ), .B(n1234), .Y(n1489) );
  OAI21X1 U1183 ( .A(n1233), .B(n1296), .C(n1489), .Y(n2194) );
  NAND2X1 U1184 ( .A(\mem<21><5> ), .B(n1234), .Y(n1490) );
  OAI21X1 U1185 ( .A(n1233), .B(n1297), .C(n1490), .Y(n2193) );
  NAND2X1 U1186 ( .A(\mem<21><6> ), .B(n1234), .Y(n1491) );
  OAI21X1 U1187 ( .A(n1233), .B(n1298), .C(n1491), .Y(n2192) );
  NAND2X1 U1188 ( .A(\mem<21><7> ), .B(n1234), .Y(n1492) );
  OAI21X1 U1189 ( .A(n1233), .B(n1299), .C(n1492), .Y(n2191) );
  NAND2X1 U1190 ( .A(\mem<21><8> ), .B(n1235), .Y(n1493) );
  OAI21X1 U1191 ( .A(n77), .B(n1300), .C(n1493), .Y(n2190) );
  NAND2X1 U1192 ( .A(\mem<21><9> ), .B(n1235), .Y(n1494) );
  OAI21X1 U1193 ( .A(n77), .B(n1301), .C(n1494), .Y(n2189) );
  NAND2X1 U1194 ( .A(\mem<21><10> ), .B(n1235), .Y(n1495) );
  OAI21X1 U1195 ( .A(n77), .B(n1302), .C(n1495), .Y(n2188) );
  NAND2X1 U1196 ( .A(\mem<21><11> ), .B(n1235), .Y(n1496) );
  OAI21X1 U1197 ( .A(n77), .B(n1303), .C(n1496), .Y(n2187) );
  NAND2X1 U1198 ( .A(\mem<21><12> ), .B(n1235), .Y(n1497) );
  OAI21X1 U1199 ( .A(n77), .B(n1304), .C(n1497), .Y(n2186) );
  NAND2X1 U1200 ( .A(\mem<21><13> ), .B(n1235), .Y(n1498) );
  OAI21X1 U1201 ( .A(n77), .B(n1305), .C(n1498), .Y(n2185) );
  NAND2X1 U1202 ( .A(\mem<21><14> ), .B(n1235), .Y(n1499) );
  OAI21X1 U1203 ( .A(n1233), .B(n1306), .C(n1499), .Y(n2184) );
  NAND2X1 U1204 ( .A(\mem<21><15> ), .B(n1235), .Y(n1500) );
  OAI21X1 U1205 ( .A(n1233), .B(n1307), .C(n1500), .Y(n2183) );
  NAND2X1 U1206 ( .A(\mem<20><0> ), .B(n1237), .Y(n1501) );
  OAI21X1 U1207 ( .A(n1236), .B(n1292), .C(n1501), .Y(n2182) );
  NAND2X1 U1208 ( .A(\mem<20><1> ), .B(n1237), .Y(n1502) );
  OAI21X1 U1209 ( .A(n1236), .B(n1293), .C(n1502), .Y(n2181) );
  NAND2X1 U1210 ( .A(\mem<20><2> ), .B(n1237), .Y(n1503) );
  OAI21X1 U1211 ( .A(n1236), .B(n1294), .C(n1503), .Y(n2180) );
  NAND2X1 U1212 ( .A(\mem<20><3> ), .B(n1237), .Y(n1504) );
  OAI21X1 U1213 ( .A(n1236), .B(n1295), .C(n1504), .Y(n2179) );
  NAND2X1 U1214 ( .A(\mem<20><4> ), .B(n1237), .Y(n1505) );
  OAI21X1 U1215 ( .A(n1236), .B(n1296), .C(n1505), .Y(n2178) );
  NAND2X1 U1216 ( .A(\mem<20><5> ), .B(n1237), .Y(n1506) );
  OAI21X1 U1217 ( .A(n1236), .B(n1297), .C(n1506), .Y(n2177) );
  NAND2X1 U1218 ( .A(\mem<20><6> ), .B(n1237), .Y(n1507) );
  OAI21X1 U1219 ( .A(n1236), .B(n1298), .C(n1507), .Y(n2176) );
  NAND2X1 U1220 ( .A(\mem<20><7> ), .B(n1237), .Y(n1508) );
  OAI21X1 U1221 ( .A(n1236), .B(n1299), .C(n1508), .Y(n2175) );
  NAND2X1 U1222 ( .A(\mem<20><8> ), .B(n1238), .Y(n1509) );
  OAI21X1 U1223 ( .A(n81), .B(n1300), .C(n1509), .Y(n2174) );
  NAND2X1 U1224 ( .A(\mem<20><9> ), .B(n1238), .Y(n1510) );
  OAI21X1 U1225 ( .A(n81), .B(n1301), .C(n1510), .Y(n2173) );
  NAND2X1 U1226 ( .A(\mem<20><10> ), .B(n1238), .Y(n1511) );
  OAI21X1 U1227 ( .A(n81), .B(n1302), .C(n1511), .Y(n2172) );
  NAND2X1 U1228 ( .A(\mem<20><11> ), .B(n1238), .Y(n1512) );
  OAI21X1 U1229 ( .A(n81), .B(n1303), .C(n1512), .Y(n2171) );
  NAND2X1 U1230 ( .A(\mem<20><12> ), .B(n1238), .Y(n1513) );
  OAI21X1 U1231 ( .A(n81), .B(n1304), .C(n1513), .Y(n2170) );
  NAND2X1 U1232 ( .A(\mem<20><13> ), .B(n1238), .Y(n1514) );
  OAI21X1 U1233 ( .A(n81), .B(n1305), .C(n1514), .Y(n2169) );
  NAND2X1 U1234 ( .A(\mem<20><14> ), .B(n1238), .Y(n1515) );
  OAI21X1 U1235 ( .A(n1236), .B(n1306), .C(n1515), .Y(n2168) );
  NAND2X1 U1236 ( .A(\mem<20><15> ), .B(n1238), .Y(n1516) );
  OAI21X1 U1237 ( .A(n1236), .B(n1307), .C(n1516), .Y(n2167) );
  NAND2X1 U1238 ( .A(\mem<19><0> ), .B(n1239), .Y(n1517) );
  OAI21X1 U1239 ( .A(n85), .B(n1292), .C(n1517), .Y(n2166) );
  NAND2X1 U1240 ( .A(\mem<19><1> ), .B(n1239), .Y(n1518) );
  OAI21X1 U1241 ( .A(n85), .B(n1293), .C(n1518), .Y(n2165) );
  NAND2X1 U1242 ( .A(\mem<19><2> ), .B(n1239), .Y(n1519) );
  OAI21X1 U1243 ( .A(n85), .B(n1294), .C(n1519), .Y(n2164) );
  NAND2X1 U1244 ( .A(\mem<19><3> ), .B(n1239), .Y(n1520) );
  OAI21X1 U1245 ( .A(n85), .B(n1295), .C(n1520), .Y(n2163) );
  NAND2X1 U1246 ( .A(\mem<19><4> ), .B(n1239), .Y(n1521) );
  OAI21X1 U1247 ( .A(n85), .B(n1296), .C(n1521), .Y(n2162) );
  NAND2X1 U1248 ( .A(\mem<19><5> ), .B(n1239), .Y(n1522) );
  OAI21X1 U1249 ( .A(n85), .B(n1297), .C(n1522), .Y(n2161) );
  NAND2X1 U1250 ( .A(\mem<19><6> ), .B(n1239), .Y(n1523) );
  OAI21X1 U1251 ( .A(n85), .B(n1298), .C(n1523), .Y(n2160) );
  NAND2X1 U1252 ( .A(\mem<19><7> ), .B(n1239), .Y(n1524) );
  OAI21X1 U1253 ( .A(n85), .B(n1299), .C(n1524), .Y(n2159) );
  NAND2X1 U1254 ( .A(\mem<19><8> ), .B(n1240), .Y(n1525) );
  OAI21X1 U1255 ( .A(n85), .B(n1300), .C(n1525), .Y(n2158) );
  NAND2X1 U1256 ( .A(\mem<19><9> ), .B(n1240), .Y(n1526) );
  OAI21X1 U1257 ( .A(n85), .B(n1301), .C(n1526), .Y(n2157) );
  NAND2X1 U1258 ( .A(\mem<19><10> ), .B(n1240), .Y(n1527) );
  OAI21X1 U1259 ( .A(n85), .B(n1302), .C(n1527), .Y(n2156) );
  NAND2X1 U1260 ( .A(\mem<19><11> ), .B(n1240), .Y(n1528) );
  OAI21X1 U1261 ( .A(n85), .B(n1303), .C(n1528), .Y(n2155) );
  NAND2X1 U1262 ( .A(\mem<19><12> ), .B(n1240), .Y(n1529) );
  OAI21X1 U1263 ( .A(n85), .B(n1304), .C(n1529), .Y(n2154) );
  NAND2X1 U1264 ( .A(\mem<19><13> ), .B(n1240), .Y(n1530) );
  OAI21X1 U1265 ( .A(n85), .B(n1305), .C(n1530), .Y(n2153) );
  NAND2X1 U1266 ( .A(\mem<19><14> ), .B(n1240), .Y(n1531) );
  OAI21X1 U1267 ( .A(n85), .B(n1306), .C(n1531), .Y(n2152) );
  NAND2X1 U1268 ( .A(\mem<19><15> ), .B(n1240), .Y(n1532) );
  OAI21X1 U1269 ( .A(n85), .B(n1307), .C(n1532), .Y(n2151) );
  NAND2X1 U1270 ( .A(\mem<18><0> ), .B(n1241), .Y(n1533) );
  OAI21X1 U1271 ( .A(n89), .B(n1292), .C(n1533), .Y(n2150) );
  NAND2X1 U1272 ( .A(\mem<18><1> ), .B(n1241), .Y(n1534) );
  OAI21X1 U1273 ( .A(n89), .B(n1293), .C(n1534), .Y(n2149) );
  NAND2X1 U1274 ( .A(\mem<18><2> ), .B(n1241), .Y(n1535) );
  OAI21X1 U1275 ( .A(n89), .B(n1294), .C(n1535), .Y(n2148) );
  NAND2X1 U1276 ( .A(\mem<18><3> ), .B(n1241), .Y(n1536) );
  OAI21X1 U1277 ( .A(n89), .B(n1295), .C(n1536), .Y(n2147) );
  NAND2X1 U1278 ( .A(\mem<18><4> ), .B(n1241), .Y(n1537) );
  OAI21X1 U1279 ( .A(n89), .B(n1296), .C(n1537), .Y(n2146) );
  NAND2X1 U1280 ( .A(\mem<18><5> ), .B(n1241), .Y(n1538) );
  OAI21X1 U1281 ( .A(n89), .B(n1297), .C(n1538), .Y(n2145) );
  NAND2X1 U1282 ( .A(\mem<18><6> ), .B(n1241), .Y(n1539) );
  OAI21X1 U1283 ( .A(n89), .B(n1298), .C(n1539), .Y(n2144) );
  NAND2X1 U1284 ( .A(\mem<18><7> ), .B(n1241), .Y(n1540) );
  OAI21X1 U1285 ( .A(n89), .B(n1299), .C(n1540), .Y(n2143) );
  NAND2X1 U1286 ( .A(\mem<18><8> ), .B(n1242), .Y(n1541) );
  OAI21X1 U1287 ( .A(n89), .B(n1300), .C(n1541), .Y(n2142) );
  NAND2X1 U1288 ( .A(\mem<18><9> ), .B(n1242), .Y(n1542) );
  OAI21X1 U1289 ( .A(n89), .B(n1301), .C(n1542), .Y(n2141) );
  NAND2X1 U1290 ( .A(\mem<18><10> ), .B(n1242), .Y(n1543) );
  OAI21X1 U1291 ( .A(n89), .B(n1302), .C(n1543), .Y(n2140) );
  NAND2X1 U1292 ( .A(\mem<18><11> ), .B(n1242), .Y(n1544) );
  OAI21X1 U1293 ( .A(n89), .B(n1303), .C(n1544), .Y(n2139) );
  NAND2X1 U1294 ( .A(\mem<18><12> ), .B(n1242), .Y(n1545) );
  OAI21X1 U1295 ( .A(n89), .B(n1304), .C(n1545), .Y(n2138) );
  NAND2X1 U1296 ( .A(\mem<18><13> ), .B(n1242), .Y(n1546) );
  OAI21X1 U1297 ( .A(n89), .B(n1305), .C(n1546), .Y(n2137) );
  NAND2X1 U1298 ( .A(\mem<18><14> ), .B(n1242), .Y(n1547) );
  OAI21X1 U1299 ( .A(n89), .B(n1306), .C(n1547), .Y(n2136) );
  NAND2X1 U1300 ( .A(\mem<18><15> ), .B(n1242), .Y(n1548) );
  OAI21X1 U1301 ( .A(n89), .B(n1307), .C(n1548), .Y(n2135) );
  NAND2X1 U1302 ( .A(\mem<17><0> ), .B(n1243), .Y(n1549) );
  OAI21X1 U1303 ( .A(n93), .B(n1292), .C(n1549), .Y(n2134) );
  NAND2X1 U1304 ( .A(\mem<17><1> ), .B(n1243), .Y(n1550) );
  OAI21X1 U1305 ( .A(n93), .B(n1293), .C(n1550), .Y(n2133) );
  NAND2X1 U1306 ( .A(\mem<17><2> ), .B(n1243), .Y(n1551) );
  OAI21X1 U1307 ( .A(n93), .B(n1294), .C(n1551), .Y(n2132) );
  NAND2X1 U1308 ( .A(\mem<17><3> ), .B(n1243), .Y(n1552) );
  OAI21X1 U1309 ( .A(n93), .B(n1295), .C(n1552), .Y(n2131) );
  NAND2X1 U1310 ( .A(\mem<17><4> ), .B(n1243), .Y(n1553) );
  OAI21X1 U1311 ( .A(n93), .B(n1296), .C(n1553), .Y(n2130) );
  NAND2X1 U1312 ( .A(\mem<17><5> ), .B(n1243), .Y(n1554) );
  OAI21X1 U1313 ( .A(n93), .B(n1297), .C(n1554), .Y(n2129) );
  NAND2X1 U1314 ( .A(\mem<17><6> ), .B(n1243), .Y(n1555) );
  OAI21X1 U1315 ( .A(n93), .B(n1298), .C(n1555), .Y(n2128) );
  NAND2X1 U1316 ( .A(\mem<17><7> ), .B(n1243), .Y(n1556) );
  OAI21X1 U1317 ( .A(n93), .B(n1299), .C(n1556), .Y(n2127) );
  NAND2X1 U1318 ( .A(\mem<17><8> ), .B(n1244), .Y(n1557) );
  OAI21X1 U1319 ( .A(n93), .B(n1300), .C(n1557), .Y(n2126) );
  NAND2X1 U1320 ( .A(\mem<17><9> ), .B(n1244), .Y(n1558) );
  OAI21X1 U1321 ( .A(n93), .B(n1301), .C(n1558), .Y(n2125) );
  NAND2X1 U1322 ( .A(\mem<17><10> ), .B(n1244), .Y(n1559) );
  OAI21X1 U1323 ( .A(n93), .B(n1302), .C(n1559), .Y(n2124) );
  NAND2X1 U1324 ( .A(\mem<17><11> ), .B(n1244), .Y(n1560) );
  OAI21X1 U1325 ( .A(n93), .B(n1303), .C(n1560), .Y(n2123) );
  NAND2X1 U1326 ( .A(\mem<17><12> ), .B(n1244), .Y(n1561) );
  OAI21X1 U1327 ( .A(n93), .B(n1304), .C(n1561), .Y(n2122) );
  NAND2X1 U1328 ( .A(\mem<17><13> ), .B(n1244), .Y(n1562) );
  OAI21X1 U1329 ( .A(n93), .B(n1305), .C(n1562), .Y(n2121) );
  NAND2X1 U1330 ( .A(\mem<17><14> ), .B(n1244), .Y(n1563) );
  OAI21X1 U1331 ( .A(n93), .B(n1306), .C(n1563), .Y(n2120) );
  NAND2X1 U1332 ( .A(\mem<17><15> ), .B(n1244), .Y(n1564) );
  OAI21X1 U1333 ( .A(n93), .B(n1307), .C(n1564), .Y(n2119) );
  NAND2X1 U1334 ( .A(\mem<16><0> ), .B(n1246), .Y(n1565) );
  OAI21X1 U1335 ( .A(n1245), .B(n1292), .C(n1565), .Y(n2118) );
  NAND2X1 U1336 ( .A(\mem<16><1> ), .B(n1246), .Y(n1566) );
  OAI21X1 U1337 ( .A(n1245), .B(n1293), .C(n1566), .Y(n2117) );
  NAND2X1 U1338 ( .A(\mem<16><2> ), .B(n1246), .Y(n1567) );
  OAI21X1 U1339 ( .A(n1245), .B(n1294), .C(n1567), .Y(n2116) );
  NAND2X1 U1340 ( .A(\mem<16><3> ), .B(n1246), .Y(n1568) );
  OAI21X1 U1341 ( .A(n1245), .B(n1295), .C(n1568), .Y(n2115) );
  NAND2X1 U1342 ( .A(\mem<16><4> ), .B(n1246), .Y(n1569) );
  OAI21X1 U1343 ( .A(n1245), .B(n1296), .C(n1569), .Y(n2114) );
  NAND2X1 U1344 ( .A(\mem<16><5> ), .B(n1246), .Y(n1570) );
  OAI21X1 U1345 ( .A(n1245), .B(n1297), .C(n1570), .Y(n2113) );
  NAND2X1 U1346 ( .A(\mem<16><6> ), .B(n1246), .Y(n1571) );
  OAI21X1 U1347 ( .A(n1245), .B(n1298), .C(n1571), .Y(n2112) );
  NAND2X1 U1348 ( .A(\mem<16><7> ), .B(n1246), .Y(n1572) );
  OAI21X1 U1349 ( .A(n1245), .B(n1299), .C(n1572), .Y(n2111) );
  NAND2X1 U1350 ( .A(\mem<16><8> ), .B(n1247), .Y(n1573) );
  OAI21X1 U1351 ( .A(n1245), .B(n1300), .C(n1573), .Y(n2110) );
  NAND2X1 U1352 ( .A(\mem<16><9> ), .B(n1247), .Y(n1574) );
  OAI21X1 U1353 ( .A(n1245), .B(n1301), .C(n1574), .Y(n2109) );
  NAND2X1 U1354 ( .A(\mem<16><10> ), .B(n1247), .Y(n1575) );
  OAI21X1 U1355 ( .A(n1245), .B(n1302), .C(n1575), .Y(n2108) );
  NAND2X1 U1356 ( .A(\mem<16><11> ), .B(n1247), .Y(n1576) );
  OAI21X1 U1357 ( .A(n1245), .B(n1303), .C(n1576), .Y(n2107) );
  NAND2X1 U1358 ( .A(\mem<16><12> ), .B(n1247), .Y(n1577) );
  OAI21X1 U1359 ( .A(n1245), .B(n1304), .C(n1577), .Y(n2106) );
  NAND2X1 U1360 ( .A(\mem<16><13> ), .B(n1247), .Y(n1578) );
  OAI21X1 U1361 ( .A(n1245), .B(n1305), .C(n1578), .Y(n2105) );
  NAND2X1 U1362 ( .A(\mem<16><14> ), .B(n1247), .Y(n1579) );
  OAI21X1 U1363 ( .A(n1245), .B(n1306), .C(n1579), .Y(n2104) );
  NAND2X1 U1364 ( .A(\mem<16><15> ), .B(n1247), .Y(n1580) );
  OAI21X1 U1365 ( .A(n1245), .B(n1307), .C(n1580), .Y(n2103) );
  NAND3X1 U1366 ( .A(n1313), .B(n2359), .C(n1316), .Y(n1581) );
  NAND2X1 U1367 ( .A(\mem<15><0> ), .B(n1250), .Y(n1582) );
  OAI21X1 U1368 ( .A(n1248), .B(n1292), .C(n1582), .Y(n2102) );
  NAND2X1 U1369 ( .A(\mem<15><1> ), .B(n1250), .Y(n1583) );
  OAI21X1 U1370 ( .A(n1248), .B(n1293), .C(n1583), .Y(n2101) );
  NAND2X1 U1371 ( .A(\mem<15><2> ), .B(n1250), .Y(n1584) );
  OAI21X1 U1372 ( .A(n1248), .B(n1294), .C(n1584), .Y(n2100) );
  NAND2X1 U1373 ( .A(\mem<15><3> ), .B(n1250), .Y(n1585) );
  OAI21X1 U1374 ( .A(n1248), .B(n1295), .C(n1585), .Y(n2099) );
  NAND2X1 U1375 ( .A(\mem<15><4> ), .B(n1250), .Y(n1586) );
  OAI21X1 U1376 ( .A(n1248), .B(n1296), .C(n1586), .Y(n2098) );
  NAND2X1 U1377 ( .A(\mem<15><5> ), .B(n1250), .Y(n1587) );
  OAI21X1 U1378 ( .A(n1248), .B(n1297), .C(n1587), .Y(n2097) );
  NAND2X1 U1379 ( .A(\mem<15><6> ), .B(n1250), .Y(n1588) );
  OAI21X1 U1380 ( .A(n1248), .B(n1298), .C(n1588), .Y(n2096) );
  NAND2X1 U1381 ( .A(\mem<15><7> ), .B(n1250), .Y(n1589) );
  OAI21X1 U1382 ( .A(n1248), .B(n1299), .C(n1589), .Y(n2095) );
  NAND2X1 U1383 ( .A(\mem<15><8> ), .B(n1251), .Y(n1590) );
  OAI21X1 U1384 ( .A(n1249), .B(n1300), .C(n1590), .Y(n2094) );
  NAND2X1 U1385 ( .A(\mem<15><9> ), .B(n1251), .Y(n1591) );
  OAI21X1 U1386 ( .A(n1249), .B(n1301), .C(n1591), .Y(n2093) );
  NAND2X1 U1387 ( .A(\mem<15><10> ), .B(n1251), .Y(n1592) );
  OAI21X1 U1388 ( .A(n1249), .B(n1302), .C(n1592), .Y(n2092) );
  NAND2X1 U1389 ( .A(\mem<15><11> ), .B(n1251), .Y(n1593) );
  OAI21X1 U1390 ( .A(n1249), .B(n1303), .C(n1593), .Y(n2091) );
  NAND2X1 U1391 ( .A(\mem<15><12> ), .B(n1251), .Y(n1594) );
  OAI21X1 U1392 ( .A(n1249), .B(n1304), .C(n1594), .Y(n2090) );
  NAND2X1 U1393 ( .A(\mem<15><13> ), .B(n1251), .Y(n1595) );
  OAI21X1 U1394 ( .A(n1249), .B(n1305), .C(n1595), .Y(n2089) );
  NAND2X1 U1395 ( .A(\mem<15><14> ), .B(n1251), .Y(n1596) );
  OAI21X1 U1396 ( .A(n1249), .B(n1306), .C(n1596), .Y(n2088) );
  NAND2X1 U1397 ( .A(\mem<15><15> ), .B(n1251), .Y(n1597) );
  OAI21X1 U1398 ( .A(n1249), .B(n1307), .C(n1597), .Y(n2087) );
  NAND2X1 U1399 ( .A(\mem<14><0> ), .B(n1252), .Y(n1598) );
  OAI21X1 U1400 ( .A(n103), .B(n1292), .C(n1598), .Y(n2086) );
  NAND2X1 U1401 ( .A(\mem<14><1> ), .B(n1252), .Y(n1599) );
  OAI21X1 U1402 ( .A(n103), .B(n1293), .C(n1599), .Y(n2085) );
  NAND2X1 U1403 ( .A(\mem<14><2> ), .B(n1252), .Y(n1600) );
  OAI21X1 U1404 ( .A(n103), .B(n1294), .C(n1600), .Y(n2084) );
  NAND2X1 U1405 ( .A(\mem<14><3> ), .B(n1252), .Y(n1601) );
  OAI21X1 U1406 ( .A(n103), .B(n1295), .C(n1601), .Y(n2083) );
  NAND2X1 U1407 ( .A(\mem<14><4> ), .B(n1252), .Y(n1602) );
  OAI21X1 U1408 ( .A(n103), .B(n1296), .C(n1602), .Y(n2082) );
  NAND2X1 U1409 ( .A(\mem<14><5> ), .B(n1252), .Y(n1603) );
  OAI21X1 U1410 ( .A(n103), .B(n1297), .C(n1603), .Y(n2081) );
  NAND2X1 U1411 ( .A(\mem<14><6> ), .B(n1252), .Y(n1604) );
  OAI21X1 U1412 ( .A(n103), .B(n1298), .C(n1604), .Y(n2080) );
  NAND2X1 U1413 ( .A(\mem<14><7> ), .B(n1252), .Y(n1605) );
  OAI21X1 U1414 ( .A(n103), .B(n1299), .C(n1605), .Y(n2079) );
  NAND2X1 U1415 ( .A(\mem<14><8> ), .B(n1253), .Y(n1606) );
  OAI21X1 U1416 ( .A(n103), .B(n1300), .C(n1606), .Y(n2078) );
  NAND2X1 U1417 ( .A(\mem<14><9> ), .B(n1253), .Y(n1607) );
  OAI21X1 U1418 ( .A(n103), .B(n1301), .C(n1607), .Y(n2077) );
  NAND2X1 U1419 ( .A(\mem<14><10> ), .B(n1253), .Y(n1608) );
  OAI21X1 U1420 ( .A(n103), .B(n1302), .C(n1608), .Y(n2076) );
  NAND2X1 U1421 ( .A(\mem<14><11> ), .B(n1253), .Y(n1609) );
  OAI21X1 U1422 ( .A(n103), .B(n1303), .C(n1609), .Y(n2075) );
  NAND2X1 U1423 ( .A(\mem<14><12> ), .B(n1253), .Y(n1610) );
  OAI21X1 U1424 ( .A(n103), .B(n1304), .C(n1610), .Y(n2074) );
  NAND2X1 U1425 ( .A(\mem<14><13> ), .B(n1253), .Y(n1611) );
  OAI21X1 U1426 ( .A(n103), .B(n1305), .C(n1611), .Y(n2073) );
  NAND2X1 U1427 ( .A(\mem<14><14> ), .B(n1253), .Y(n1612) );
  OAI21X1 U1428 ( .A(n103), .B(n1306), .C(n1612), .Y(n2072) );
  NAND2X1 U1429 ( .A(\mem<14><15> ), .B(n1253), .Y(n1613) );
  OAI21X1 U1430 ( .A(n103), .B(n1307), .C(n1613), .Y(n2071) );
  NAND2X1 U1431 ( .A(\mem<13><0> ), .B(n1255), .Y(n1614) );
  OAI21X1 U1432 ( .A(n1254), .B(n1292), .C(n1614), .Y(n2070) );
  NAND2X1 U1433 ( .A(\mem<13><1> ), .B(n1255), .Y(n1615) );
  OAI21X1 U1434 ( .A(n1254), .B(n1293), .C(n1615), .Y(n2069) );
  NAND2X1 U1435 ( .A(\mem<13><2> ), .B(n1255), .Y(n1616) );
  OAI21X1 U1436 ( .A(n1254), .B(n1294), .C(n1616), .Y(n2068) );
  NAND2X1 U1437 ( .A(\mem<13><3> ), .B(n1255), .Y(n1617) );
  OAI21X1 U1438 ( .A(n1254), .B(n1295), .C(n1617), .Y(n2067) );
  NAND2X1 U1439 ( .A(\mem<13><4> ), .B(n1255), .Y(n1618) );
  OAI21X1 U1440 ( .A(n1254), .B(n1296), .C(n1618), .Y(n2066) );
  NAND2X1 U1441 ( .A(\mem<13><5> ), .B(n1255), .Y(n1619) );
  OAI21X1 U1442 ( .A(n1254), .B(n1297), .C(n1619), .Y(n2065) );
  NAND2X1 U1443 ( .A(\mem<13><6> ), .B(n1255), .Y(n1620) );
  OAI21X1 U1444 ( .A(n1254), .B(n1298), .C(n1620), .Y(n2064) );
  NAND2X1 U1445 ( .A(\mem<13><7> ), .B(n1255), .Y(n1621) );
  OAI21X1 U1446 ( .A(n1254), .B(n1299), .C(n1621), .Y(n2063) );
  NAND2X1 U1447 ( .A(\mem<13><8> ), .B(n1256), .Y(n1622) );
  OAI21X1 U1448 ( .A(n107), .B(n1300), .C(n1622), .Y(n2062) );
  NAND2X1 U1449 ( .A(\mem<13><9> ), .B(n1256), .Y(n1623) );
  OAI21X1 U1450 ( .A(n107), .B(n1301), .C(n1623), .Y(n2061) );
  NAND2X1 U1451 ( .A(\mem<13><10> ), .B(n1256), .Y(n1624) );
  OAI21X1 U1452 ( .A(n107), .B(n1302), .C(n1624), .Y(n2060) );
  NAND2X1 U1453 ( .A(\mem<13><11> ), .B(n1256), .Y(n1625) );
  OAI21X1 U1454 ( .A(n107), .B(n1303), .C(n1625), .Y(n2059) );
  NAND2X1 U1455 ( .A(\mem<13><12> ), .B(n1256), .Y(n1626) );
  OAI21X1 U1456 ( .A(n107), .B(n1304), .C(n1626), .Y(n2058) );
  NAND2X1 U1457 ( .A(\mem<13><13> ), .B(n1256), .Y(n1627) );
  OAI21X1 U1458 ( .A(n107), .B(n1305), .C(n1627), .Y(n2057) );
  NAND2X1 U1459 ( .A(\mem<13><14> ), .B(n1256), .Y(n1628) );
  OAI21X1 U1460 ( .A(n1254), .B(n1306), .C(n1628), .Y(n2056) );
  NAND2X1 U1461 ( .A(\mem<13><15> ), .B(n1256), .Y(n1629) );
  OAI21X1 U1462 ( .A(n1254), .B(n1307), .C(n1629), .Y(n2055) );
  NAND2X1 U1463 ( .A(\mem<12><0> ), .B(n1258), .Y(n1630) );
  OAI21X1 U1464 ( .A(n1257), .B(n1292), .C(n1630), .Y(n2054) );
  NAND2X1 U1465 ( .A(\mem<12><1> ), .B(n1258), .Y(n1631) );
  OAI21X1 U1466 ( .A(n1257), .B(n1293), .C(n1631), .Y(n2053) );
  NAND2X1 U1467 ( .A(\mem<12><2> ), .B(n1258), .Y(n1632) );
  OAI21X1 U1468 ( .A(n1257), .B(n1294), .C(n1632), .Y(n2052) );
  NAND2X1 U1469 ( .A(\mem<12><3> ), .B(n1258), .Y(n1633) );
  OAI21X1 U1470 ( .A(n1257), .B(n1295), .C(n1633), .Y(n2051) );
  NAND2X1 U1471 ( .A(\mem<12><4> ), .B(n1258), .Y(n1634) );
  OAI21X1 U1472 ( .A(n1257), .B(n1296), .C(n1634), .Y(n2050) );
  NAND2X1 U1473 ( .A(\mem<12><5> ), .B(n1258), .Y(n1635) );
  OAI21X1 U1474 ( .A(n1257), .B(n1297), .C(n1635), .Y(n2049) );
  NAND2X1 U1475 ( .A(\mem<12><6> ), .B(n1258), .Y(n1636) );
  OAI21X1 U1476 ( .A(n1257), .B(n1298), .C(n1636), .Y(n2048) );
  NAND2X1 U1477 ( .A(\mem<12><7> ), .B(n1258), .Y(n1637) );
  OAI21X1 U1478 ( .A(n1257), .B(n1299), .C(n1637), .Y(n2047) );
  NAND2X1 U1479 ( .A(\mem<12><8> ), .B(n1259), .Y(n1638) );
  OAI21X1 U1480 ( .A(n111), .B(n1300), .C(n1638), .Y(n2046) );
  NAND2X1 U1481 ( .A(\mem<12><9> ), .B(n1259), .Y(n1639) );
  OAI21X1 U1482 ( .A(n111), .B(n1301), .C(n1639), .Y(n2045) );
  NAND2X1 U1483 ( .A(\mem<12><10> ), .B(n1259), .Y(n1640) );
  OAI21X1 U1484 ( .A(n111), .B(n1302), .C(n1640), .Y(n2044) );
  NAND2X1 U1485 ( .A(\mem<12><11> ), .B(n1259), .Y(n1641) );
  OAI21X1 U1486 ( .A(n111), .B(n1303), .C(n1641), .Y(n2043) );
  NAND2X1 U1487 ( .A(\mem<12><12> ), .B(n1259), .Y(n1642) );
  OAI21X1 U1488 ( .A(n111), .B(n1304), .C(n1642), .Y(n2042) );
  NAND2X1 U1489 ( .A(\mem<12><13> ), .B(n1259), .Y(n1643) );
  OAI21X1 U1490 ( .A(n111), .B(n1305), .C(n1643), .Y(n2041) );
  NAND2X1 U1491 ( .A(\mem<12><14> ), .B(n1259), .Y(n1644) );
  OAI21X1 U1492 ( .A(n1257), .B(n1306), .C(n1644), .Y(n2040) );
  NAND2X1 U1493 ( .A(\mem<12><15> ), .B(n1259), .Y(n1645) );
  OAI21X1 U1494 ( .A(n1257), .B(n1307), .C(n1645), .Y(n2039) );
  NAND2X1 U1495 ( .A(\mem<11><0> ), .B(n1260), .Y(n1646) );
  OAI21X1 U1496 ( .A(n115), .B(n1292), .C(n1646), .Y(n2038) );
  NAND2X1 U1497 ( .A(\mem<11><1> ), .B(n1260), .Y(n1647) );
  OAI21X1 U1498 ( .A(n115), .B(n1293), .C(n1647), .Y(n2037) );
  NAND2X1 U1499 ( .A(\mem<11><2> ), .B(n1260), .Y(n1648) );
  OAI21X1 U1500 ( .A(n115), .B(n1294), .C(n1648), .Y(n2036) );
  NAND2X1 U1501 ( .A(\mem<11><3> ), .B(n1260), .Y(n1649) );
  OAI21X1 U1502 ( .A(n115), .B(n1295), .C(n1649), .Y(n2035) );
  NAND2X1 U1503 ( .A(\mem<11><4> ), .B(n1260), .Y(n1650) );
  OAI21X1 U1504 ( .A(n115), .B(n1296), .C(n1650), .Y(n2034) );
  NAND2X1 U1505 ( .A(\mem<11><5> ), .B(n1260), .Y(n1651) );
  OAI21X1 U1506 ( .A(n115), .B(n1297), .C(n1651), .Y(n2033) );
  NAND2X1 U1507 ( .A(\mem<11><6> ), .B(n1260), .Y(n1652) );
  OAI21X1 U1508 ( .A(n115), .B(n1298), .C(n1652), .Y(n2032) );
  NAND2X1 U1509 ( .A(\mem<11><7> ), .B(n1260), .Y(n1653) );
  OAI21X1 U1510 ( .A(n115), .B(n1299), .C(n1653), .Y(n2031) );
  NAND2X1 U1511 ( .A(\mem<11><8> ), .B(n1261), .Y(n1654) );
  OAI21X1 U1512 ( .A(n115), .B(n1300), .C(n1654), .Y(n2030) );
  NAND2X1 U1513 ( .A(\mem<11><9> ), .B(n1261), .Y(n1655) );
  OAI21X1 U1514 ( .A(n115), .B(n1301), .C(n1655), .Y(n2029) );
  NAND2X1 U1515 ( .A(\mem<11><10> ), .B(n1261), .Y(n1656) );
  OAI21X1 U1516 ( .A(n115), .B(n1302), .C(n1656), .Y(n2028) );
  NAND2X1 U1517 ( .A(\mem<11><11> ), .B(n1261), .Y(n1657) );
  OAI21X1 U1518 ( .A(n115), .B(n1303), .C(n1657), .Y(n2027) );
  NAND2X1 U1519 ( .A(\mem<11><12> ), .B(n1261), .Y(n1658) );
  OAI21X1 U1520 ( .A(n115), .B(n1304), .C(n1658), .Y(n2026) );
  NAND2X1 U1521 ( .A(\mem<11><13> ), .B(n1261), .Y(n1659) );
  OAI21X1 U1522 ( .A(n115), .B(n1305), .C(n1659), .Y(n2025) );
  NAND2X1 U1523 ( .A(\mem<11><14> ), .B(n1261), .Y(n1660) );
  OAI21X1 U1524 ( .A(n115), .B(n1306), .C(n1660), .Y(n2024) );
  NAND2X1 U1525 ( .A(\mem<11><15> ), .B(n1261), .Y(n1661) );
  OAI21X1 U1526 ( .A(n115), .B(n1307), .C(n1661), .Y(n2023) );
  NAND2X1 U1527 ( .A(\mem<10><0> ), .B(n1262), .Y(n1662) );
  OAI21X1 U1528 ( .A(n119), .B(n1292), .C(n1662), .Y(n2022) );
  NAND2X1 U1529 ( .A(\mem<10><1> ), .B(n1262), .Y(n1663) );
  OAI21X1 U1530 ( .A(n119), .B(n1293), .C(n1663), .Y(n2021) );
  NAND2X1 U1531 ( .A(\mem<10><2> ), .B(n1262), .Y(n1664) );
  OAI21X1 U1532 ( .A(n119), .B(n1294), .C(n1664), .Y(n2020) );
  NAND2X1 U1533 ( .A(\mem<10><3> ), .B(n1262), .Y(n1665) );
  OAI21X1 U1534 ( .A(n119), .B(n1295), .C(n1665), .Y(n2019) );
  NAND2X1 U1535 ( .A(\mem<10><4> ), .B(n1262), .Y(n1666) );
  OAI21X1 U1536 ( .A(n119), .B(n1296), .C(n1666), .Y(n2018) );
  NAND2X1 U1537 ( .A(\mem<10><5> ), .B(n1262), .Y(n1667) );
  OAI21X1 U1538 ( .A(n119), .B(n1297), .C(n1667), .Y(n2017) );
  NAND2X1 U1539 ( .A(\mem<10><6> ), .B(n1262), .Y(n1668) );
  OAI21X1 U1540 ( .A(n119), .B(n1298), .C(n1668), .Y(n2016) );
  NAND2X1 U1541 ( .A(\mem<10><7> ), .B(n1262), .Y(n1669) );
  OAI21X1 U1542 ( .A(n119), .B(n1299), .C(n1669), .Y(n2015) );
  NAND2X1 U1543 ( .A(\mem<10><8> ), .B(n1263), .Y(n1670) );
  OAI21X1 U1544 ( .A(n119), .B(n1300), .C(n1670), .Y(n2014) );
  NAND2X1 U1545 ( .A(\mem<10><9> ), .B(n1263), .Y(n1671) );
  OAI21X1 U1546 ( .A(n119), .B(n1301), .C(n1671), .Y(n2013) );
  NAND2X1 U1547 ( .A(\mem<10><10> ), .B(n1263), .Y(n1672) );
  OAI21X1 U1548 ( .A(n119), .B(n1302), .C(n1672), .Y(n2012) );
  NAND2X1 U1549 ( .A(\mem<10><11> ), .B(n1263), .Y(n1673) );
  OAI21X1 U1550 ( .A(n119), .B(n1303), .C(n1673), .Y(n2011) );
  NAND2X1 U1551 ( .A(\mem<10><12> ), .B(n1263), .Y(n1674) );
  OAI21X1 U1552 ( .A(n119), .B(n1304), .C(n1674), .Y(n2010) );
  NAND2X1 U1553 ( .A(\mem<10><13> ), .B(n1263), .Y(n1675) );
  OAI21X1 U1554 ( .A(n119), .B(n1305), .C(n1675), .Y(n2009) );
  NAND2X1 U1555 ( .A(\mem<10><14> ), .B(n1263), .Y(n1676) );
  OAI21X1 U1556 ( .A(n119), .B(n1306), .C(n1676), .Y(n2008) );
  NAND2X1 U1557 ( .A(\mem<10><15> ), .B(n1263), .Y(n1677) );
  OAI21X1 U1558 ( .A(n119), .B(n1307), .C(n1677), .Y(n2007) );
  NAND2X1 U1559 ( .A(\mem<9><0> ), .B(n1264), .Y(n1678) );
  OAI21X1 U1560 ( .A(n123), .B(n1292), .C(n1678), .Y(n2006) );
  NAND2X1 U1561 ( .A(\mem<9><1> ), .B(n1264), .Y(n1679) );
  OAI21X1 U1562 ( .A(n123), .B(n1293), .C(n1679), .Y(n2005) );
  NAND2X1 U1563 ( .A(\mem<9><2> ), .B(n1264), .Y(n1680) );
  OAI21X1 U1564 ( .A(n123), .B(n1294), .C(n1680), .Y(n2004) );
  NAND2X1 U1565 ( .A(\mem<9><3> ), .B(n1264), .Y(n1681) );
  OAI21X1 U1566 ( .A(n123), .B(n1295), .C(n1681), .Y(n2003) );
  NAND2X1 U1567 ( .A(\mem<9><4> ), .B(n1264), .Y(n1682) );
  OAI21X1 U1568 ( .A(n123), .B(n1296), .C(n1682), .Y(n2002) );
  NAND2X1 U1569 ( .A(\mem<9><5> ), .B(n1264), .Y(n1683) );
  OAI21X1 U1570 ( .A(n123), .B(n1297), .C(n1683), .Y(n2001) );
  NAND2X1 U1571 ( .A(\mem<9><6> ), .B(n1264), .Y(n1684) );
  OAI21X1 U1572 ( .A(n123), .B(n1298), .C(n1684), .Y(n2000) );
  NAND2X1 U1573 ( .A(\mem<9><7> ), .B(n1264), .Y(n1685) );
  OAI21X1 U1574 ( .A(n123), .B(n1299), .C(n1685), .Y(n1999) );
  NAND2X1 U1575 ( .A(\mem<9><8> ), .B(n1265), .Y(n1686) );
  OAI21X1 U1576 ( .A(n123), .B(n1300), .C(n1686), .Y(n1998) );
  NAND2X1 U1577 ( .A(\mem<9><9> ), .B(n1265), .Y(n1687) );
  OAI21X1 U1578 ( .A(n123), .B(n1301), .C(n1687), .Y(n1997) );
  NAND2X1 U1579 ( .A(\mem<9><10> ), .B(n1265), .Y(n1688) );
  OAI21X1 U1580 ( .A(n123), .B(n1302), .C(n1688), .Y(n1996) );
  NAND2X1 U1581 ( .A(\mem<9><11> ), .B(n1265), .Y(n1689) );
  OAI21X1 U1582 ( .A(n123), .B(n1303), .C(n1689), .Y(n1995) );
  NAND2X1 U1583 ( .A(\mem<9><12> ), .B(n1265), .Y(n1690) );
  OAI21X1 U1584 ( .A(n123), .B(n1304), .C(n1690), .Y(n1994) );
  NAND2X1 U1585 ( .A(\mem<9><13> ), .B(n1265), .Y(n1691) );
  OAI21X1 U1586 ( .A(n123), .B(n1305), .C(n1691), .Y(n1993) );
  NAND2X1 U1587 ( .A(\mem<9><14> ), .B(n1265), .Y(n1692) );
  OAI21X1 U1588 ( .A(n123), .B(n1306), .C(n1692), .Y(n1992) );
  NAND2X1 U1589 ( .A(\mem<9><15> ), .B(n1265), .Y(n1693) );
  OAI21X1 U1590 ( .A(n123), .B(n1307), .C(n1693), .Y(n1991) );
  NAND2X1 U1591 ( .A(\mem<8><0> ), .B(n1266), .Y(n1695) );
  OAI21X1 U1592 ( .A(n35), .B(n1292), .C(n1695), .Y(n1990) );
  NAND2X1 U1593 ( .A(\mem<8><1> ), .B(n1266), .Y(n1696) );
  OAI21X1 U1594 ( .A(n35), .B(n1293), .C(n1696), .Y(n1989) );
  NAND2X1 U1595 ( .A(\mem<8><2> ), .B(n1266), .Y(n1697) );
  OAI21X1 U1596 ( .A(n35), .B(n1294), .C(n1697), .Y(n1988) );
  NAND2X1 U1597 ( .A(\mem<8><3> ), .B(n1266), .Y(n1698) );
  OAI21X1 U1598 ( .A(n35), .B(n1295), .C(n1698), .Y(n1987) );
  NAND2X1 U1599 ( .A(\mem<8><4> ), .B(n1266), .Y(n1699) );
  OAI21X1 U1600 ( .A(n35), .B(n1296), .C(n1699), .Y(n1986) );
  NAND2X1 U1601 ( .A(\mem<8><5> ), .B(n1266), .Y(n1700) );
  OAI21X1 U1602 ( .A(n35), .B(n1297), .C(n1700), .Y(n1985) );
  NAND2X1 U1603 ( .A(\mem<8><6> ), .B(n1266), .Y(n1701) );
  OAI21X1 U1604 ( .A(n35), .B(n1298), .C(n1701), .Y(n1984) );
  NAND2X1 U1605 ( .A(\mem<8><7> ), .B(n1266), .Y(n1702) );
  OAI21X1 U1606 ( .A(n35), .B(n1299), .C(n1702), .Y(n1983) );
  NAND2X1 U1607 ( .A(\mem<8><8> ), .B(n1267), .Y(n1703) );
  OAI21X1 U1608 ( .A(n35), .B(n1300), .C(n1703), .Y(n1982) );
  NAND2X1 U1609 ( .A(\mem<8><9> ), .B(n1267), .Y(n1704) );
  OAI21X1 U1610 ( .A(n35), .B(n1301), .C(n1704), .Y(n1981) );
  NAND2X1 U1611 ( .A(\mem<8><10> ), .B(n1267), .Y(n1705) );
  OAI21X1 U1612 ( .A(n35), .B(n1302), .C(n1705), .Y(n1980) );
  NAND2X1 U1613 ( .A(\mem<8><11> ), .B(n1267), .Y(n1706) );
  OAI21X1 U1614 ( .A(n35), .B(n1303), .C(n1706), .Y(n1979) );
  NAND2X1 U1615 ( .A(\mem<8><12> ), .B(n1267), .Y(n1707) );
  OAI21X1 U1616 ( .A(n35), .B(n1304), .C(n1707), .Y(n1978) );
  NAND2X1 U1617 ( .A(\mem<8><13> ), .B(n1267), .Y(n1708) );
  OAI21X1 U1618 ( .A(n35), .B(n1305), .C(n1708), .Y(n1977) );
  NAND2X1 U1619 ( .A(\mem<8><14> ), .B(n1267), .Y(n1709) );
  OAI21X1 U1620 ( .A(n35), .B(n1306), .C(n1709), .Y(n1976) );
  NAND2X1 U1621 ( .A(\mem<8><15> ), .B(n1267), .Y(n1710) );
  OAI21X1 U1622 ( .A(n35), .B(n1307), .C(n1710), .Y(n1975) );
  NAND3X1 U1623 ( .A(n1314), .B(n2359), .C(n1316), .Y(n1711) );
  NAND2X1 U1624 ( .A(\mem<7><0> ), .B(n1270), .Y(n1712) );
  OAI21X1 U1625 ( .A(n1268), .B(n1292), .C(n1712), .Y(n1974) );
  NAND2X1 U1626 ( .A(\mem<7><1> ), .B(n1270), .Y(n1713) );
  OAI21X1 U1627 ( .A(n1268), .B(n1293), .C(n1713), .Y(n1973) );
  NAND2X1 U1628 ( .A(\mem<7><2> ), .B(n1270), .Y(n1714) );
  OAI21X1 U1629 ( .A(n1268), .B(n1294), .C(n1714), .Y(n1972) );
  NAND2X1 U1630 ( .A(\mem<7><3> ), .B(n1270), .Y(n1715) );
  OAI21X1 U1631 ( .A(n1268), .B(n1295), .C(n1715), .Y(n1971) );
  NAND2X1 U1632 ( .A(\mem<7><4> ), .B(n1270), .Y(n1716) );
  OAI21X1 U1633 ( .A(n1268), .B(n1296), .C(n1716), .Y(n1970) );
  NAND2X1 U1634 ( .A(\mem<7><5> ), .B(n1270), .Y(n1717) );
  OAI21X1 U1635 ( .A(n1268), .B(n1297), .C(n1717), .Y(n1969) );
  NAND2X1 U1636 ( .A(\mem<7><6> ), .B(n1270), .Y(n1718) );
  OAI21X1 U1637 ( .A(n1268), .B(n1298), .C(n1718), .Y(n1968) );
  NAND2X1 U1638 ( .A(\mem<7><7> ), .B(n1270), .Y(n1719) );
  OAI21X1 U1639 ( .A(n1268), .B(n1299), .C(n1719), .Y(n1967) );
  NAND2X1 U1640 ( .A(\mem<7><8> ), .B(n1271), .Y(n1720) );
  OAI21X1 U1641 ( .A(n1269), .B(n1300), .C(n1720), .Y(n1966) );
  NAND2X1 U1642 ( .A(\mem<7><9> ), .B(n1271), .Y(n1721) );
  OAI21X1 U1643 ( .A(n1269), .B(n1301), .C(n1721), .Y(n1965) );
  NAND2X1 U1644 ( .A(\mem<7><10> ), .B(n1271), .Y(n1722) );
  OAI21X1 U1645 ( .A(n1269), .B(n1302), .C(n1722), .Y(n1964) );
  NAND2X1 U1646 ( .A(\mem<7><11> ), .B(n1271), .Y(n1723) );
  OAI21X1 U1647 ( .A(n1269), .B(n1303), .C(n1723), .Y(n1963) );
  NAND2X1 U1648 ( .A(\mem<7><12> ), .B(n1271), .Y(n1724) );
  OAI21X1 U1649 ( .A(n1269), .B(n1304), .C(n1724), .Y(n1962) );
  NAND2X1 U1650 ( .A(\mem<7><13> ), .B(n1271), .Y(n1725) );
  OAI21X1 U1651 ( .A(n1269), .B(n1305), .C(n1725), .Y(n1961) );
  NAND2X1 U1652 ( .A(\mem<7><14> ), .B(n1271), .Y(n1726) );
  OAI21X1 U1653 ( .A(n1269), .B(n1306), .C(n1726), .Y(n1960) );
  NAND2X1 U1654 ( .A(\mem<7><15> ), .B(n1271), .Y(n1727) );
  OAI21X1 U1655 ( .A(n1269), .B(n1307), .C(n1727), .Y(n1959) );
  NAND2X1 U1656 ( .A(\mem<6><0> ), .B(n1272), .Y(n1728) );
  OAI21X1 U1657 ( .A(n133), .B(n1292), .C(n1728), .Y(n1958) );
  NAND2X1 U1658 ( .A(\mem<6><1> ), .B(n1272), .Y(n1729) );
  OAI21X1 U1659 ( .A(n133), .B(n1293), .C(n1729), .Y(n1957) );
  NAND2X1 U1660 ( .A(\mem<6><2> ), .B(n1272), .Y(n1730) );
  OAI21X1 U1661 ( .A(n133), .B(n1294), .C(n1730), .Y(n1956) );
  NAND2X1 U1662 ( .A(\mem<6><3> ), .B(n1272), .Y(n1731) );
  OAI21X1 U1663 ( .A(n133), .B(n1295), .C(n1731), .Y(n1955) );
  NAND2X1 U1664 ( .A(\mem<6><4> ), .B(n1272), .Y(n1732) );
  OAI21X1 U1665 ( .A(n133), .B(n1296), .C(n1732), .Y(n1954) );
  NAND2X1 U1666 ( .A(\mem<6><5> ), .B(n1272), .Y(n1733) );
  OAI21X1 U1667 ( .A(n133), .B(n1297), .C(n1733), .Y(n1953) );
  NAND2X1 U1668 ( .A(\mem<6><6> ), .B(n1272), .Y(n1734) );
  OAI21X1 U1669 ( .A(n133), .B(n1298), .C(n1734), .Y(n1952) );
  NAND2X1 U1670 ( .A(\mem<6><7> ), .B(n1272), .Y(n1735) );
  OAI21X1 U1671 ( .A(n133), .B(n1299), .C(n1735), .Y(n1951) );
  NAND2X1 U1672 ( .A(\mem<6><8> ), .B(n1273), .Y(n1736) );
  OAI21X1 U1673 ( .A(n133), .B(n1300), .C(n1736), .Y(n1950) );
  NAND2X1 U1674 ( .A(\mem<6><9> ), .B(n1273), .Y(n1737) );
  OAI21X1 U1675 ( .A(n133), .B(n1301), .C(n1737), .Y(n1949) );
  NAND2X1 U1676 ( .A(\mem<6><10> ), .B(n1273), .Y(n1738) );
  OAI21X1 U1677 ( .A(n133), .B(n1302), .C(n1738), .Y(n1948) );
  NAND2X1 U1678 ( .A(\mem<6><11> ), .B(n1273), .Y(n1739) );
  OAI21X1 U1679 ( .A(n133), .B(n1303), .C(n1739), .Y(n1947) );
  NAND2X1 U1680 ( .A(\mem<6><12> ), .B(n1273), .Y(n1740) );
  OAI21X1 U1681 ( .A(n133), .B(n1304), .C(n1740), .Y(n1946) );
  NAND2X1 U1682 ( .A(\mem<6><13> ), .B(n1273), .Y(n1741) );
  OAI21X1 U1683 ( .A(n133), .B(n1305), .C(n1741), .Y(n1945) );
  NAND2X1 U1684 ( .A(\mem<6><14> ), .B(n1273), .Y(n1742) );
  OAI21X1 U1685 ( .A(n133), .B(n1306), .C(n1742), .Y(n1944) );
  NAND2X1 U1686 ( .A(\mem<6><15> ), .B(n1273), .Y(n1743) );
  OAI21X1 U1687 ( .A(n133), .B(n1307), .C(n1743), .Y(n1943) );
  NAND2X1 U1688 ( .A(\mem<5><0> ), .B(n1275), .Y(n1745) );
  OAI21X1 U1689 ( .A(n1274), .B(n1292), .C(n1745), .Y(n1942) );
  NAND2X1 U1690 ( .A(\mem<5><1> ), .B(n1275), .Y(n1746) );
  OAI21X1 U1691 ( .A(n1274), .B(n1293), .C(n1746), .Y(n1941) );
  NAND2X1 U1692 ( .A(\mem<5><2> ), .B(n1275), .Y(n1747) );
  OAI21X1 U1693 ( .A(n1274), .B(n1294), .C(n1747), .Y(n1940) );
  NAND2X1 U1694 ( .A(\mem<5><3> ), .B(n1275), .Y(n1748) );
  OAI21X1 U1695 ( .A(n1274), .B(n1295), .C(n1748), .Y(n1939) );
  NAND2X1 U1696 ( .A(\mem<5><4> ), .B(n1275), .Y(n1749) );
  OAI21X1 U1697 ( .A(n1274), .B(n1296), .C(n1749), .Y(n1938) );
  NAND2X1 U1698 ( .A(\mem<5><5> ), .B(n1275), .Y(n1750) );
  OAI21X1 U1699 ( .A(n1274), .B(n1297), .C(n1750), .Y(n1937) );
  NAND2X1 U1700 ( .A(\mem<5><6> ), .B(n1275), .Y(n1751) );
  OAI21X1 U1701 ( .A(n1274), .B(n1298), .C(n1751), .Y(n1936) );
  NAND2X1 U1702 ( .A(\mem<5><7> ), .B(n1275), .Y(n1752) );
  OAI21X1 U1703 ( .A(n1274), .B(n1299), .C(n1752), .Y(n1935) );
  NAND2X1 U1704 ( .A(\mem<5><8> ), .B(n1276), .Y(n1753) );
  OAI21X1 U1705 ( .A(n137), .B(n1300), .C(n1753), .Y(n1934) );
  NAND2X1 U1706 ( .A(\mem<5><9> ), .B(n1276), .Y(n1754) );
  OAI21X1 U1707 ( .A(n137), .B(n1301), .C(n1754), .Y(n1933) );
  NAND2X1 U1708 ( .A(\mem<5><10> ), .B(n1276), .Y(n1755) );
  OAI21X1 U1709 ( .A(n137), .B(n1302), .C(n1755), .Y(n1932) );
  NAND2X1 U1710 ( .A(\mem<5><11> ), .B(n1276), .Y(n1756) );
  OAI21X1 U1711 ( .A(n137), .B(n1303), .C(n1756), .Y(n1931) );
  NAND2X1 U1712 ( .A(\mem<5><12> ), .B(n1276), .Y(n1757) );
  OAI21X1 U1713 ( .A(n137), .B(n1304), .C(n1757), .Y(n1930) );
  NAND2X1 U1714 ( .A(\mem<5><13> ), .B(n1276), .Y(n1758) );
  OAI21X1 U1715 ( .A(n137), .B(n1305), .C(n1758), .Y(n1929) );
  NAND2X1 U1716 ( .A(\mem<5><14> ), .B(n1276), .Y(n1759) );
  OAI21X1 U1717 ( .A(n1274), .B(n1306), .C(n1759), .Y(n1928) );
  NAND2X1 U1718 ( .A(\mem<5><15> ), .B(n1276), .Y(n1760) );
  OAI21X1 U1719 ( .A(n1274), .B(n1307), .C(n1760), .Y(n1927) );
  NAND2X1 U1720 ( .A(\mem<4><0> ), .B(n1278), .Y(n1762) );
  OAI21X1 U1721 ( .A(n1277), .B(n1292), .C(n1762), .Y(n1926) );
  NAND2X1 U1722 ( .A(\mem<4><1> ), .B(n1278), .Y(n1763) );
  OAI21X1 U1723 ( .A(n1277), .B(n1293), .C(n1763), .Y(n1925) );
  NAND2X1 U1724 ( .A(\mem<4><2> ), .B(n1278), .Y(n1764) );
  OAI21X1 U1725 ( .A(n1277), .B(n1294), .C(n1764), .Y(n1924) );
  NAND2X1 U1726 ( .A(\mem<4><3> ), .B(n1278), .Y(n1765) );
  OAI21X1 U1727 ( .A(n1277), .B(n1295), .C(n1765), .Y(n1923) );
  NAND2X1 U1728 ( .A(\mem<4><4> ), .B(n1278), .Y(n1766) );
  OAI21X1 U1729 ( .A(n1277), .B(n1296), .C(n1766), .Y(n1922) );
  NAND2X1 U1730 ( .A(\mem<4><5> ), .B(n1278), .Y(n1767) );
  OAI21X1 U1731 ( .A(n1277), .B(n1297), .C(n1767), .Y(n1921) );
  NAND2X1 U1732 ( .A(\mem<4><6> ), .B(n1278), .Y(n1768) );
  OAI21X1 U1733 ( .A(n1277), .B(n1298), .C(n1768), .Y(n1920) );
  NAND2X1 U1734 ( .A(\mem<4><7> ), .B(n1278), .Y(n1769) );
  OAI21X1 U1735 ( .A(n1277), .B(n1299), .C(n1769), .Y(n1919) );
  NAND2X1 U1736 ( .A(\mem<4><8> ), .B(n1279), .Y(n1770) );
  OAI21X1 U1737 ( .A(n141), .B(n1300), .C(n1770), .Y(n1918) );
  NAND2X1 U1738 ( .A(\mem<4><9> ), .B(n1279), .Y(n1771) );
  OAI21X1 U1739 ( .A(n141), .B(n1301), .C(n1771), .Y(n1917) );
  NAND2X1 U1740 ( .A(\mem<4><10> ), .B(n1279), .Y(n1772) );
  OAI21X1 U1741 ( .A(n141), .B(n1302), .C(n1772), .Y(n1916) );
  NAND2X1 U1742 ( .A(\mem<4><11> ), .B(n1279), .Y(n1773) );
  OAI21X1 U1743 ( .A(n141), .B(n1303), .C(n1773), .Y(n1915) );
  NAND2X1 U1744 ( .A(\mem<4><12> ), .B(n1279), .Y(n1774) );
  OAI21X1 U1745 ( .A(n141), .B(n1304), .C(n1774), .Y(n1914) );
  NAND2X1 U1746 ( .A(\mem<4><13> ), .B(n1279), .Y(n1775) );
  OAI21X1 U1747 ( .A(n141), .B(n1305), .C(n1775), .Y(n1913) );
  NAND2X1 U1748 ( .A(\mem<4><14> ), .B(n1279), .Y(n1776) );
  OAI21X1 U1749 ( .A(n1277), .B(n1306), .C(n1776), .Y(n1912) );
  NAND2X1 U1750 ( .A(\mem<4><15> ), .B(n1279), .Y(n1777) );
  OAI21X1 U1751 ( .A(n1277), .B(n1307), .C(n1777), .Y(n1911) );
  NAND2X1 U1752 ( .A(\mem<3><0> ), .B(n1280), .Y(n1779) );
  OAI21X1 U1753 ( .A(n145), .B(n1292), .C(n1779), .Y(n1910) );
  NAND2X1 U1754 ( .A(\mem<3><1> ), .B(n1280), .Y(n1780) );
  OAI21X1 U1755 ( .A(n145), .B(n1293), .C(n1780), .Y(n1909) );
  NAND2X1 U1756 ( .A(\mem<3><2> ), .B(n1280), .Y(n1781) );
  OAI21X1 U1757 ( .A(n145), .B(n1294), .C(n1781), .Y(n1908) );
  NAND2X1 U1758 ( .A(\mem<3><3> ), .B(n1280), .Y(n1782) );
  OAI21X1 U1759 ( .A(n145), .B(n1295), .C(n1782), .Y(n1907) );
  NAND2X1 U1760 ( .A(\mem<3><4> ), .B(n1280), .Y(n1783) );
  OAI21X1 U1761 ( .A(n145), .B(n1296), .C(n1783), .Y(n1906) );
  NAND2X1 U1762 ( .A(\mem<3><5> ), .B(n1280), .Y(n1784) );
  OAI21X1 U1763 ( .A(n145), .B(n1297), .C(n1784), .Y(n1905) );
  NAND2X1 U1764 ( .A(\mem<3><6> ), .B(n1280), .Y(n1785) );
  OAI21X1 U1765 ( .A(n145), .B(n1298), .C(n1785), .Y(n1904) );
  NAND2X1 U1766 ( .A(\mem<3><7> ), .B(n1280), .Y(n1786) );
  OAI21X1 U1767 ( .A(n145), .B(n1299), .C(n1786), .Y(n1903) );
  NAND2X1 U1768 ( .A(\mem<3><8> ), .B(n1281), .Y(n1787) );
  OAI21X1 U1769 ( .A(n145), .B(n1300), .C(n1787), .Y(n1902) );
  NAND2X1 U1770 ( .A(\mem<3><9> ), .B(n1281), .Y(n1788) );
  OAI21X1 U1771 ( .A(n145), .B(n1301), .C(n1788), .Y(n1901) );
  NAND2X1 U1772 ( .A(\mem<3><10> ), .B(n1281), .Y(n1789) );
  OAI21X1 U1773 ( .A(n145), .B(n1302), .C(n1789), .Y(n1900) );
  NAND2X1 U1774 ( .A(\mem<3><11> ), .B(n1281), .Y(n1790) );
  OAI21X1 U1775 ( .A(n145), .B(n1303), .C(n1790), .Y(n1899) );
  NAND2X1 U1776 ( .A(\mem<3><12> ), .B(n1281), .Y(n1791) );
  OAI21X1 U1777 ( .A(n145), .B(n1304), .C(n1791), .Y(n1898) );
  NAND2X1 U1778 ( .A(\mem<3><13> ), .B(n1281), .Y(n1792) );
  OAI21X1 U1779 ( .A(n145), .B(n1305), .C(n1792), .Y(n1897) );
  NAND2X1 U1780 ( .A(\mem<3><14> ), .B(n1281), .Y(n1793) );
  OAI21X1 U1781 ( .A(n145), .B(n1306), .C(n1793), .Y(n1896) );
  NAND2X1 U1782 ( .A(\mem<3><15> ), .B(n1281), .Y(n1794) );
  OAI21X1 U1783 ( .A(n145), .B(n1307), .C(n1794), .Y(n1895) );
  NAND2X1 U1784 ( .A(\mem<2><0> ), .B(n1282), .Y(n1796) );
  OAI21X1 U1785 ( .A(n149), .B(n1292), .C(n1796), .Y(n1894) );
  NAND2X1 U1786 ( .A(\mem<2><1> ), .B(n1282), .Y(n1797) );
  OAI21X1 U1787 ( .A(n149), .B(n1293), .C(n1797), .Y(n1893) );
  NAND2X1 U1788 ( .A(\mem<2><2> ), .B(n1282), .Y(n1798) );
  OAI21X1 U1789 ( .A(n149), .B(n1294), .C(n1798), .Y(n1892) );
  NAND2X1 U1790 ( .A(\mem<2><3> ), .B(n1282), .Y(n1799) );
  OAI21X1 U1791 ( .A(n149), .B(n1295), .C(n1799), .Y(n1891) );
  NAND2X1 U1792 ( .A(\mem<2><4> ), .B(n1282), .Y(n1800) );
  OAI21X1 U1793 ( .A(n149), .B(n1296), .C(n1800), .Y(n1890) );
  NAND2X1 U1794 ( .A(\mem<2><5> ), .B(n1282), .Y(n1801) );
  OAI21X1 U1795 ( .A(n149), .B(n1297), .C(n1801), .Y(n1889) );
  NAND2X1 U1796 ( .A(\mem<2><6> ), .B(n1282), .Y(n1802) );
  OAI21X1 U1797 ( .A(n149), .B(n1298), .C(n1802), .Y(n1888) );
  NAND2X1 U1798 ( .A(\mem<2><7> ), .B(n1282), .Y(n1803) );
  OAI21X1 U1799 ( .A(n149), .B(n1299), .C(n1803), .Y(n1887) );
  NAND2X1 U1800 ( .A(\mem<2><8> ), .B(n1283), .Y(n1804) );
  OAI21X1 U1801 ( .A(n149), .B(n1300), .C(n1804), .Y(n1886) );
  NAND2X1 U1802 ( .A(\mem<2><9> ), .B(n1283), .Y(n1805) );
  OAI21X1 U1803 ( .A(n149), .B(n1301), .C(n1805), .Y(n1885) );
  NAND2X1 U1804 ( .A(\mem<2><10> ), .B(n1283), .Y(n1806) );
  OAI21X1 U1805 ( .A(n149), .B(n1302), .C(n1806), .Y(n1884) );
  NAND2X1 U1806 ( .A(\mem<2><11> ), .B(n1283), .Y(n1807) );
  OAI21X1 U1807 ( .A(n149), .B(n1303), .C(n1807), .Y(n1883) );
  NAND2X1 U1808 ( .A(\mem<2><12> ), .B(n1283), .Y(n1808) );
  OAI21X1 U1809 ( .A(n149), .B(n1304), .C(n1808), .Y(n1882) );
  NAND2X1 U1810 ( .A(\mem<2><13> ), .B(n1283), .Y(n1809) );
  OAI21X1 U1811 ( .A(n149), .B(n1305), .C(n1809), .Y(n1881) );
  NAND2X1 U1812 ( .A(\mem<2><14> ), .B(n1283), .Y(n1810) );
  OAI21X1 U1813 ( .A(n149), .B(n1306), .C(n1810), .Y(n1880) );
  NAND2X1 U1814 ( .A(\mem<2><15> ), .B(n1283), .Y(n1811) );
  OAI21X1 U1815 ( .A(n149), .B(n1307), .C(n1811), .Y(n1879) );
  NAND2X1 U1816 ( .A(\mem<1><0> ), .B(n1284), .Y(n1813) );
  OAI21X1 U1817 ( .A(n153), .B(n1292), .C(n1813), .Y(n1878) );
  NAND2X1 U1818 ( .A(\mem<1><1> ), .B(n1284), .Y(n1814) );
  OAI21X1 U1819 ( .A(n153), .B(n1293), .C(n1814), .Y(n1877) );
  NAND2X1 U1820 ( .A(\mem<1><2> ), .B(n1284), .Y(n1815) );
  OAI21X1 U1821 ( .A(n153), .B(n1294), .C(n1815), .Y(n1876) );
  NAND2X1 U1822 ( .A(\mem<1><3> ), .B(n1284), .Y(n1816) );
  OAI21X1 U1823 ( .A(n153), .B(n1295), .C(n1816), .Y(n1875) );
  NAND2X1 U1824 ( .A(\mem<1><4> ), .B(n1284), .Y(n1817) );
  OAI21X1 U1825 ( .A(n153), .B(n1296), .C(n1817), .Y(n1874) );
  NAND2X1 U1826 ( .A(\mem<1><5> ), .B(n1284), .Y(n1818) );
  OAI21X1 U1827 ( .A(n153), .B(n1297), .C(n1818), .Y(n1873) );
  NAND2X1 U1828 ( .A(\mem<1><6> ), .B(n1284), .Y(n1819) );
  OAI21X1 U1829 ( .A(n153), .B(n1298), .C(n1819), .Y(n1872) );
  NAND2X1 U1830 ( .A(\mem<1><7> ), .B(n1284), .Y(n1820) );
  OAI21X1 U1831 ( .A(n153), .B(n1299), .C(n1820), .Y(n1871) );
  NAND2X1 U1832 ( .A(\mem<1><8> ), .B(n1285), .Y(n1821) );
  OAI21X1 U1833 ( .A(n153), .B(n1300), .C(n1821), .Y(n1870) );
  NAND2X1 U1834 ( .A(\mem<1><9> ), .B(n1285), .Y(n1822) );
  OAI21X1 U1835 ( .A(n153), .B(n1301), .C(n1822), .Y(n1869) );
  NAND2X1 U1836 ( .A(\mem<1><10> ), .B(n1285), .Y(n1823) );
  OAI21X1 U1837 ( .A(n153), .B(n1302), .C(n1823), .Y(n1868) );
  NAND2X1 U1838 ( .A(\mem<1><11> ), .B(n1285), .Y(n1824) );
  OAI21X1 U1839 ( .A(n153), .B(n1303), .C(n1824), .Y(n1867) );
  NAND2X1 U1840 ( .A(\mem<1><12> ), .B(n1285), .Y(n1825) );
  OAI21X1 U1841 ( .A(n153), .B(n1304), .C(n1825), .Y(n1866) );
  NAND2X1 U1842 ( .A(\mem<1><13> ), .B(n1285), .Y(n1826) );
  OAI21X1 U1843 ( .A(n153), .B(n1305), .C(n1826), .Y(n1865) );
  NAND2X1 U1844 ( .A(\mem<1><14> ), .B(n1285), .Y(n1827) );
  OAI21X1 U1845 ( .A(n153), .B(n1306), .C(n1827), .Y(n1864) );
  NAND2X1 U1846 ( .A(\mem<1><15> ), .B(n1285), .Y(n1828) );
  OAI21X1 U1847 ( .A(n153), .B(n1307), .C(n1828), .Y(n1863) );
  NAND2X1 U1848 ( .A(\mem<0><0> ), .B(n1286), .Y(n1831) );
  OAI21X1 U1849 ( .A(n37), .B(n1292), .C(n1831), .Y(n1862) );
  NAND2X1 U1850 ( .A(\mem<0><1> ), .B(n1286), .Y(n1832) );
  OAI21X1 U1851 ( .A(n37), .B(n1293), .C(n1832), .Y(n1861) );
  NAND2X1 U1852 ( .A(\mem<0><2> ), .B(n1286), .Y(n1833) );
  OAI21X1 U1853 ( .A(n37), .B(n1294), .C(n1833), .Y(n1860) );
  NAND2X1 U1854 ( .A(\mem<0><3> ), .B(n1286), .Y(n1834) );
  OAI21X1 U1855 ( .A(n37), .B(n1295), .C(n1834), .Y(n1859) );
  NAND2X1 U1856 ( .A(\mem<0><4> ), .B(n1286), .Y(n1835) );
  OAI21X1 U1857 ( .A(n37), .B(n1296), .C(n1835), .Y(n1858) );
  NAND2X1 U1858 ( .A(\mem<0><5> ), .B(n1286), .Y(n1836) );
  OAI21X1 U1859 ( .A(n37), .B(n1297), .C(n1836), .Y(n1857) );
  NAND2X1 U1860 ( .A(\mem<0><6> ), .B(n1286), .Y(n1837) );
  OAI21X1 U1861 ( .A(n37), .B(n1298), .C(n1837), .Y(n1856) );
  NAND2X1 U1862 ( .A(\mem<0><7> ), .B(n1286), .Y(n1838) );
  OAI21X1 U1863 ( .A(n37), .B(n1299), .C(n1838), .Y(n1855) );
  NAND2X1 U1864 ( .A(\mem<0><8> ), .B(n1287), .Y(n1839) );
  OAI21X1 U1865 ( .A(n37), .B(n1300), .C(n1839), .Y(n1854) );
  NAND2X1 U1866 ( .A(\mem<0><9> ), .B(n1287), .Y(n1840) );
  OAI21X1 U1867 ( .A(n37), .B(n1301), .C(n1840), .Y(n1853) );
  NAND2X1 U1868 ( .A(\mem<0><10> ), .B(n1287), .Y(n1841) );
  OAI21X1 U1869 ( .A(n37), .B(n1302), .C(n1841), .Y(n1852) );
  NAND2X1 U1870 ( .A(\mem<0><11> ), .B(n1287), .Y(n1842) );
  OAI21X1 U1871 ( .A(n37), .B(n1303), .C(n1842), .Y(n1851) );
  NAND2X1 U1872 ( .A(\mem<0><12> ), .B(n1287), .Y(n1843) );
  OAI21X1 U1873 ( .A(n37), .B(n1304), .C(n1843), .Y(n1850) );
  NAND2X1 U1874 ( .A(\mem<0><13> ), .B(n1287), .Y(n1844) );
  OAI21X1 U1875 ( .A(n37), .B(n1305), .C(n1844), .Y(n1849) );
  NAND2X1 U1876 ( .A(\mem<0><14> ), .B(n1287), .Y(n1845) );
  OAI21X1 U1877 ( .A(n37), .B(n1306), .C(n1845), .Y(n1848) );
  NAND2X1 U1878 ( .A(\mem<0><15> ), .B(n1287), .Y(n1846) );
  OAI21X1 U1879 ( .A(n37), .B(n1307), .C(n1846), .Y(n1847) );
endmodule


module memc_Size5_0 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n58, n59, n60, n61, n62, n63, n64, n66, n67, n68, n69, n70,
         n71, n74, n75, n76, n77, n78, n79, n82, n83, n84, n85, n86, n87, n88,
         n90, n91, n92, n93, n94, n95, n96, n98, n99, n100, n101, n102, n103,
         n106, n107, n108, n109, n110, n111, n112, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n130, n131, n132,
         n133, n134, n137, n138, n139, n140, n141, n142, n144, n145, n146,
         n147, n148, n149, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n165, n166, n167, n168, n169, n170,
         n171, n173, n175, n176, n177, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n189, n190, n191, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n230, n231, n232,
         n233, n234, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n251, n252, n253, n254, n255, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n267, n268, n269, n270, n271,
         n272, n274, n275, n276, n278, n279, n280, n281, n282, n283, n284,
         n285, n287, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n467, n469,
         n471, n473, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n814), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n815), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n816), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n817), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n818), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n819), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n820), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n821), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n822), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n823), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n824), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n825), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n826), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n827), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n828), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n829), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n830), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n831), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n832), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n833), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n834), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n835), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n836), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n837), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n838), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n839), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n840), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n841), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n842), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n843), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n844), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n845), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n846), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n847), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n848), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n849), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n850), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n851), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n852), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n853), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n854), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n855), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n856), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n857), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n858), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n859), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n860), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n861), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n862), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n863), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n864), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n865), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n866), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n867), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n868), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n869), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n870), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n871), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n872), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n873), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n874), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n875), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n876), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n877), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n878), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n879), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n880), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n881), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n882), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n883), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n884), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n885), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n886), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n887), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n888), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n889), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n890), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n891), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n892), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n893), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n894), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n895), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n896), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n897), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n898), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n899), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n900), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n901), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n902), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n903), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n904), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n905), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n906), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n907), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n908), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n909), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n910), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n911), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n912), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n913), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n914), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n915), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n916), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n917), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n918), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n919), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n920), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n921), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n922), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n923), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n924), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n925), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n926), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n927), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n928), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n929), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n930), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n931), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n932), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n933), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n934), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n935), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n936), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n937), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n938), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n939), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n940), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n941), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n942), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n943), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n944), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n945), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n946), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n947), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n948), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n949), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n950), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n951), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n952), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n953), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n954), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n955), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n956), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n957), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n958), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n959), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n960), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n961), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n962), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n963), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n964), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n965), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n966), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n967), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n968), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n969), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n970), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n971), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n972), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n973), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(write), .B(n653), .Y(n1010) );
  OAI21X1 U50 ( .A(n561), .B(n632), .C(n463), .Y(n973) );
  OAI21X1 U52 ( .A(n561), .B(n631), .C(n461), .Y(n972) );
  OAI21X1 U54 ( .A(n561), .B(n630), .C(n459), .Y(n971) );
  OAI21X1 U56 ( .A(n561), .B(n629), .C(n457), .Y(n970) );
  OAI21X1 U58 ( .A(n561), .B(n628), .C(n1011), .Y(n969) );
  NAND2X1 U59 ( .A(\mem<31><4> ), .B(n559), .Y(n1011) );
  OAI21X1 U62 ( .A(n632), .B(n623), .C(n455), .Y(n968) );
  OAI21X1 U64 ( .A(n631), .B(n623), .C(n453), .Y(n967) );
  OAI21X1 U66 ( .A(n630), .B(n623), .C(n451), .Y(n966) );
  OAI21X1 U68 ( .A(n629), .B(n623), .C(n449), .Y(n965) );
  OAI21X1 U70 ( .A(n628), .B(n623), .C(n287), .Y(n964) );
  OAI21X1 U74 ( .A(n632), .B(n621), .C(n284), .Y(n963) );
  OAI21X1 U76 ( .A(n631), .B(n621), .C(n282), .Y(n962) );
  OAI21X1 U78 ( .A(n630), .B(n621), .C(n280), .Y(n961) );
  OAI21X1 U80 ( .A(n629), .B(n621), .C(n278), .Y(n960) );
  OAI21X1 U82 ( .A(n628), .B(n621), .C(n1007), .Y(n959) );
  NAND2X1 U83 ( .A(\mem<29><4> ), .B(n555), .Y(n1007) );
  OAI21X1 U86 ( .A(n632), .B(n619), .C(n275), .Y(n958) );
  OAI21X1 U88 ( .A(n631), .B(n619), .C(n272), .Y(n957) );
  OAI21X1 U90 ( .A(n630), .B(n619), .C(n270), .Y(n956) );
  OAI21X1 U92 ( .A(n629), .B(n619), .C(n268), .Y(n955) );
  OAI21X1 U94 ( .A(n628), .B(n619), .C(n1005), .Y(n954) );
  NAND2X1 U95 ( .A(\mem<28><4> ), .B(n553), .Y(n1005) );
  OAI21X1 U98 ( .A(n632), .B(n617), .C(n265), .Y(n953) );
  OAI21X1 U100 ( .A(n631), .B(n617), .C(n263), .Y(n952) );
  OAI21X1 U102 ( .A(n630), .B(n617), .C(n261), .Y(n951) );
  OAI21X1 U104 ( .A(n629), .B(n617), .C(n259), .Y(n950) );
  OAI21X1 U106 ( .A(n628), .B(n617), .C(n257), .Y(n949) );
  OAI21X1 U110 ( .A(n632), .B(n615), .C(n254), .Y(n948) );
  OAI21X1 U112 ( .A(n631), .B(n615), .C(n252), .Y(n947) );
  OAI21X1 U114 ( .A(n630), .B(n615), .C(n486), .Y(n946) );
  OAI21X1 U116 ( .A(n629), .B(n615), .C(n248), .Y(n945) );
  OAI21X1 U118 ( .A(n628), .B(n615), .C(n246), .Y(n944) );
  OAI21X1 U122 ( .A(n632), .B(n613), .C(n244), .Y(n943) );
  OAI21X1 U124 ( .A(n631), .B(n613), .C(n242), .Y(n942) );
  OAI21X1 U126 ( .A(n630), .B(n613), .C(n240), .Y(n941) );
  OAI21X1 U128 ( .A(n629), .B(n613), .C(n238), .Y(n940) );
  OAI21X1 U130 ( .A(n628), .B(n613), .C(n1001), .Y(n939) );
  NAND2X1 U131 ( .A(\mem<25><4> ), .B(n547), .Y(n1001) );
  OAI21X1 U134 ( .A(n632), .B(n611), .C(n234), .Y(n938) );
  OAI21X1 U136 ( .A(n631), .B(n611), .C(n232), .Y(n937) );
  OAI21X1 U138 ( .A(n630), .B(n611), .C(n484), .Y(n936) );
  OAI21X1 U140 ( .A(n629), .B(n611), .C(n230), .Y(n935) );
  OAI21X1 U142 ( .A(n628), .B(n611), .C(n227), .Y(n934) );
  NAND3X1 U146 ( .A(n649), .B(n997), .C(n651), .Y(n998) );
  OAI21X1 U147 ( .A(n632), .B(n609), .C(n225), .Y(n933) );
  OAI21X1 U149 ( .A(n631), .B(n609), .C(n223), .Y(n932) );
  OAI21X1 U151 ( .A(n630), .B(n609), .C(n221), .Y(n931) );
  OAI21X1 U153 ( .A(n629), .B(n609), .C(n219), .Y(n930) );
  OAI21X1 U155 ( .A(n628), .B(n609), .C(n996), .Y(n929) );
  NAND2X1 U156 ( .A(\mem<23><4> ), .B(n543), .Y(n996) );
  OAI21X1 U159 ( .A(n632), .B(n607), .C(n217), .Y(n928) );
  OAI21X1 U161 ( .A(n631), .B(n607), .C(n215), .Y(n927) );
  OAI21X1 U163 ( .A(n630), .B(n607), .C(n213), .Y(n926) );
  OAI21X1 U165 ( .A(n629), .B(n607), .C(n211), .Y(n925) );
  OAI21X1 U167 ( .A(n628), .B(n607), .C(n995), .Y(n924) );
  NAND2X1 U168 ( .A(\mem<22><4> ), .B(n541), .Y(n995) );
  OAI21X1 U171 ( .A(n632), .B(n605), .C(n209), .Y(n923) );
  OAI21X1 U173 ( .A(n631), .B(n605), .C(n206), .Y(n922) );
  OAI21X1 U175 ( .A(n630), .B(n605), .C(n204), .Y(n921) );
  OAI21X1 U177 ( .A(n629), .B(n605), .C(n994), .Y(n920) );
  NAND2X1 U178 ( .A(\mem<21><3> ), .B(n539), .Y(n994) );
  OAI21X1 U179 ( .A(n628), .B(n605), .C(n993), .Y(n919) );
  NAND2X1 U180 ( .A(\mem<21><4> ), .B(n539), .Y(n993) );
  OAI21X1 U183 ( .A(n632), .B(n603), .C(n202), .Y(n918) );
  OAI21X1 U185 ( .A(n631), .B(n603), .C(n200), .Y(n917) );
  OAI21X1 U187 ( .A(n630), .B(n603), .C(n198), .Y(n916) );
  OAI21X1 U189 ( .A(n629), .B(n603), .C(n196), .Y(n915) );
  OAI21X1 U191 ( .A(n628), .B(n603), .C(n992), .Y(n914) );
  NAND2X1 U192 ( .A(\mem<20><4> ), .B(n537), .Y(n992) );
  OAI21X1 U195 ( .A(n632), .B(n601), .C(n194), .Y(n913) );
  OAI21X1 U197 ( .A(n631), .B(n601), .C(n191), .Y(n912) );
  OAI21X1 U199 ( .A(n630), .B(n601), .C(n189), .Y(n911) );
  OAI21X1 U201 ( .A(n629), .B(n601), .C(n186), .Y(n910) );
  OAI21X1 U203 ( .A(n628), .B(n601), .C(n991), .Y(n909) );
  NAND2X1 U204 ( .A(\mem<19><4> ), .B(n535), .Y(n991) );
  OAI21X1 U207 ( .A(n632), .B(n598), .C(n184), .Y(n908) );
  OAI21X1 U209 ( .A(n631), .B(n598), .C(n182), .Y(n907) );
  OAI21X1 U211 ( .A(n630), .B(n598), .C(n482), .Y(n906) );
  OAI21X1 U213 ( .A(n629), .B(n598), .C(n180), .Y(n905) );
  OAI21X1 U215 ( .A(n628), .B(n598), .C(n177), .Y(n904) );
  OAI21X1 U219 ( .A(n632), .B(n597), .C(n175), .Y(n903) );
  OAI21X1 U221 ( .A(n631), .B(n597), .C(n171), .Y(n902) );
  OAI21X1 U223 ( .A(n630), .B(n597), .C(n169), .Y(n901) );
  OAI21X1 U225 ( .A(n629), .B(n597), .C(n167), .Y(n900) );
  OAI21X1 U227 ( .A(n628), .B(n597), .C(n990), .Y(n899) );
  NAND2X1 U228 ( .A(\mem<17><4> ), .B(n531), .Y(n990) );
  OAI21X1 U231 ( .A(n632), .B(n595), .C(n165), .Y(n898) );
  OAI21X1 U233 ( .A(n631), .B(n595), .C(n162), .Y(n897) );
  OAI21X1 U235 ( .A(n630), .B(n595), .C(n160), .Y(n896) );
  OAI21X1 U237 ( .A(n629), .B(n595), .C(n158), .Y(n895) );
  OAI21X1 U239 ( .A(n628), .B(n595), .C(n156), .Y(n894) );
  NAND3X1 U243 ( .A(n997), .B(n650), .C(n651), .Y(n989) );
  OAI21X1 U244 ( .A(n632), .B(n593), .C(n988), .Y(n893) );
  NAND2X1 U245 ( .A(\mem<15><0> ), .B(n527), .Y(n988) );
  OAI21X1 U246 ( .A(n631), .B(n593), .C(n154), .Y(n892) );
  OAI21X1 U248 ( .A(n630), .B(n593), .C(n152), .Y(n891) );
  OAI21X1 U250 ( .A(n629), .B(n593), .C(n987), .Y(n890) );
  NAND2X1 U251 ( .A(\mem<15><3> ), .B(n527), .Y(n987) );
  OAI21X1 U252 ( .A(n628), .B(n593), .C(n149), .Y(n889) );
  OAI21X1 U256 ( .A(n632), .B(n591), .C(n147), .Y(n888) );
  OAI21X1 U258 ( .A(n631), .B(n591), .C(n145), .Y(n887) );
  OAI21X1 U260 ( .A(n630), .B(n591), .C(n142), .Y(n886) );
  OAI21X1 U262 ( .A(n629), .B(n591), .C(n140), .Y(n885) );
  OAI21X1 U264 ( .A(n628), .B(n591), .C(n138), .Y(n884) );
  OAI21X1 U268 ( .A(n632), .B(n589), .C(n986), .Y(n883) );
  NAND2X1 U269 ( .A(\mem<13><0> ), .B(n523), .Y(n986) );
  OAI21X1 U270 ( .A(n631), .B(n589), .C(n134), .Y(n882) );
  OAI21X1 U272 ( .A(n630), .B(n589), .C(n132), .Y(n881) );
  OAI21X1 U274 ( .A(n629), .B(n589), .C(n985), .Y(n880) );
  NAND2X1 U275 ( .A(\mem<13><3> ), .B(n523), .Y(n985) );
  OAI21X1 U276 ( .A(n628), .B(n589), .C(n130), .Y(n879) );
  OAI21X1 U280 ( .A(n632), .B(n586), .C(n127), .Y(n878) );
  OAI21X1 U282 ( .A(n631), .B(n586), .C(n125), .Y(n877) );
  OAI21X1 U284 ( .A(n630), .B(n586), .C(n123), .Y(n876) );
  OAI21X1 U286 ( .A(n629), .B(n586), .C(n120), .Y(n875) );
  OAI21X1 U288 ( .A(n628), .B(n586), .C(n118), .Y(n874) );
  OAI21X1 U292 ( .A(n632), .B(n584), .C(n116), .Y(n873) );
  OAI21X1 U294 ( .A(n631), .B(n584), .C(n111), .Y(n872) );
  OAI21X1 U296 ( .A(n630), .B(n584), .C(n109), .Y(n871) );
  OAI21X1 U298 ( .A(n629), .B(n584), .C(n107), .Y(n870) );
  OAI21X1 U300 ( .A(n628), .B(n584), .C(n984), .Y(n869) );
  NAND2X1 U301 ( .A(\mem<11><4> ), .B(n519), .Y(n984) );
  OAI21X1 U304 ( .A(n632), .B(n582), .C(n103), .Y(n868) );
  OAI21X1 U306 ( .A(n631), .B(n582), .C(n480), .Y(n867) );
  OAI21X1 U308 ( .A(n630), .B(n582), .C(n101), .Y(n866) );
  OAI21X1 U310 ( .A(n629), .B(n582), .C(n99), .Y(n865) );
  OAI21X1 U312 ( .A(n628), .B(n582), .C(n96), .Y(n864) );
  OAI21X1 U316 ( .A(n632), .B(n581), .C(n94), .Y(n863) );
  OAI21X1 U318 ( .A(n631), .B(n581), .C(n92), .Y(n862) );
  OAI21X1 U320 ( .A(n630), .B(n581), .C(n90), .Y(n861) );
  OAI21X1 U322 ( .A(n629), .B(n581), .C(n87), .Y(n860) );
  OAI21X1 U324 ( .A(n628), .B(n581), .C(n85), .Y(n859) );
  OAI21X1 U328 ( .A(n632), .B(n579), .C(n83), .Y(n858) );
  OAI21X1 U330 ( .A(n631), .B(n579), .C(n79), .Y(n857) );
  OAI21X1 U332 ( .A(n630), .B(n579), .C(n77), .Y(n856) );
  OAI21X1 U334 ( .A(n629), .B(n579), .C(n75), .Y(n855) );
  OAI21X1 U336 ( .A(n628), .B(n579), .C(n71), .Y(n854) );
  NAND3X1 U340 ( .A(n997), .B(n652), .C(n649), .Y(n983) );
  OAI21X1 U341 ( .A(n632), .B(n577), .C(n69), .Y(n853) );
  OAI21X1 U343 ( .A(n631), .B(n577), .C(n67), .Y(n852) );
  OAI21X1 U345 ( .A(n630), .B(n577), .C(n64), .Y(n851) );
  OAI21X1 U347 ( .A(n629), .B(n577), .C(n982), .Y(n850) );
  NAND2X1 U348 ( .A(\mem<7><3> ), .B(n511), .Y(n982) );
  OAI21X1 U349 ( .A(n628), .B(n577), .C(n981), .Y(n849) );
  NAND2X1 U350 ( .A(\mem<7><4> ), .B(n511), .Y(n981) );
  NOR3X1 U353 ( .A(n645), .B(n640), .C(n648), .Y(n1009) );
  OAI21X1 U354 ( .A(n632), .B(n575), .C(n62), .Y(n848) );
  OAI21X1 U356 ( .A(n631), .B(n575), .C(n60), .Y(n847) );
  OAI21X1 U358 ( .A(n630), .B(n575), .C(n58), .Y(n846) );
  OAI21X1 U360 ( .A(n629), .B(n575), .C(n53), .Y(n845) );
  OAI21X1 U362 ( .A(n628), .B(n575), .C(n51), .Y(n844) );
  NOR3X1 U366 ( .A(n646), .B(n636), .C(n648), .Y(n1008) );
  OAI21X1 U367 ( .A(n632), .B(n573), .C(n49), .Y(n843) );
  OAI21X1 U369 ( .A(n631), .B(n573), .C(n47), .Y(n842) );
  OAI21X1 U371 ( .A(n630), .B(n573), .C(n45), .Y(n841) );
  OAI21X1 U373 ( .A(n629), .B(n573), .C(n980), .Y(n840) );
  NAND2X1 U374 ( .A(\mem<5><3> ), .B(n507), .Y(n980) );
  OAI21X1 U375 ( .A(n628), .B(n573), .C(n979), .Y(n839) );
  NAND2X1 U376 ( .A(\mem<5><4> ), .B(n507), .Y(n979) );
  NOR3X1 U379 ( .A(n625), .B(n644), .C(n648), .Y(n1006) );
  OAI21X1 U380 ( .A(n632), .B(n570), .C(n43), .Y(n838) );
  OAI21X1 U382 ( .A(n631), .B(n570), .C(n41), .Y(n837) );
  OAI21X1 U384 ( .A(n630), .B(n570), .C(n39), .Y(n836) );
  OAI21X1 U386 ( .A(n629), .B(n570), .C(n978), .Y(n835) );
  NAND2X1 U387 ( .A(\mem<4><3> ), .B(n505), .Y(n978) );
  OAI21X1 U388 ( .A(n628), .B(n570), .C(n37), .Y(n834) );
  NOR3X1 U392 ( .A(n633), .B(n644), .C(n464), .Y(n1004) );
  OAI21X1 U393 ( .A(n632), .B(n568), .C(n35), .Y(n833) );
  OAI21X1 U395 ( .A(n631), .B(n568), .C(n33), .Y(n832) );
  OAI21X1 U397 ( .A(n630), .B(n568), .C(n31), .Y(n831) );
  OAI21X1 U399 ( .A(n629), .B(n568), .C(n29), .Y(n830) );
  OAI21X1 U401 ( .A(n628), .B(n568), .C(n27), .Y(n829) );
  NOR3X1 U405 ( .A(n626), .B(n647), .C(n646), .Y(n1003) );
  OAI21X1 U406 ( .A(n632), .B(n566), .C(n977), .Y(n828) );
  NAND2X1 U407 ( .A(\mem<2><0> ), .B(n501), .Y(n977) );
  OAI21X1 U408 ( .A(n631), .B(n566), .C(n478), .Y(n827) );
  OAI21X1 U410 ( .A(n630), .B(n566), .C(n25), .Y(n826) );
  OAI21X1 U412 ( .A(n629), .B(n566), .C(n23), .Y(n825) );
  OAI21X1 U414 ( .A(n628), .B(n566), .C(n21), .Y(n824) );
  NOR3X1 U418 ( .A(n2), .B(n647), .C(n646), .Y(n1002) );
  OAI21X1 U419 ( .A(n632), .B(n565), .C(n976), .Y(n823) );
  NAND2X1 U420 ( .A(\mem<1><0> ), .B(n499), .Y(n976) );
  OAI21X1 U421 ( .A(n631), .B(n565), .C(n19), .Y(n822) );
  OAI21X1 U423 ( .A(n630), .B(n565), .C(n17), .Y(n821) );
  OAI21X1 U425 ( .A(n629), .B(n565), .C(n975), .Y(n820) );
  NAND2X1 U426 ( .A(\mem<1><3> ), .B(n499), .Y(n975) );
  OAI21X1 U427 ( .A(n628), .B(n565), .C(n15), .Y(n819) );
  NOR3X1 U431 ( .A(n644), .B(n647), .C(n639), .Y(n1000) );
  OAI21X1 U432 ( .A(n632), .B(n563), .C(n13), .Y(n818) );
  OAI21X1 U435 ( .A(n631), .B(n563), .C(n476), .Y(n817) );
  OAI21X1 U438 ( .A(n630), .B(n563), .C(n11), .Y(n816) );
  OAI21X1 U441 ( .A(n629), .B(n563), .C(n9), .Y(n815) );
  OAI21X1 U444 ( .A(n628), .B(n563), .C(n7), .Y(n814) );
  NOR3X1 U448 ( .A(n644), .B(n647), .C(n635), .Y(n999) );
  NAND3X1 U449 ( .A(n650), .B(n652), .C(n997), .Y(n974) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n997) );
  INVX1 U3 ( .A(n652), .Y(n651) );
  INVX1 U4 ( .A(n638), .Y(n626) );
  INVX1 U5 ( .A(n641), .Y(n3) );
  INVX1 U6 ( .A(n649), .Y(n1) );
  INVX1 U7 ( .A(n467), .Y(\data_out<1> ) );
  OR2X1 U8 ( .A(n715), .B(n808), .Y(n467) );
  INVX1 U9 ( .A(n469), .Y(\data_out<2> ) );
  OR2X1 U10 ( .A(n746), .B(n808), .Y(n469) );
  AND2X1 U11 ( .A(\mem<31><0> ), .B(n559), .Y(n462) );
  AND2X1 U12 ( .A(\mem<31><1> ), .B(n559), .Y(n460) );
  AND2X1 U13 ( .A(\mem<30><4> ), .B(n557), .Y(n285) );
  AND2X1 U14 ( .A(\mem<29><1> ), .B(n555), .Y(n281) );
  AND2X1 U15 ( .A(\mem<28><0> ), .B(n553), .Y(n274) );
  AND2X1 U16 ( .A(\mem<27><3> ), .B(n551), .Y(n258) );
  AND2X1 U17 ( .A(\mem<27><4> ), .B(n551), .Y(n255) );
  AND2X1 U18 ( .A(\mem<25><3> ), .B(n547), .Y(n237) );
  AND2X1 U19 ( .A(\mem<23><3> ), .B(n543), .Y(n218) );
  AND2X1 U20 ( .A(\mem<20><2> ), .B(n537), .Y(n197) );
  AND2X1 U21 ( .A(\mem<20><3> ), .B(n537), .Y(n195) );
  AND2X1 U22 ( .A(\mem<19><0> ), .B(n535), .Y(n193) );
  AND2X1 U23 ( .A(\mem<19><1> ), .B(n535), .Y(n190) );
  AND2X1 U24 ( .A(\mem<17><0> ), .B(n531), .Y(n173) );
  AND2X1 U25 ( .A(\mem<17><1> ), .B(n531), .Y(n170) );
  AND2X1 U26 ( .A(\mem<17><3> ), .B(n531), .Y(n166) );
  AND2X1 U27 ( .A(\mem<16><4> ), .B(n529), .Y(n155) );
  AND2X1 U28 ( .A(\mem<15><2> ), .B(n527), .Y(n151) );
  AND2X1 U29 ( .A(\mem<15><4> ), .B(n527), .Y(n148) );
  AND2X1 U30 ( .A(\mem<14><0> ), .B(n525), .Y(n146) );
  AND2X1 U31 ( .A(\mem<14><3> ), .B(n525), .Y(n139) );
  AND2X1 U32 ( .A(\mem<14><4> ), .B(n525), .Y(n137) );
  AND2X1 U33 ( .A(\mem<13><2> ), .B(n523), .Y(n131) );
  AND2X1 U34 ( .A(\mem<13><4> ), .B(n523), .Y(n128) );
  AND2X1 U35 ( .A(\mem<12><0> ), .B(n521), .Y(n126) );
  AND2X1 U36 ( .A(\mem<12><3> ), .B(n521), .Y(n119) );
  AND2X1 U37 ( .A(\mem<12><4> ), .B(n521), .Y(n117) );
  AND2X1 U38 ( .A(\mem<11><3> ), .B(n519), .Y(n106) );
  AND2X1 U39 ( .A(\mem<10><0> ), .B(n517), .Y(n102) );
  AND2X1 U40 ( .A(\mem<10><4> ), .B(n517), .Y(n95) );
  AND2X1 U41 ( .A(\mem<9><0> ), .B(n515), .Y(n93) );
  AND2X1 U42 ( .A(\mem<9><3> ), .B(n515), .Y(n86) );
  AND2X1 U43 ( .A(\mem<9><4> ), .B(n515), .Y(n84) );
  AND2X1 U44 ( .A(\mem<8><4> ), .B(n513), .Y(n70) );
  AND2X1 U45 ( .A(\mem<7><0> ), .B(n511), .Y(n68) );
  AND2X1 U46 ( .A(\mem<7><2> ), .B(n511), .Y(n63) );
  AND2X1 U47 ( .A(\mem<6><3> ), .B(n509), .Y(n52) );
  AND2X1 U48 ( .A(\mem<6><4> ), .B(n509), .Y(n50) );
  AND2X1 U49 ( .A(\mem<5><0> ), .B(n507), .Y(n48) );
  AND2X1 U51 ( .A(\mem<5><2> ), .B(n507), .Y(n44) );
  AND2X1 U53 ( .A(\mem<4><2> ), .B(n505), .Y(n38) );
  AND2X1 U55 ( .A(\mem<4><4> ), .B(n505), .Y(n36) );
  AND2X1 U57 ( .A(\mem<3><0> ), .B(n503), .Y(n34) );
  AND2X1 U60 ( .A(\mem<3><3> ), .B(n503), .Y(n28) );
  AND2X1 U61 ( .A(\mem<3><4> ), .B(n503), .Y(n26) );
  AND2X1 U63 ( .A(\mem<2><4> ), .B(n501), .Y(n20) );
  AND2X1 U65 ( .A(\mem<1><2> ), .B(n499), .Y(n16) );
  AND2X1 U67 ( .A(\mem<1><4> ), .B(n499), .Y(n14) );
  AND2X1 U69 ( .A(\mem<0><0> ), .B(n497), .Y(n12) );
  AND2X1 U71 ( .A(\mem<0><3> ), .B(n497), .Y(n8) );
  AND2X1 U72 ( .A(\mem<0><4> ), .B(n497), .Y(n6) );
  INVX4 U73 ( .A(N12), .Y(n4) );
  INVX1 U75 ( .A(N12), .Y(n5) );
  INVX1 U77 ( .A(rst), .Y(n653) );
  INVX1 U79 ( .A(n647), .Y(n464) );
  MUX2X1 U81 ( .B(\mem<11><4> ), .A(\mem<10><4> ), .S(n639), .Y(n784) );
  MUX2X1 U84 ( .B(n790), .A(n791), .S(n1), .Y(n807) );
  MUX2X1 U85 ( .B(n806), .A(n807), .S(n652), .Y(n809) );
  OR2X1 U87 ( .A(n809), .B(n808), .Y(n473) );
  MUX2X1 U89 ( .B(n686), .A(n685), .S(N11), .Y(n690) );
  INVX8 U91 ( .A(n627), .Y(n2) );
  MUX2X1 U93 ( .B(n691), .A(n692), .S(n3), .Y(n696) );
  MUX2X1 U96 ( .B(\mem<5><1> ), .A(\mem<4><1> ), .S(n634), .Y(n688) );
  MUX2X1 U97 ( .B(n703), .A(n704), .S(n4), .Y(n712) );
  MUX2X1 U99 ( .B(n689), .A(n690), .S(n4), .Y(n698) );
  MUX2X1 U101 ( .B(n695), .A(n696), .S(n5), .Y(n697) );
  INVX1 U103 ( .A(n6), .Y(n7) );
  INVX1 U105 ( .A(n8), .Y(n9) );
  AND2X2 U107 ( .A(\mem<0><2> ), .B(n497), .Y(n10) );
  INVX1 U108 ( .A(n10), .Y(n11) );
  INVX1 U109 ( .A(n12), .Y(n13) );
  INVX1 U111 ( .A(n14), .Y(n15) );
  INVX1 U113 ( .A(n16), .Y(n17) );
  AND2X2 U115 ( .A(\mem<1><1> ), .B(n499), .Y(n18) );
  INVX1 U117 ( .A(n18), .Y(n19) );
  INVX1 U119 ( .A(n20), .Y(n21) );
  AND2X2 U120 ( .A(\mem<2><3> ), .B(n501), .Y(n22) );
  INVX1 U121 ( .A(n22), .Y(n23) );
  AND2X2 U123 ( .A(\mem<2><2> ), .B(n501), .Y(n24) );
  INVX1 U125 ( .A(n24), .Y(n25) );
  INVX1 U127 ( .A(n26), .Y(n27) );
  INVX1 U129 ( .A(n28), .Y(n29) );
  AND2X2 U132 ( .A(\mem<3><2> ), .B(n503), .Y(n30) );
  INVX1 U133 ( .A(n30), .Y(n31) );
  AND2X2 U135 ( .A(\mem<3><1> ), .B(n503), .Y(n32) );
  INVX1 U137 ( .A(n32), .Y(n33) );
  INVX1 U139 ( .A(n34), .Y(n35) );
  INVX1 U141 ( .A(n36), .Y(n37) );
  INVX1 U143 ( .A(n38), .Y(n39) );
  AND2X2 U144 ( .A(\mem<4><1> ), .B(n505), .Y(n40) );
  INVX1 U145 ( .A(n40), .Y(n41) );
  AND2X2 U148 ( .A(\mem<4><0> ), .B(n505), .Y(n42) );
  INVX1 U150 ( .A(n42), .Y(n43) );
  INVX1 U152 ( .A(n44), .Y(n45) );
  AND2X2 U154 ( .A(\mem<5><1> ), .B(n507), .Y(n46) );
  INVX1 U157 ( .A(n46), .Y(n47) );
  INVX1 U158 ( .A(n48), .Y(n49) );
  INVX1 U160 ( .A(n50), .Y(n51) );
  INVX1 U162 ( .A(n52), .Y(n53) );
  AND2X2 U164 ( .A(\mem<6><2> ), .B(n509), .Y(n54) );
  INVX1 U166 ( .A(n54), .Y(n58) );
  AND2X2 U169 ( .A(\mem<6><1> ), .B(n509), .Y(n59) );
  INVX1 U170 ( .A(n59), .Y(n60) );
  AND2X2 U172 ( .A(\mem<6><0> ), .B(n509), .Y(n61) );
  INVX1 U174 ( .A(n61), .Y(n62) );
  INVX1 U176 ( .A(n63), .Y(n64) );
  AND2X2 U181 ( .A(\mem<7><1> ), .B(n511), .Y(n66) );
  INVX1 U182 ( .A(n66), .Y(n67) );
  INVX1 U184 ( .A(n68), .Y(n69) );
  INVX1 U186 ( .A(n70), .Y(n71) );
  AND2X2 U188 ( .A(\mem<8><3> ), .B(n513), .Y(n74) );
  INVX1 U190 ( .A(n74), .Y(n75) );
  AND2X2 U193 ( .A(\mem<8><2> ), .B(n513), .Y(n76) );
  INVX1 U194 ( .A(n76), .Y(n77) );
  AND2X2 U196 ( .A(\mem<8><1> ), .B(n513), .Y(n78) );
  INVX1 U198 ( .A(n78), .Y(n79) );
  AND2X2 U200 ( .A(\mem<8><0> ), .B(n513), .Y(n82) );
  INVX1 U202 ( .A(n82), .Y(n83) );
  INVX1 U205 ( .A(n84), .Y(n85) );
  INVX1 U206 ( .A(n86), .Y(n87) );
  AND2X2 U208 ( .A(\mem<9><2> ), .B(n515), .Y(n88) );
  INVX1 U210 ( .A(n88), .Y(n90) );
  AND2X2 U212 ( .A(\mem<9><1> ), .B(n515), .Y(n91) );
  INVX1 U214 ( .A(n91), .Y(n92) );
  INVX1 U216 ( .A(n93), .Y(n94) );
  INVX1 U217 ( .A(n95), .Y(n96) );
  AND2X2 U218 ( .A(\mem<10><3> ), .B(n517), .Y(n98) );
  INVX1 U220 ( .A(n98), .Y(n99) );
  AND2X2 U222 ( .A(\mem<10><2> ), .B(n517), .Y(n100) );
  INVX1 U224 ( .A(n100), .Y(n101) );
  INVX1 U226 ( .A(n102), .Y(n103) );
  INVX1 U229 ( .A(n106), .Y(n107) );
  AND2X2 U230 ( .A(\mem<11><2> ), .B(n519), .Y(n108) );
  INVX1 U232 ( .A(n108), .Y(n109) );
  AND2X2 U234 ( .A(\mem<11><1> ), .B(n519), .Y(n110) );
  INVX1 U236 ( .A(n110), .Y(n111) );
  AND2X2 U238 ( .A(\mem<11><0> ), .B(n519), .Y(n112) );
  INVX1 U240 ( .A(n112), .Y(n116) );
  INVX1 U241 ( .A(n117), .Y(n118) );
  INVX1 U242 ( .A(n119), .Y(n120) );
  AND2X2 U247 ( .A(\mem<12><2> ), .B(n521), .Y(n121) );
  INVX1 U249 ( .A(n121), .Y(n123) );
  AND2X2 U253 ( .A(\mem<12><1> ), .B(n521), .Y(n124) );
  INVX1 U254 ( .A(n124), .Y(n125) );
  INVX1 U255 ( .A(n126), .Y(n127) );
  INVX1 U257 ( .A(n128), .Y(n130) );
  INVX1 U259 ( .A(n131), .Y(n132) );
  AND2X2 U261 ( .A(\mem<13><1> ), .B(n523), .Y(n133) );
  INVX1 U263 ( .A(n133), .Y(n134) );
  INVX1 U265 ( .A(n137), .Y(n138) );
  INVX1 U266 ( .A(n139), .Y(n140) );
  AND2X2 U267 ( .A(\mem<14><2> ), .B(n525), .Y(n141) );
  INVX1 U271 ( .A(n141), .Y(n142) );
  AND2X2 U273 ( .A(\mem<14><1> ), .B(n525), .Y(n144) );
  INVX1 U277 ( .A(n144), .Y(n145) );
  INVX1 U278 ( .A(n146), .Y(n147) );
  INVX1 U279 ( .A(n148), .Y(n149) );
  INVX1 U281 ( .A(n151), .Y(n152) );
  AND2X2 U283 ( .A(\mem<15><1> ), .B(n527), .Y(n153) );
  INVX1 U285 ( .A(n153), .Y(n154) );
  INVX1 U287 ( .A(n155), .Y(n156) );
  AND2X2 U289 ( .A(\mem<16><3> ), .B(n529), .Y(n157) );
  INVX1 U290 ( .A(n157), .Y(n158) );
  AND2X2 U291 ( .A(\mem<16><2> ), .B(n529), .Y(n159) );
  INVX1 U293 ( .A(n159), .Y(n160) );
  AND2X2 U295 ( .A(\mem<16><1> ), .B(n529), .Y(n161) );
  INVX1 U297 ( .A(n161), .Y(n162) );
  AND2X2 U299 ( .A(\mem<16><0> ), .B(n529), .Y(n163) );
  INVX1 U302 ( .A(n163), .Y(n165) );
  INVX1 U303 ( .A(n166), .Y(n167) );
  AND2X2 U305 ( .A(\mem<17><2> ), .B(n531), .Y(n168) );
  INVX1 U307 ( .A(n168), .Y(n169) );
  INVX1 U309 ( .A(n170), .Y(n171) );
  INVX1 U311 ( .A(n173), .Y(n175) );
  AND2X2 U313 ( .A(\mem<18><4> ), .B(n533), .Y(n176) );
  INVX1 U314 ( .A(n176), .Y(n177) );
  AND2X2 U315 ( .A(\mem<18><3> ), .B(n533), .Y(n179) );
  INVX1 U317 ( .A(n179), .Y(n180) );
  AND2X2 U319 ( .A(\mem<18><1> ), .B(n533), .Y(n181) );
  INVX1 U321 ( .A(n181), .Y(n182) );
  AND2X2 U323 ( .A(\mem<18><0> ), .B(n533), .Y(n183) );
  INVX1 U325 ( .A(n183), .Y(n184) );
  AND2X2 U326 ( .A(\mem<19><3> ), .B(n535), .Y(n185) );
  INVX1 U327 ( .A(n185), .Y(n186) );
  AND2X2 U329 ( .A(\mem<19><2> ), .B(n535), .Y(n187) );
  INVX1 U331 ( .A(n187), .Y(n189) );
  INVX1 U333 ( .A(n190), .Y(n191) );
  INVX1 U335 ( .A(n193), .Y(n194) );
  INVX1 U337 ( .A(n195), .Y(n196) );
  INVX1 U338 ( .A(n197), .Y(n198) );
  AND2X2 U339 ( .A(\mem<20><1> ), .B(n537), .Y(n199) );
  INVX1 U342 ( .A(n199), .Y(n200) );
  AND2X2 U344 ( .A(\mem<20><0> ), .B(n537), .Y(n201) );
  INVX1 U346 ( .A(n201), .Y(n202) );
  AND2X2 U351 ( .A(\mem<21><2> ), .B(n539), .Y(n203) );
  INVX1 U352 ( .A(n203), .Y(n204) );
  AND2X2 U355 ( .A(\mem<21><1> ), .B(n539), .Y(n205) );
  INVX1 U357 ( .A(n205), .Y(n206) );
  AND2X2 U359 ( .A(\mem<21><0> ), .B(n539), .Y(n208) );
  INVX1 U361 ( .A(n208), .Y(n209) );
  AND2X2 U363 ( .A(\mem<22><3> ), .B(n541), .Y(n210) );
  INVX1 U364 ( .A(n210), .Y(n211) );
  AND2X2 U365 ( .A(\mem<22><2> ), .B(n541), .Y(n212) );
  INVX1 U368 ( .A(n212), .Y(n213) );
  AND2X2 U370 ( .A(\mem<22><1> ), .B(n541), .Y(n214) );
  INVX1 U372 ( .A(n214), .Y(n215) );
  AND2X2 U377 ( .A(\mem<22><0> ), .B(n541), .Y(n216) );
  INVX1 U378 ( .A(n216), .Y(n217) );
  INVX1 U381 ( .A(n218), .Y(n219) );
  AND2X2 U383 ( .A(\mem<23><2> ), .B(n543), .Y(n220) );
  INVX1 U385 ( .A(n220), .Y(n221) );
  AND2X2 U389 ( .A(\mem<23><1> ), .B(n543), .Y(n222) );
  INVX1 U390 ( .A(n222), .Y(n223) );
  AND2X2 U391 ( .A(\mem<23><0> ), .B(n543), .Y(n224) );
  INVX1 U394 ( .A(n224), .Y(n225) );
  AND2X2 U396 ( .A(\mem<24><4> ), .B(n545), .Y(n226) );
  INVX1 U398 ( .A(n226), .Y(n227) );
  AND2X2 U400 ( .A(\mem<24><3> ), .B(n545), .Y(n228) );
  INVX1 U402 ( .A(n228), .Y(n230) );
  AND2X2 U403 ( .A(\mem<24><1> ), .B(n545), .Y(n231) );
  INVX1 U404 ( .A(n231), .Y(n232) );
  AND2X2 U409 ( .A(\mem<24><0> ), .B(n545), .Y(n233) );
  INVX1 U411 ( .A(n233), .Y(n234) );
  INVX1 U413 ( .A(n237), .Y(n238) );
  AND2X2 U415 ( .A(\mem<25><2> ), .B(n547), .Y(n239) );
  INVX1 U416 ( .A(n239), .Y(n240) );
  AND2X2 U417 ( .A(\mem<25><1> ), .B(n547), .Y(n241) );
  INVX1 U422 ( .A(n241), .Y(n242) );
  AND2X2 U424 ( .A(\mem<25><0> ), .B(n547), .Y(n243) );
  INVX1 U428 ( .A(n243), .Y(n244) );
  AND2X2 U429 ( .A(\mem<26><4> ), .B(n549), .Y(n245) );
  INVX1 U430 ( .A(n245), .Y(n246) );
  AND2X2 U433 ( .A(\mem<26><3> ), .B(n549), .Y(n247) );
  INVX1 U434 ( .A(n247), .Y(n248) );
  AND2X2 U436 ( .A(\mem<26><1> ), .B(n549), .Y(n251) );
  INVX1 U437 ( .A(n251), .Y(n252) );
  AND2X2 U439 ( .A(\mem<26><0> ), .B(n549), .Y(n253) );
  INVX1 U440 ( .A(n253), .Y(n254) );
  INVX1 U442 ( .A(n255), .Y(n257) );
  INVX1 U443 ( .A(n258), .Y(n259) );
  AND2X2 U445 ( .A(\mem<27><2> ), .B(n551), .Y(n260) );
  INVX1 U446 ( .A(n260), .Y(n261) );
  AND2X2 U447 ( .A(\mem<27><1> ), .B(n551), .Y(n262) );
  INVX1 U451 ( .A(n262), .Y(n263) );
  AND2X2 U452 ( .A(\mem<27><0> ), .B(n551), .Y(n264) );
  INVX1 U453 ( .A(n264), .Y(n265) );
  AND2X2 U454 ( .A(\mem<28><3> ), .B(n553), .Y(n267) );
  INVX1 U455 ( .A(n267), .Y(n268) );
  AND2X2 U456 ( .A(\mem<28><2> ), .B(n553), .Y(n269) );
  INVX1 U457 ( .A(n269), .Y(n270) );
  AND2X2 U458 ( .A(\mem<28><1> ), .B(n553), .Y(n271) );
  INVX1 U459 ( .A(n271), .Y(n272) );
  INVX1 U460 ( .A(n274), .Y(n275) );
  AND2X2 U461 ( .A(\mem<29><3> ), .B(n555), .Y(n276) );
  INVX1 U462 ( .A(n276), .Y(n278) );
  AND2X2 U463 ( .A(\mem<29><2> ), .B(n555), .Y(n279) );
  INVX1 U464 ( .A(n279), .Y(n280) );
  INVX1 U465 ( .A(n281), .Y(n282) );
  AND2X2 U466 ( .A(\mem<29><0> ), .B(n555), .Y(n283) );
  INVX1 U467 ( .A(n283), .Y(n284) );
  INVX1 U468 ( .A(n285), .Y(n287) );
  AND2X2 U469 ( .A(\mem<30><3> ), .B(n557), .Y(n448) );
  INVX1 U470 ( .A(n448), .Y(n449) );
  AND2X2 U471 ( .A(\mem<30><2> ), .B(n557), .Y(n450) );
  INVX1 U472 ( .A(n450), .Y(n451) );
  AND2X2 U473 ( .A(\mem<30><1> ), .B(n557), .Y(n452) );
  INVX1 U474 ( .A(n452), .Y(n453) );
  AND2X2 U475 ( .A(\mem<30><0> ), .B(n557), .Y(n454) );
  INVX1 U476 ( .A(n454), .Y(n455) );
  AND2X2 U477 ( .A(\mem<31><3> ), .B(n559), .Y(n456) );
  INVX1 U478 ( .A(n456), .Y(n457) );
  AND2X2 U479 ( .A(\mem<31><2> ), .B(n559), .Y(n458) );
  INVX1 U480 ( .A(n458), .Y(n459) );
  INVX1 U481 ( .A(n460), .Y(n461) );
  INVX1 U482 ( .A(n462), .Y(n463) );
  OR2X1 U483 ( .A(n777), .B(n808), .Y(n471) );
  INVX8 U484 ( .A(n634), .Y(n636) );
  MUX2X1 U485 ( .B(n788), .A(n789), .S(n464), .Y(n790) );
  MUX2X1 U486 ( .B(n675), .A(n674), .S(N11), .Y(n679) );
  INVX4 U487 ( .A(n638), .Y(n624) );
  MUX2X1 U488 ( .B(n680), .A(n681), .S(n650), .Y(n682) );
  INVX4 U489 ( .A(n627), .Y(n633) );
  INVX8 U490 ( .A(n645), .Y(n641) );
  OR2X1 U491 ( .A(n684), .B(n808), .Y(n465) );
  MUX2X1 U492 ( .B(n666), .A(n667), .S(n650), .Y(n683) );
  INVX8 U493 ( .A(n650), .Y(n649) );
  MUX2X1 U494 ( .B(n672), .A(n673), .S(n4), .Y(n681) );
  MUX2X1 U495 ( .B(n698), .A(n697), .S(N13), .Y(n714) );
  INVX8 U496 ( .A(N13), .Y(n650) );
  INVX1 U497 ( .A(n465), .Y(\data_out<0> ) );
  INVX1 U498 ( .A(n471), .Y(\data_out<3> ) );
  INVX1 U499 ( .A(n473), .Y(\data_out<4> ) );
  AND2X2 U500 ( .A(\mem<0><1> ), .B(n497), .Y(n475) );
  INVX1 U501 ( .A(n475), .Y(n476) );
  AND2X2 U502 ( .A(\mem<2><1> ), .B(n501), .Y(n477) );
  INVX1 U503 ( .A(n477), .Y(n478) );
  AND2X2 U504 ( .A(\mem<10><1> ), .B(n517), .Y(n479) );
  INVX1 U505 ( .A(n479), .Y(n480) );
  AND2X2 U506 ( .A(\mem<18><2> ), .B(n533), .Y(n481) );
  INVX1 U507 ( .A(n481), .Y(n482) );
  AND2X2 U508 ( .A(\mem<24><2> ), .B(n545), .Y(n483) );
  INVX1 U509 ( .A(n483), .Y(n484) );
  AND2X2 U510 ( .A(\mem<26><2> ), .B(n549), .Y(n485) );
  INVX1 U511 ( .A(n485), .Y(n486) );
  AND2X1 U512 ( .A(\data_in<4> ), .B(n1010), .Y(n487) );
  AND2X1 U513 ( .A(\data_in<3> ), .B(n1010), .Y(n488) );
  AND2X1 U514 ( .A(\data_in<2> ), .B(n1010), .Y(n489) );
  AND2X1 U515 ( .A(\data_in<1> ), .B(n1010), .Y(n490) );
  AND2X1 U516 ( .A(\data_in<0> ), .B(n1010), .Y(n491) );
  BUFX2 U517 ( .A(n974), .Y(n492) );
  INVX1 U518 ( .A(n492), .Y(n810) );
  BUFX2 U519 ( .A(n983), .Y(n493) );
  INVX1 U520 ( .A(n493), .Y(n813) );
  BUFX2 U521 ( .A(n989), .Y(n494) );
  INVX1 U522 ( .A(n494), .Y(n811) );
  BUFX2 U523 ( .A(n998), .Y(n495) );
  INVX1 U524 ( .A(n495), .Y(n812) );
  INVX1 U525 ( .A(n487), .Y(n628) );
  INVX1 U526 ( .A(n488), .Y(n629) );
  INVX1 U527 ( .A(n489), .Y(n630) );
  INVX1 U528 ( .A(n490), .Y(n631) );
  INVX1 U529 ( .A(n491), .Y(n632) );
  AND2X1 U530 ( .A(n562), .B(n1010), .Y(n496) );
  INVX1 U531 ( .A(n496), .Y(n497) );
  AND2X1 U532 ( .A(n564), .B(n1010), .Y(n498) );
  INVX1 U533 ( .A(n498), .Y(n499) );
  AND2X1 U534 ( .A(n567), .B(n1010), .Y(n500) );
  INVX1 U535 ( .A(n500), .Y(n501) );
  AND2X1 U536 ( .A(n569), .B(n1010), .Y(n502) );
  INVX1 U537 ( .A(n502), .Y(n503) );
  AND2X1 U538 ( .A(n571), .B(n1010), .Y(n504) );
  INVX1 U539 ( .A(n504), .Y(n505) );
  AND2X1 U540 ( .A(n572), .B(n1010), .Y(n506) );
  INVX1 U541 ( .A(n506), .Y(n507) );
  AND2X1 U542 ( .A(n574), .B(n1010), .Y(n508) );
  INVX1 U543 ( .A(n508), .Y(n509) );
  AND2X1 U544 ( .A(n576), .B(n1010), .Y(n510) );
  INVX1 U545 ( .A(n510), .Y(n511) );
  AND2X1 U546 ( .A(n578), .B(n1010), .Y(n512) );
  INVX1 U547 ( .A(n512), .Y(n513) );
  AND2X1 U548 ( .A(n580), .B(n1010), .Y(n514) );
  INVX1 U549 ( .A(n514), .Y(n515) );
  AND2X1 U550 ( .A(n583), .B(n1010), .Y(n516) );
  INVX1 U551 ( .A(n516), .Y(n517) );
  AND2X1 U552 ( .A(n585), .B(n1010), .Y(n518) );
  INVX1 U553 ( .A(n518), .Y(n519) );
  AND2X1 U554 ( .A(n587), .B(n1010), .Y(n520) );
  INVX1 U555 ( .A(n520), .Y(n521) );
  AND2X1 U556 ( .A(n588), .B(n1010), .Y(n522) );
  INVX1 U557 ( .A(n522), .Y(n523) );
  AND2X1 U558 ( .A(n590), .B(n1010), .Y(n524) );
  INVX1 U559 ( .A(n524), .Y(n525) );
  AND2X1 U560 ( .A(n592), .B(n1010), .Y(n526) );
  INVX1 U561 ( .A(n526), .Y(n527) );
  AND2X1 U562 ( .A(n594), .B(n1010), .Y(n528) );
  INVX1 U563 ( .A(n528), .Y(n529) );
  AND2X1 U564 ( .A(n596), .B(n1010), .Y(n530) );
  INVX1 U565 ( .A(n530), .Y(n531) );
  AND2X1 U566 ( .A(n599), .B(n1010), .Y(n532) );
  INVX1 U567 ( .A(n532), .Y(n533) );
  AND2X1 U568 ( .A(n600), .B(n1010), .Y(n534) );
  INVX1 U569 ( .A(n534), .Y(n535) );
  AND2X1 U570 ( .A(n602), .B(n1010), .Y(n536) );
  INVX1 U571 ( .A(n536), .Y(n537) );
  AND2X1 U572 ( .A(n604), .B(n1010), .Y(n538) );
  INVX1 U573 ( .A(n538), .Y(n539) );
  AND2X1 U574 ( .A(n606), .B(n1010), .Y(n540) );
  INVX1 U575 ( .A(n540), .Y(n541) );
  AND2X1 U576 ( .A(n608), .B(n1010), .Y(n542) );
  INVX1 U577 ( .A(n542), .Y(n543) );
  AND2X1 U578 ( .A(n610), .B(n1010), .Y(n544) );
  INVX1 U579 ( .A(n544), .Y(n545) );
  AND2X1 U580 ( .A(n612), .B(n1010), .Y(n546) );
  INVX1 U581 ( .A(n546), .Y(n547) );
  AND2X1 U582 ( .A(n614), .B(n1010), .Y(n548) );
  INVX1 U583 ( .A(n548), .Y(n549) );
  AND2X1 U584 ( .A(n616), .B(n1010), .Y(n550) );
  INVX1 U585 ( .A(n550), .Y(n551) );
  AND2X1 U586 ( .A(n618), .B(n1010), .Y(n552) );
  INVX1 U587 ( .A(n552), .Y(n553) );
  AND2X1 U588 ( .A(n620), .B(n1010), .Y(n554) );
  INVX1 U589 ( .A(n554), .Y(n555) );
  AND2X1 U590 ( .A(n622), .B(n1010), .Y(n556) );
  INVX1 U591 ( .A(n556), .Y(n557) );
  AND2X1 U592 ( .A(n560), .B(n1010), .Y(n558) );
  INVX1 U593 ( .A(n558), .Y(n559) );
  AND2X1 U594 ( .A(n1009), .B(n812), .Y(n560) );
  INVX1 U595 ( .A(n560), .Y(n561) );
  AND2X1 U596 ( .A(n810), .B(n999), .Y(n562) );
  INVX1 U597 ( .A(n562), .Y(n563) );
  AND2X1 U598 ( .A(n810), .B(n1000), .Y(n564) );
  INVX1 U599 ( .A(n564), .Y(n565) );
  INVX1 U600 ( .A(n567), .Y(n566) );
  AND2X1 U601 ( .A(n810), .B(n1002), .Y(n567) );
  INVX1 U602 ( .A(n569), .Y(n568) );
  AND2X1 U603 ( .A(n810), .B(n1003), .Y(n569) );
  INVX1 U604 ( .A(n571), .Y(n570) );
  AND2X1 U605 ( .A(n810), .B(n1004), .Y(n571) );
  AND2X1 U606 ( .A(n810), .B(n1006), .Y(n572) );
  INVX1 U607 ( .A(n572), .Y(n573) );
  AND2X1 U608 ( .A(n810), .B(n1008), .Y(n574) );
  INVX1 U609 ( .A(n574), .Y(n575) );
  AND2X1 U610 ( .A(n810), .B(n1009), .Y(n576) );
  INVX1 U611 ( .A(n576), .Y(n577) );
  AND2X1 U612 ( .A(n813), .B(n999), .Y(n578) );
  INVX1 U613 ( .A(n578), .Y(n579) );
  AND2X1 U614 ( .A(n813), .B(n1000), .Y(n580) );
  INVX1 U615 ( .A(n580), .Y(n581) );
  INVX1 U616 ( .A(n583), .Y(n582) );
  AND2X1 U617 ( .A(n813), .B(n1002), .Y(n583) );
  INVX1 U618 ( .A(n585), .Y(n584) );
  AND2X1 U619 ( .A(n813), .B(n1003), .Y(n585) );
  INVX1 U620 ( .A(n587), .Y(n586) );
  AND2X1 U621 ( .A(n813), .B(n1004), .Y(n587) );
  AND2X1 U622 ( .A(n813), .B(n1006), .Y(n588) );
  INVX1 U623 ( .A(n588), .Y(n589) );
  AND2X1 U624 ( .A(n813), .B(n1008), .Y(n590) );
  INVX1 U625 ( .A(n590), .Y(n591) );
  AND2X1 U626 ( .A(n813), .B(n1009), .Y(n592) );
  INVX1 U627 ( .A(n592), .Y(n593) );
  AND2X1 U628 ( .A(n811), .B(n999), .Y(n594) );
  INVX1 U629 ( .A(n594), .Y(n595) );
  AND2X1 U630 ( .A(n811), .B(n1000), .Y(n596) );
  INVX1 U631 ( .A(n596), .Y(n597) );
  INVX1 U632 ( .A(n599), .Y(n598) );
  AND2X1 U633 ( .A(n811), .B(n1002), .Y(n599) );
  AND2X1 U634 ( .A(n811), .B(n1003), .Y(n600) );
  INVX1 U635 ( .A(n600), .Y(n601) );
  AND2X1 U636 ( .A(n811), .B(n1004), .Y(n602) );
  INVX1 U637 ( .A(n602), .Y(n603) );
  AND2X1 U638 ( .A(n811), .B(n1006), .Y(n604) );
  INVX1 U639 ( .A(n604), .Y(n605) );
  AND2X1 U640 ( .A(n811), .B(n1008), .Y(n606) );
  INVX1 U641 ( .A(n606), .Y(n607) );
  AND2X1 U642 ( .A(n811), .B(n1009), .Y(n608) );
  INVX1 U643 ( .A(n608), .Y(n609) );
  AND2X1 U644 ( .A(n999), .B(n812), .Y(n610) );
  INVX1 U645 ( .A(n610), .Y(n611) );
  AND2X1 U646 ( .A(n1000), .B(n812), .Y(n612) );
  INVX1 U647 ( .A(n612), .Y(n613) );
  AND2X1 U648 ( .A(n1002), .B(n812), .Y(n614) );
  INVX1 U649 ( .A(n614), .Y(n615) );
  AND2X1 U650 ( .A(n1003), .B(n812), .Y(n616) );
  INVX1 U651 ( .A(n616), .Y(n617) );
  AND2X1 U652 ( .A(n1004), .B(n812), .Y(n618) );
  INVX1 U653 ( .A(n618), .Y(n619) );
  AND2X1 U654 ( .A(n1006), .B(n812), .Y(n620) );
  INVX1 U655 ( .A(n620), .Y(n621) );
  AND2X1 U656 ( .A(n1008), .B(n812), .Y(n622) );
  INVX1 U657 ( .A(n622), .Y(n623) );
  MUX2X1 U658 ( .B(n744), .A(n745), .S(n652), .Y(n746) );
  MUX2X1 U659 ( .B(n676), .A(n677), .S(n645), .Y(n678) );
  MUX2X1 U660 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2), .Y(n702) );
  MUX2X1 U661 ( .B(\mem<7><1> ), .A(\mem<6><1> ), .S(n634), .Y(n687) );
  MUX2X1 U662 ( .B(n784), .A(n785), .S(n646), .Y(n789) );
  INVX4 U663 ( .A(N10), .Y(n634) );
  INVX1 U664 ( .A(n638), .Y(n625) );
  INVX8 U665 ( .A(N10), .Y(n627) );
  INVX1 U666 ( .A(n637), .Y(n640) );
  MUX2X1 U667 ( .B(n771), .A(n772), .S(n5), .Y(n773) );
  INVX1 U668 ( .A(n2), .Y(n639) );
  MUX2X1 U669 ( .B(\mem<3><0> ), .A(\mem<2><0> ), .S(n624), .Y(n654) );
  MUX2X1 U670 ( .B(n682), .A(n683), .S(n652), .Y(n684) );
  MUX2X1 U671 ( .B(\mem<11><0> ), .A(\mem<10><0> ), .S(n624), .Y(n660) );
  MUX2X1 U672 ( .B(\mem<29><0> ), .A(\mem<28><0> ), .S(n625), .Y(n677) );
  MUX2X1 U673 ( .B(n658), .A(n659), .S(n648), .Y(n667) );
  MUX2X1 U674 ( .B(n775), .A(n776), .S(n652), .Y(n777) );
  MUX2X1 U675 ( .B(\mem<21><2> ), .A(\mem<20><2> ), .S(n626), .Y(n733) );
  MUX2X1 U676 ( .B(n774), .A(n773), .S(N13), .Y(n775) );
  INVX8 U677 ( .A(n627), .Y(n635) );
  INVX8 U678 ( .A(n634), .Y(n637) );
  INVX8 U679 ( .A(n627), .Y(n638) );
  INVX8 U680 ( .A(n645), .Y(n642) );
  INVX8 U681 ( .A(n646), .Y(n643) );
  INVX8 U682 ( .A(n645), .Y(n644) );
  INVX8 U683 ( .A(N11), .Y(n645) );
  INVX8 U684 ( .A(N11), .Y(n646) );
  INVX8 U685 ( .A(n648), .Y(n647) );
  INVX8 U686 ( .A(N12), .Y(n648) );
  INVX8 U687 ( .A(N14), .Y(n652) );
  OR2X2 U688 ( .A(write), .B(rst), .Y(n808) );
  MUX2X1 U689 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n637), .Y(n655) );
  MUX2X1 U690 ( .B(n655), .A(n654), .S(n641), .Y(n659) );
  MUX2X1 U691 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n637), .Y(n657) );
  MUX2X1 U692 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n636), .Y(n656) );
  MUX2X1 U693 ( .B(n657), .A(n656), .S(n641), .Y(n658) );
  MUX2X1 U694 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n637), .Y(n661) );
  MUX2X1 U695 ( .B(n661), .A(n660), .S(n641), .Y(n665) );
  MUX2X1 U696 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n635), .Y(n663) );
  MUX2X1 U697 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n636), .Y(n662) );
  MUX2X1 U698 ( .B(n663), .A(n662), .S(n641), .Y(n664) );
  MUX2X1 U699 ( .B(n665), .A(n664), .S(N12), .Y(n666) );
  MUX2X1 U700 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n2), .Y(n669) );
  MUX2X1 U701 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n635), .Y(n668) );
  MUX2X1 U702 ( .B(n669), .A(n668), .S(n641), .Y(n673) );
  MUX2X1 U703 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n2), .Y(n671) );
  MUX2X1 U704 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n638), .Y(n670) );
  MUX2X1 U705 ( .B(n671), .A(n670), .S(n641), .Y(n672) );
  MUX2X1 U706 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n636), .Y(n675) );
  MUX2X1 U707 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n635), .Y(n674) );
  MUX2X1 U708 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n636), .Y(n676) );
  MUX2X1 U709 ( .B(n679), .A(n678), .S(N12), .Y(n680) );
  MUX2X1 U710 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n636), .Y(n686) );
  MUX2X1 U711 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n633), .Y(n685) );
  MUX2X1 U712 ( .B(n688), .A(n687), .S(n641), .Y(n689) );
  MUX2X1 U713 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2), .Y(n692) );
  MUX2X1 U714 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n635), .Y(n691) );
  MUX2X1 U715 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n638), .Y(n694) );
  MUX2X1 U716 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n638), .Y(n693) );
  MUX2X1 U717 ( .B(n694), .A(n693), .S(n641), .Y(n695) );
  MUX2X1 U718 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n635), .Y(n700) );
  MUX2X1 U719 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n637), .Y(n699) );
  MUX2X1 U720 ( .B(n700), .A(n699), .S(n642), .Y(n704) );
  MUX2X1 U721 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n635), .Y(n701) );
  MUX2X1 U722 ( .B(n702), .A(n701), .S(n642), .Y(n703) );
  MUX2X1 U723 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n2), .Y(n706) );
  MUX2X1 U724 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n635), .Y(n705) );
  MUX2X1 U725 ( .B(n706), .A(n705), .S(n642), .Y(n710) );
  MUX2X1 U726 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n636), .Y(n708) );
  MUX2X1 U727 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n636), .Y(n707) );
  MUX2X1 U728 ( .B(n708), .A(n707), .S(n642), .Y(n709) );
  MUX2X1 U729 ( .B(n710), .A(n709), .S(N12), .Y(n711) );
  MUX2X1 U730 ( .B(n712), .A(n711), .S(n649), .Y(n713) );
  MUX2X1 U731 ( .B(n714), .A(n713), .S(n651), .Y(n715) );
  MUX2X1 U732 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2), .Y(n717) );
  MUX2X1 U733 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n633), .Y(n716) );
  MUX2X1 U734 ( .B(n717), .A(n716), .S(n642), .Y(n721) );
  MUX2X1 U735 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n633), .Y(n719) );
  MUX2X1 U736 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n637), .Y(n718) );
  MUX2X1 U737 ( .B(n719), .A(n718), .S(n642), .Y(n720) );
  MUX2X1 U738 ( .B(n721), .A(n720), .S(N12), .Y(n729) );
  MUX2X1 U739 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n637), .Y(n723) );
  MUX2X1 U740 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n635), .Y(n722) );
  MUX2X1 U741 ( .B(n723), .A(n722), .S(n642), .Y(n727) );
  MUX2X1 U742 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n637), .Y(n725) );
  MUX2X1 U743 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2), .Y(n724) );
  MUX2X1 U744 ( .B(n725), .A(n724), .S(n642), .Y(n726) );
  MUX2X1 U745 ( .B(n727), .A(n726), .S(N12), .Y(n728) );
  MUX2X1 U746 ( .B(n729), .A(n728), .S(n649), .Y(n745) );
  MUX2X1 U747 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n638), .Y(n731) );
  MUX2X1 U748 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n638), .Y(n730) );
  MUX2X1 U749 ( .B(n731), .A(n730), .S(n642), .Y(n735) );
  MUX2X1 U750 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2), .Y(n732) );
  MUX2X1 U751 ( .B(n733), .A(n732), .S(n642), .Y(n734) );
  MUX2X1 U752 ( .B(n735), .A(n734), .S(N12), .Y(n743) );
  MUX2X1 U753 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n638), .Y(n737) );
  MUX2X1 U754 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n638), .Y(n736) );
  MUX2X1 U755 ( .B(n737), .A(n736), .S(n642), .Y(n741) );
  MUX2X1 U756 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n2), .Y(n739) );
  MUX2X1 U757 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2), .Y(n738) );
  MUX2X1 U758 ( .B(n739), .A(n738), .S(n642), .Y(n740) );
  MUX2X1 U759 ( .B(n741), .A(n740), .S(N12), .Y(n742) );
  MUX2X1 U760 ( .B(n743), .A(n742), .S(n649), .Y(n744) );
  MUX2X1 U761 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2), .Y(n748) );
  MUX2X1 U762 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n2), .Y(n747) );
  MUX2X1 U763 ( .B(n748), .A(n747), .S(n643), .Y(n752) );
  MUX2X1 U764 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n635), .Y(n750) );
  MUX2X1 U765 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n637), .Y(n749) );
  MUX2X1 U766 ( .B(n750), .A(n749), .S(n643), .Y(n751) );
  MUX2X1 U767 ( .B(n752), .A(n751), .S(n647), .Y(n760) );
  MUX2X1 U768 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n635), .Y(n754) );
  MUX2X1 U769 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n633), .Y(n753) );
  MUX2X1 U770 ( .B(n754), .A(n753), .S(n643), .Y(n758) );
  MUX2X1 U771 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n636), .Y(n756) );
  MUX2X1 U772 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n2), .Y(n755) );
  MUX2X1 U773 ( .B(n756), .A(n755), .S(n643), .Y(n757) );
  MUX2X1 U774 ( .B(n758), .A(n757), .S(n647), .Y(n759) );
  MUX2X1 U775 ( .B(n760), .A(n759), .S(n649), .Y(n776) );
  MUX2X1 U776 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n633), .Y(n762) );
  MUX2X1 U777 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n635), .Y(n761) );
  MUX2X1 U778 ( .B(n762), .A(n761), .S(n643), .Y(n766) );
  MUX2X1 U779 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n636), .Y(n764) );
  MUX2X1 U780 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n635), .Y(n763) );
  MUX2X1 U781 ( .B(n764), .A(n763), .S(n643), .Y(n765) );
  MUX2X1 U782 ( .B(n766), .A(n765), .S(n647), .Y(n774) );
  MUX2X1 U783 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n636), .Y(n768) );
  MUX2X1 U784 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2), .Y(n767) );
  MUX2X1 U785 ( .B(n768), .A(n767), .S(n643), .Y(n772) );
  MUX2X1 U786 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n635), .Y(n770) );
  MUX2X1 U787 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n633), .Y(n769) );
  MUX2X1 U788 ( .B(n770), .A(n769), .S(n643), .Y(n771) );
  MUX2X1 U789 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n633), .Y(n779) );
  MUX2X1 U790 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n635), .Y(n778) );
  MUX2X1 U791 ( .B(n779), .A(n778), .S(n643), .Y(n783) );
  MUX2X1 U792 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2), .Y(n781) );
  MUX2X1 U793 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n636), .Y(n780) );
  MUX2X1 U794 ( .B(n781), .A(n780), .S(n643), .Y(n782) );
  MUX2X1 U795 ( .B(n783), .A(n782), .S(n647), .Y(n791) );
  MUX2X1 U796 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n636), .Y(n785) );
  MUX2X1 U797 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n637), .Y(n787) );
  MUX2X1 U798 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2), .Y(n786) );
  MUX2X1 U799 ( .B(n787), .A(n786), .S(n643), .Y(n788) );
  MUX2X1 U800 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n637), .Y(n793) );
  MUX2X1 U801 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n635), .Y(n792) );
  MUX2X1 U802 ( .B(n793), .A(n792), .S(n644), .Y(n797) );
  MUX2X1 U803 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2), .Y(n795) );
  MUX2X1 U804 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n636), .Y(n794) );
  MUX2X1 U805 ( .B(n795), .A(n794), .S(n644), .Y(n796) );
  MUX2X1 U806 ( .B(n797), .A(n796), .S(n647), .Y(n805) );
  MUX2X1 U807 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n635), .Y(n799) );
  MUX2X1 U808 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n637), .Y(n798) );
  MUX2X1 U809 ( .B(n799), .A(n798), .S(n644), .Y(n803) );
  MUX2X1 U810 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n635), .Y(n801) );
  MUX2X1 U811 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n633), .Y(n800) );
  MUX2X1 U812 ( .B(n801), .A(n800), .S(n644), .Y(n802) );
  MUX2X1 U813 ( .B(n803), .A(n802), .S(n647), .Y(n804) );
  MUX2X1 U814 ( .B(n805), .A(n804), .S(n649), .Y(n806) );
endmodule


module memc_Size1_0 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n214), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n215), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n216), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n217), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n218), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n219), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n220), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n221), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n222), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n223), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n224), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n225), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n226), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n227), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n228), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n229), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n230), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n231), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n232), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n233), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n234), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n235), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n236), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n238), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n239), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n240), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n241), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n242), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n243), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n244), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n245), .CLK(clk), .Q(\mem<31><0> ) );
  INVX2 U2 ( .A(n9), .Y(n7) );
  INVX1 U3 ( .A(rst), .Y(n168) );
  INVX1 U4 ( .A(n153), .Y(N17) );
  INVX1 U5 ( .A(n161), .Y(n154) );
  INVX1 U6 ( .A(N12), .Y(n163) );
  INVX1 U7 ( .A(n107), .Y(n198) );
  INVX1 U8 ( .A(n108), .Y(n201) );
  INVX1 U9 ( .A(n109), .Y(n204) );
  INVX1 U10 ( .A(n110), .Y(n207) );
  INVX1 U11 ( .A(n111), .Y(n210) );
  INVX2 U12 ( .A(n159), .Y(n155) );
  AND2X1 U13 ( .A(n159), .B(n98), .Y(n115) );
  INVX1 U14 ( .A(n167), .Y(n166) );
  INVX1 U15 ( .A(n11), .Y(n1) );
  BUFX2 U16 ( .A(write), .Y(n2) );
  INVX1 U17 ( .A(n120), .Y(n3) );
  INVX1 U18 ( .A(n8), .Y(n4) );
  INVX1 U19 ( .A(n1), .Y(n5) );
  INVX1 U20 ( .A(n1), .Y(n6) );
  AND2X2 U21 ( .A(\data_in<0> ), .B(n156), .Y(n118) );
  AND2X2 U22 ( .A(\data_in<0> ), .B(n1), .Y(n104) );
  AND2X2 U23 ( .A(\data_in<0> ), .B(n4), .Y(n103) );
  OR2X2 U24 ( .A(n101), .B(n2), .Y(n95) );
  OR2X2 U25 ( .A(n165), .B(n10), .Y(n8) );
  INVX1 U26 ( .A(n8), .Y(n9) );
  OR2X2 U27 ( .A(n121), .B(n12), .Y(n10) );
  OR2X2 U28 ( .A(n122), .B(n10), .Y(n11) );
  OR2X2 U29 ( .A(\addr<5> ), .B(n93), .Y(n12) );
  INVX1 U30 ( .A(n12), .Y(n13) );
  AND2X2 U31 ( .A(n94), .B(n117), .Y(n14) );
  INVX1 U32 ( .A(n14), .Y(n15) );
  AND2X2 U33 ( .A(n113), .B(n94), .Y(n16) );
  INVX1 U34 ( .A(n16), .Y(n17) );
  AND2X2 U35 ( .A(n198), .B(n94), .Y(n18) );
  INVX1 U36 ( .A(n18), .Y(n19) );
  AND2X2 U37 ( .A(n201), .B(n94), .Y(n20) );
  INVX1 U38 ( .A(n20), .Y(n21) );
  AND2X2 U39 ( .A(n204), .B(n94), .Y(n22) );
  INVX1 U40 ( .A(n22), .Y(n23) );
  AND2X2 U41 ( .A(n207), .B(n94), .Y(n24) );
  INVX1 U42 ( .A(n24), .Y(n25) );
  AND2X2 U43 ( .A(n210), .B(n94), .Y(n26) );
  INVX1 U44 ( .A(n26), .Y(n27) );
  AND2X2 U45 ( .A(n115), .B(n94), .Y(n28) );
  INVX1 U46 ( .A(n28), .Y(n29) );
  AND2X2 U47 ( .A(n117), .B(n103), .Y(n30) );
  AND2X2 U48 ( .A(n113), .B(n103), .Y(n31) );
  INVX1 U49 ( .A(n31), .Y(n32) );
  AND2X2 U50 ( .A(n198), .B(n103), .Y(n33) );
  INVX1 U51 ( .A(n33), .Y(n34) );
  AND2X2 U52 ( .A(n201), .B(n103), .Y(n35) );
  INVX1 U53 ( .A(n35), .Y(n36) );
  AND2X2 U54 ( .A(n204), .B(n103), .Y(n37) );
  INVX1 U55 ( .A(n37), .Y(n38) );
  AND2X2 U56 ( .A(n207), .B(n103), .Y(n39) );
  INVX1 U57 ( .A(n39), .Y(n40) );
  AND2X2 U58 ( .A(n210), .B(n103), .Y(n41) );
  INVX1 U59 ( .A(n41), .Y(n42) );
  AND2X2 U60 ( .A(n115), .B(n103), .Y(n43) );
  INVX1 U61 ( .A(n43), .Y(n44) );
  AND2X2 U62 ( .A(n117), .B(n104), .Y(n45) );
  INVX1 U63 ( .A(n45), .Y(n46) );
  AND2X2 U64 ( .A(n113), .B(n104), .Y(n47) );
  INVX1 U65 ( .A(n47), .Y(n48) );
  AND2X2 U66 ( .A(n198), .B(n104), .Y(n49) );
  INVX1 U67 ( .A(n49), .Y(n50) );
  AND2X2 U68 ( .A(n201), .B(n104), .Y(n51) );
  INVX1 U69 ( .A(n51), .Y(n52) );
  AND2X2 U70 ( .A(n204), .B(n104), .Y(n53) );
  INVX1 U71 ( .A(n53), .Y(n54) );
  AND2X2 U72 ( .A(n207), .B(n104), .Y(n55) );
  INVX1 U73 ( .A(n55), .Y(n56) );
  AND2X2 U74 ( .A(n210), .B(n104), .Y(n57) );
  INVX1 U75 ( .A(n57), .Y(n58) );
  AND2X2 U76 ( .A(n115), .B(n104), .Y(n59) );
  INVX1 U77 ( .A(n59), .Y(n60) );
  BUFX2 U78 ( .A(n169), .Y(n93) );
  AND2X2 U79 ( .A(\data_in<0> ), .B(n120), .Y(n94) );
  INVX1 U80 ( .A(n163), .Y(n162) );
  INVX1 U81 ( .A(n161), .Y(n160) );
  INVX1 U82 ( .A(n159), .Y(n158) );
  INVX1 U83 ( .A(n95), .Y(\data_out<0> ) );
  OR2X1 U84 ( .A(n160), .B(n162), .Y(n97) );
  INVX1 U85 ( .A(n97), .Y(n98) );
  INVX1 U86 ( .A(n30), .Y(n99) );
  AND2X1 U87 ( .A(N17), .B(n168), .Y(n100) );
  INVX1 U88 ( .A(n100), .Y(n101) );
  AND2X1 U89 ( .A(n162), .B(n160), .Y(n102) );
  OR2X1 U90 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n105) );
  INVX1 U91 ( .A(n105), .Y(n106) );
  BUFX2 U92 ( .A(n199), .Y(n107) );
  BUFX2 U93 ( .A(n202), .Y(n108) );
  BUFX2 U94 ( .A(n205), .Y(n109) );
  BUFX2 U95 ( .A(n208), .Y(n110) );
  BUFX2 U96 ( .A(n211), .Y(n111) );
  INVX1 U97 ( .A(n113), .Y(n112) );
  AND2X1 U98 ( .A(n159), .B(n102), .Y(n113) );
  INVX1 U99 ( .A(n115), .Y(n114) );
  INVX1 U100 ( .A(n117), .Y(n116) );
  AND2X1 U101 ( .A(n158), .B(n102), .Y(n117) );
  INVX1 U102 ( .A(n118), .Y(n119) );
  INVX1 U103 ( .A(n186), .Y(n120) );
  INVX1 U104 ( .A(n167), .Y(n121) );
  INVX1 U105 ( .A(n165), .Y(n122) );
  INVX1 U106 ( .A(N13), .Y(n165) );
  INVX1 U107 ( .A(N14), .Y(n167) );
  MUX2X1 U108 ( .B(n124), .A(n125), .S(n154), .Y(n123) );
  MUX2X1 U109 ( .B(n127), .A(n128), .S(n154), .Y(n126) );
  MUX2X1 U110 ( .B(n130), .A(n131), .S(n154), .Y(n129) );
  MUX2X1 U111 ( .B(n133), .A(n134), .S(n154), .Y(n132) );
  MUX2X1 U112 ( .B(n136), .A(n137), .S(n164), .Y(n135) );
  MUX2X1 U113 ( .B(n139), .A(n140), .S(n154), .Y(n138) );
  MUX2X1 U114 ( .B(n142), .A(n143), .S(n154), .Y(n141) );
  MUX2X1 U115 ( .B(n145), .A(n146), .S(n154), .Y(n144) );
  MUX2X1 U116 ( .B(n148), .A(n149), .S(n154), .Y(n147) );
  MUX2X1 U117 ( .B(n151), .A(n152), .S(n164), .Y(n150) );
  MUX2X1 U118 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n155), .Y(n125) );
  MUX2X1 U119 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n155), .Y(n124) );
  MUX2X1 U120 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n155), .Y(n128) );
  MUX2X1 U121 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n155), .Y(n127) );
  MUX2X1 U122 ( .B(n126), .A(n123), .S(n162), .Y(n137) );
  MUX2X1 U123 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n155), .Y(n131) );
  MUX2X1 U124 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n155), .Y(n130) );
  MUX2X1 U125 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n155), .Y(n134) );
  MUX2X1 U126 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n155), .Y(n133) );
  MUX2X1 U127 ( .B(n132), .A(n129), .S(n162), .Y(n136) );
  MUX2X1 U128 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n155), .Y(n140) );
  MUX2X1 U129 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n155), .Y(n139) );
  MUX2X1 U130 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n155), .Y(n143) );
  MUX2X1 U131 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n155), .Y(n142) );
  MUX2X1 U132 ( .B(n141), .A(n138), .S(n162), .Y(n152) );
  MUX2X1 U133 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n155), .Y(n146) );
  MUX2X1 U134 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n155), .Y(n145) );
  MUX2X1 U135 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n155), .Y(n149) );
  MUX2X1 U136 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n155), .Y(n148) );
  MUX2X1 U137 ( .B(n147), .A(n144), .S(n162), .Y(n151) );
  MUX2X1 U138 ( .B(n150), .A(n135), .S(n166), .Y(n153) );
  INVX1 U139 ( .A(N11), .Y(n161) );
  INVX1 U140 ( .A(n13), .Y(n157) );
  INVX1 U141 ( .A(N10), .Y(n159) );
  NOR3X1 U142 ( .A(n167), .B(n165), .C(n157), .Y(n156) );
  INVX2 U143 ( .A(n156), .Y(n177) );
  INVX1 U144 ( .A(n165), .Y(n164) );
  NAND3X1 U145 ( .A(n168), .B(n106), .C(write), .Y(n169) );
  OAI21X1 U146 ( .A(n177), .B(n116), .C(\mem<31><0> ), .Y(n170) );
  OAI21X1 U147 ( .A(n119), .B(n116), .C(n170), .Y(n245) );
  OAI21X1 U148 ( .A(n112), .B(n177), .C(\mem<30><0> ), .Y(n171) );
  OAI21X1 U149 ( .A(n112), .B(n119), .C(n171), .Y(n244) );
  NAND3X1 U150 ( .A(n158), .B(n162), .C(n161), .Y(n199) );
  OAI21X1 U151 ( .A(n107), .B(n177), .C(\mem<29><0> ), .Y(n172) );
  OAI21X1 U152 ( .A(n107), .B(n119), .C(n172), .Y(n243) );
  NAND3X1 U153 ( .A(n162), .B(n161), .C(n159), .Y(n202) );
  OAI21X1 U154 ( .A(n108), .B(n177), .C(\mem<28><0> ), .Y(n173) );
  OAI21X1 U155 ( .A(n108), .B(n119), .C(n173), .Y(n242) );
  NAND3X1 U156 ( .A(n158), .B(n160), .C(n163), .Y(n205) );
  OAI21X1 U157 ( .A(n109), .B(n177), .C(\mem<27><0> ), .Y(n174) );
  OAI21X1 U158 ( .A(n109), .B(n119), .C(n174), .Y(n241) );
  NAND3X1 U159 ( .A(n163), .B(n160), .C(n159), .Y(n208) );
  OAI21X1 U160 ( .A(n110), .B(n177), .C(\mem<26><0> ), .Y(n175) );
  OAI21X1 U161 ( .A(n110), .B(n119), .C(n175), .Y(n240) );
  NAND3X1 U162 ( .A(n158), .B(n163), .C(n161), .Y(n211) );
  OAI21X1 U163 ( .A(n111), .B(n177), .C(\mem<25><0> ), .Y(n176) );
  OAI21X1 U164 ( .A(n111), .B(n119), .C(n176), .Y(n239) );
  OAI21X1 U165 ( .A(n114), .B(n177), .C(\mem<24><0> ), .Y(n178) );
  OAI21X1 U166 ( .A(n114), .B(n119), .C(n178), .Y(n238) );
  NAND3X1 U167 ( .A(n166), .B(n13), .C(n165), .Y(n186) );
  OAI21X1 U168 ( .A(n3), .B(n116), .C(\mem<23><0> ), .Y(n179) );
  NAND2X1 U169 ( .A(n15), .B(n179), .Y(n237) );
  OAI21X1 U170 ( .A(n3), .B(n112), .C(\mem<22><0> ), .Y(n180) );
  NAND2X1 U171 ( .A(n17), .B(n180), .Y(n236) );
  OAI21X1 U172 ( .A(n3), .B(n107), .C(\mem<21><0> ), .Y(n181) );
  NAND2X1 U173 ( .A(n19), .B(n181), .Y(n235) );
  OAI21X1 U174 ( .A(n3), .B(n108), .C(\mem<20><0> ), .Y(n182) );
  NAND2X1 U175 ( .A(n21), .B(n182), .Y(n234) );
  OAI21X1 U176 ( .A(n3), .B(n109), .C(\mem<19><0> ), .Y(n183) );
  NAND2X1 U177 ( .A(n23), .B(n183), .Y(n233) );
  OAI21X1 U178 ( .A(n3), .B(n110), .C(\mem<18><0> ), .Y(n184) );
  NAND2X1 U179 ( .A(n25), .B(n184), .Y(n232) );
  OAI21X1 U180 ( .A(n3), .B(n111), .C(\mem<17><0> ), .Y(n185) );
  NAND2X1 U181 ( .A(n27), .B(n185), .Y(n231) );
  OAI21X1 U182 ( .A(n3), .B(n114), .C(\mem<16><0> ), .Y(n187) );
  NAND2X1 U183 ( .A(n29), .B(n187), .Y(n230) );
  OAI21X1 U184 ( .A(n7), .B(n116), .C(\mem<15><0> ), .Y(n188) );
  NAND2X1 U185 ( .A(n99), .B(n188), .Y(n229) );
  OAI21X1 U186 ( .A(n7), .B(n112), .C(\mem<14><0> ), .Y(n189) );
  NAND2X1 U187 ( .A(n32), .B(n189), .Y(n228) );
  OAI21X1 U188 ( .A(n7), .B(n107), .C(\mem<13><0> ), .Y(n190) );
  NAND2X1 U189 ( .A(n34), .B(n190), .Y(n227) );
  OAI21X1 U190 ( .A(n7), .B(n108), .C(\mem<12><0> ), .Y(n191) );
  NAND2X1 U191 ( .A(n36), .B(n191), .Y(n226) );
  OAI21X1 U192 ( .A(n7), .B(n109), .C(\mem<11><0> ), .Y(n192) );
  NAND2X1 U193 ( .A(n38), .B(n192), .Y(n225) );
  OAI21X1 U194 ( .A(n7), .B(n110), .C(\mem<10><0> ), .Y(n193) );
  NAND2X1 U195 ( .A(n40), .B(n193), .Y(n224) );
  OAI21X1 U196 ( .A(n7), .B(n111), .C(\mem<9><0> ), .Y(n194) );
  NAND2X1 U197 ( .A(n42), .B(n194), .Y(n223) );
  OAI21X1 U198 ( .A(n7), .B(n114), .C(\mem<8><0> ), .Y(n195) );
  NAND2X1 U199 ( .A(n44), .B(n195), .Y(n222) );
  OAI21X1 U200 ( .A(n6), .B(n116), .C(\mem<7><0> ), .Y(n196) );
  NAND2X1 U201 ( .A(n46), .B(n196), .Y(n221) );
  OAI21X1 U202 ( .A(n5), .B(n112), .C(\mem<6><0> ), .Y(n197) );
  NAND2X1 U203 ( .A(n48), .B(n197), .Y(n220) );
  OAI21X1 U204 ( .A(n6), .B(n107), .C(\mem<5><0> ), .Y(n200) );
  NAND2X1 U205 ( .A(n50), .B(n200), .Y(n219) );
  OAI21X1 U206 ( .A(n5), .B(n108), .C(\mem<4><0> ), .Y(n203) );
  NAND2X1 U207 ( .A(n52), .B(n203), .Y(n218) );
  OAI21X1 U208 ( .A(n6), .B(n109), .C(\mem<3><0> ), .Y(n206) );
  NAND2X1 U209 ( .A(n54), .B(n206), .Y(n217) );
  OAI21X1 U210 ( .A(n5), .B(n110), .C(\mem<2><0> ), .Y(n209) );
  NAND2X1 U211 ( .A(n56), .B(n209), .Y(n216) );
  OAI21X1 U212 ( .A(n6), .B(n111), .C(\mem<1><0> ), .Y(n212) );
  NAND2X1 U213 ( .A(n58), .B(n212), .Y(n215) );
  OAI21X1 U214 ( .A(n5), .B(n114), .C(\mem<0><0> ), .Y(n213) );
  NAND2X1 U215 ( .A(n60), .B(n213), .Y(n214) );
endmodule


module memv_0 ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n43, n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62,
         n63, n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83,
         n84, n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149,
         n150, n152, n169, n171, n187, n189, n205, n207, n223, n225, n241,
         n242, n244, n260, n262, n278, n280, n296, n298, n314, n315, n317,
         n333, n335, n351, n353, n354, n360, n362, n369, n374, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n1052), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n1053), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n1054), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n1055), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n1056), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n1057), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n1058), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n1059), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n1060), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n1061), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n1062), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n1063), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n1064), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n1065), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n1066), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n1067), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n1068), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n1069), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n1070), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n1071), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n1072), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n1073), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n1074), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n1075), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n1076), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n1077), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n1078), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n1079), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n1080), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n1081), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n1082), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n1083), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n1084), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n1085), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n1086), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n1087), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n1088), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n1089), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n1090), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n1091), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n1092), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n1093), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n1094), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n1095), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n1096), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n1097), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n1098), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n1099), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n1100), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n1101), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n1102), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n1103), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n1104), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n1105), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n1106), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n1107), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n1108), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n1109), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n1110), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n1111), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n1112), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n1113), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n1114), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n1115), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n1116), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n1117), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n1118), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n1119), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n1120), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n1121), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n1122), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n1123), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n1124), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n1125), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n1126), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n1127), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n1128), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n1129), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n1130), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n1131), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n1132), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n1133), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n1134), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n1135), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n1136), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n1137), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n1138), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n1139), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n1140), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n1141), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n1142), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n1143), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n1144), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n1145), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n1146), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n1147), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n1148), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n1149), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n1150), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n1151), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n1152), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n1153), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n1154), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n1155), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n1156), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n1157), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n1158), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n1159), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n1160), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n1161), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n1162), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n1163), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n1164), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n1165), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n1166), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n1167), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n1168), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n1169), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n1170), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n1171), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n1172), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n1173), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n1174), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n1175), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n1176), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n1177), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n1178), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n1179), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n1180), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n1181), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n1182), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n1183), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n1184), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n1185), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n1186), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n1187), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n1188), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n1189), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n1190), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n1191), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n1192), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n1193), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n1194), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n1195), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n1196), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n1197), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n1198), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n1199), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n1200), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n1201), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n1202), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n1203), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n1204), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n1205), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n1206), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n1207), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n1208), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n1209), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n1210), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n1211), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n1212), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n1213), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n1214), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n1215), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n1216), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n1217), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n1218), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n1219), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n1220), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n1221), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n1222), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n1223), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n1224), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n1225), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n1226), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n1227), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n1228), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n1229), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n1230), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n1231), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n1232), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n1233), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n1234), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n1235), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n1236), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n1237), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n1238), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n1239), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n1240), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n1241), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n1242), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n1243), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n1244), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n1245), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n1246), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n1247), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n1248), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n1249), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n1250), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n1251), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n1252), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n1253), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n1254), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n1255), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n1256), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n1257), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n1258), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n1259), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n1260), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n1261), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n1262), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n1263), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n1264), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n1265), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n1266), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n1267), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n1268), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n1269), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n1270), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n1271), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n1272), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n1273), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n1274), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n1275), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n1276), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n1277), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n1278), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n1279), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n1280), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n1281), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n1282), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n1283), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n1284), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n1285), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n1286), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n1287), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n1288), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n1289), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n1290), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n1291), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n1292), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n1293), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n1294), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n1295), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n1296), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n1297), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n1298), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n1299), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n1300), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n1301), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n1302), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n1303), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n1304), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n1305), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n1306), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n1307), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U6 ( .A(n797), .B(n794), .Y(n1326) );
  AND2X2 U7 ( .A(n797), .B(n795), .Y(n1319) );
  AND2X2 U8 ( .A(n789), .B(n683), .Y(n1325) );
  AND2X2 U9 ( .A(n789), .B(n782), .Y(n1323) );
  OAI21X1 U49 ( .A(n262), .B(n770), .C(n1572), .Y(n1307) );
  OAI21X1 U50 ( .A(n69), .B(n768), .C(\mem<255> ), .Y(n1572) );
  OAI21X1 U51 ( .A(n771), .B(n244), .C(n1571), .Y(n1306) );
  OAI21X1 U52 ( .A(n769), .B(n66), .C(\mem<254> ), .Y(n1571) );
  OAI21X1 U53 ( .A(n771), .B(n720), .C(n1570), .Y(n1305) );
  OAI21X1 U54 ( .A(n769), .B(n63), .C(\mem<253> ), .Y(n1570) );
  OAI21X1 U55 ( .A(n771), .B(n719), .C(n1569), .Y(n1304) );
  OAI21X1 U56 ( .A(n769), .B(n60), .C(\mem<252> ), .Y(n1569) );
  OAI21X1 U57 ( .A(n771), .B(n241), .C(n1568), .Y(n1303) );
  OAI21X1 U58 ( .A(n769), .B(n57), .C(\mem<251> ), .Y(n1568) );
  OAI21X1 U59 ( .A(n771), .B(n223), .C(n1567), .Y(n1302) );
  OAI21X1 U60 ( .A(n769), .B(n54), .C(\mem<250> ), .Y(n1567) );
  OAI21X1 U61 ( .A(n771), .B(n205), .C(n1566), .Y(n1301) );
  OAI21X1 U62 ( .A(n769), .B(n51), .C(\mem<249> ), .Y(n1566) );
  OAI21X1 U63 ( .A(n771), .B(n187), .C(n1565), .Y(n1300) );
  OAI21X1 U64 ( .A(n769), .B(n48), .C(\mem<248> ), .Y(n1565) );
  OAI21X1 U65 ( .A(n771), .B(n718), .C(n1564), .Y(n1299) );
  OAI21X1 U66 ( .A(n769), .B(n45), .C(\mem<247> ), .Y(n1564) );
  OAI21X1 U67 ( .A(n770), .B(n717), .C(n1563), .Y(n1298) );
  OAI21X1 U68 ( .A(n768), .B(n43), .C(\mem<246> ), .Y(n1563) );
  OAI21X1 U69 ( .A(n770), .B(n716), .C(n1562), .Y(n1297) );
  OAI21X1 U70 ( .A(n768), .B(n40), .C(\mem<245> ), .Y(n1562) );
  OAI21X1 U71 ( .A(n770), .B(n715), .C(n1561), .Y(n1296) );
  OAI21X1 U72 ( .A(n768), .B(n38), .C(\mem<244> ), .Y(n1561) );
  OAI21X1 U73 ( .A(n770), .B(n714), .C(n1560), .Y(n1295) );
  OAI21X1 U74 ( .A(n768), .B(n36), .C(\mem<243> ), .Y(n1560) );
  OAI21X1 U75 ( .A(n770), .B(n713), .C(n1559), .Y(n1294) );
  OAI21X1 U76 ( .A(n768), .B(n34), .C(\mem<242> ), .Y(n1559) );
  OAI21X1 U77 ( .A(n770), .B(n712), .C(n1558), .Y(n1293) );
  OAI21X1 U78 ( .A(n768), .B(n32), .C(\mem<241> ), .Y(n1558) );
  OAI21X1 U79 ( .A(n770), .B(n706), .C(n1557), .Y(n1292) );
  OAI21X1 U80 ( .A(n768), .B(n30), .C(\mem<240> ), .Y(n1557) );
  OAI21X1 U83 ( .A(n262), .B(n767), .C(n1553), .Y(n1291) );
  OAI21X1 U84 ( .A(n69), .B(n765), .C(\mem<239> ), .Y(n1553) );
  OAI21X1 U85 ( .A(n244), .B(n767), .C(n1552), .Y(n1290) );
  OAI21X1 U86 ( .A(n66), .B(n765), .C(\mem<238> ), .Y(n1552) );
  OAI21X1 U87 ( .A(n720), .B(n767), .C(n1551), .Y(n1289) );
  OAI21X1 U88 ( .A(n63), .B(n765), .C(\mem<237> ), .Y(n1551) );
  OAI21X1 U89 ( .A(n719), .B(n767), .C(n1550), .Y(n1288) );
  OAI21X1 U90 ( .A(n60), .B(n765), .C(\mem<236> ), .Y(n1550) );
  OAI21X1 U91 ( .A(n241), .B(n767), .C(n1549), .Y(n1287) );
  OAI21X1 U92 ( .A(n57), .B(n765), .C(\mem<235> ), .Y(n1549) );
  OAI21X1 U93 ( .A(n223), .B(n767), .C(n1548), .Y(n1286) );
  OAI21X1 U94 ( .A(n54), .B(n765), .C(\mem<234> ), .Y(n1548) );
  OAI21X1 U95 ( .A(n205), .B(n767), .C(n1547), .Y(n1285) );
  OAI21X1 U96 ( .A(n51), .B(n765), .C(\mem<233> ), .Y(n1547) );
  OAI21X1 U97 ( .A(n187), .B(n767), .C(n1546), .Y(n1284) );
  OAI21X1 U98 ( .A(n48), .B(n765), .C(\mem<232> ), .Y(n1546) );
  OAI21X1 U99 ( .A(n718), .B(n766), .C(n1545), .Y(n1283) );
  OAI21X1 U100 ( .A(n45), .B(n764), .C(\mem<231> ), .Y(n1545) );
  OAI21X1 U101 ( .A(n717), .B(n766), .C(n1544), .Y(n1282) );
  OAI21X1 U102 ( .A(n43), .B(n764), .C(\mem<230> ), .Y(n1544) );
  OAI21X1 U103 ( .A(n716), .B(n766), .C(n1543), .Y(n1281) );
  OAI21X1 U104 ( .A(n40), .B(n764), .C(\mem<229> ), .Y(n1543) );
  OAI21X1 U105 ( .A(n715), .B(n766), .C(n1542), .Y(n1280) );
  OAI21X1 U106 ( .A(n38), .B(n764), .C(\mem<228> ), .Y(n1542) );
  OAI21X1 U107 ( .A(n714), .B(n766), .C(n1541), .Y(n1279) );
  OAI21X1 U108 ( .A(n36), .B(n764), .C(\mem<227> ), .Y(n1541) );
  OAI21X1 U109 ( .A(n713), .B(n766), .C(n1540), .Y(n1278) );
  OAI21X1 U110 ( .A(n34), .B(n764), .C(\mem<226> ), .Y(n1540) );
  OAI21X1 U111 ( .A(n712), .B(n766), .C(n1539), .Y(n1277) );
  OAI21X1 U112 ( .A(n32), .B(n764), .C(\mem<225> ), .Y(n1539) );
  OAI21X1 U113 ( .A(n706), .B(n766), .C(n1538), .Y(n1276) );
  OAI21X1 U114 ( .A(n30), .B(n764), .C(\mem<224> ), .Y(n1538) );
  OAI21X1 U117 ( .A(n262), .B(n763), .C(n1536), .Y(n1275) );
  OAI21X1 U118 ( .A(n69), .B(n761), .C(\mem<223> ), .Y(n1536) );
  OAI21X1 U119 ( .A(n244), .B(n763), .C(n1535), .Y(n1274) );
  OAI21X1 U120 ( .A(n66), .B(n761), .C(\mem<222> ), .Y(n1535) );
  OAI21X1 U121 ( .A(n720), .B(n763), .C(n1534), .Y(n1273) );
  OAI21X1 U122 ( .A(n63), .B(n761), .C(\mem<221> ), .Y(n1534) );
  OAI21X1 U123 ( .A(n719), .B(n763), .C(n1533), .Y(n1272) );
  OAI21X1 U124 ( .A(n60), .B(n761), .C(\mem<220> ), .Y(n1533) );
  OAI21X1 U125 ( .A(n241), .B(n763), .C(n1532), .Y(n1271) );
  OAI21X1 U126 ( .A(n57), .B(n761), .C(\mem<219> ), .Y(n1532) );
  OAI21X1 U127 ( .A(n223), .B(n763), .C(n1531), .Y(n1270) );
  OAI21X1 U128 ( .A(n54), .B(n761), .C(\mem<218> ), .Y(n1531) );
  OAI21X1 U129 ( .A(n205), .B(n763), .C(n1530), .Y(n1269) );
  OAI21X1 U130 ( .A(n51), .B(n761), .C(\mem<217> ), .Y(n1530) );
  OAI21X1 U131 ( .A(n187), .B(n763), .C(n1529), .Y(n1268) );
  OAI21X1 U132 ( .A(n48), .B(n761), .C(\mem<216> ), .Y(n1529) );
  OAI21X1 U133 ( .A(n718), .B(n762), .C(n1528), .Y(n1267) );
  OAI21X1 U134 ( .A(n45), .B(n761), .C(\mem<215> ), .Y(n1528) );
  OAI21X1 U135 ( .A(n717), .B(n762), .C(n1527), .Y(n1266) );
  OAI21X1 U136 ( .A(n43), .B(n761), .C(\mem<214> ), .Y(n1527) );
  OAI21X1 U137 ( .A(n716), .B(n762), .C(n1526), .Y(n1265) );
  OAI21X1 U138 ( .A(n40), .B(n761), .C(\mem<213> ), .Y(n1526) );
  OAI21X1 U139 ( .A(n715), .B(n762), .C(n1525), .Y(n1264) );
  OAI21X1 U140 ( .A(n38), .B(n761), .C(\mem<212> ), .Y(n1525) );
  OAI21X1 U141 ( .A(n714), .B(n762), .C(n1524), .Y(n1263) );
  OAI21X1 U142 ( .A(n36), .B(n761), .C(\mem<211> ), .Y(n1524) );
  OAI21X1 U143 ( .A(n713), .B(n762), .C(n1523), .Y(n1262) );
  OAI21X1 U144 ( .A(n34), .B(n761), .C(\mem<210> ), .Y(n1523) );
  OAI21X1 U145 ( .A(n712), .B(n762), .C(n1522), .Y(n1261) );
  OAI21X1 U146 ( .A(n32), .B(n761), .C(\mem<209> ), .Y(n1522) );
  OAI21X1 U147 ( .A(n706), .B(n762), .C(n1521), .Y(n1260) );
  OAI21X1 U148 ( .A(n30), .B(n761), .C(\mem<208> ), .Y(n1521) );
  OAI21X1 U151 ( .A(n262), .B(n760), .C(n1520), .Y(n1259) );
  OAI21X1 U152 ( .A(n69), .B(n758), .C(\mem<207> ), .Y(n1520) );
  OAI21X1 U153 ( .A(n244), .B(n760), .C(n1519), .Y(n1258) );
  OAI21X1 U154 ( .A(n66), .B(n758), .C(\mem<206> ), .Y(n1519) );
  OAI21X1 U155 ( .A(n720), .B(n760), .C(n1518), .Y(n1257) );
  OAI21X1 U156 ( .A(n63), .B(n758), .C(\mem<205> ), .Y(n1518) );
  OAI21X1 U157 ( .A(n719), .B(n760), .C(n1517), .Y(n1256) );
  OAI21X1 U158 ( .A(n60), .B(n758), .C(\mem<204> ), .Y(n1517) );
  OAI21X1 U159 ( .A(n241), .B(n760), .C(n1516), .Y(n1255) );
  OAI21X1 U160 ( .A(n57), .B(n758), .C(\mem<203> ), .Y(n1516) );
  OAI21X1 U161 ( .A(n223), .B(n760), .C(n1515), .Y(n1254) );
  OAI21X1 U162 ( .A(n54), .B(n758), .C(\mem<202> ), .Y(n1515) );
  OAI21X1 U163 ( .A(n205), .B(n760), .C(n1514), .Y(n1253) );
  OAI21X1 U164 ( .A(n51), .B(n758), .C(\mem<201> ), .Y(n1514) );
  OAI21X1 U165 ( .A(n187), .B(n760), .C(n1513), .Y(n1252) );
  OAI21X1 U166 ( .A(n48), .B(n758), .C(\mem<200> ), .Y(n1513) );
  OAI21X1 U167 ( .A(n718), .B(n759), .C(n1512), .Y(n1251) );
  OAI21X1 U168 ( .A(n45), .B(n758), .C(\mem<199> ), .Y(n1512) );
  OAI21X1 U169 ( .A(n717), .B(n759), .C(n1511), .Y(n1250) );
  OAI21X1 U170 ( .A(n43), .B(n758), .C(\mem<198> ), .Y(n1511) );
  OAI21X1 U171 ( .A(n716), .B(n759), .C(n1510), .Y(n1249) );
  OAI21X1 U172 ( .A(n40), .B(n758), .C(\mem<197> ), .Y(n1510) );
  OAI21X1 U173 ( .A(n715), .B(n759), .C(n1509), .Y(n1248) );
  OAI21X1 U174 ( .A(n38), .B(n758), .C(\mem<196> ), .Y(n1509) );
  OAI21X1 U175 ( .A(n714), .B(n759), .C(n1508), .Y(n1247) );
  OAI21X1 U176 ( .A(n36), .B(n758), .C(\mem<195> ), .Y(n1508) );
  OAI21X1 U177 ( .A(n713), .B(n759), .C(n1507), .Y(n1246) );
  OAI21X1 U178 ( .A(n34), .B(n758), .C(\mem<194> ), .Y(n1507) );
  OAI21X1 U179 ( .A(n712), .B(n759), .C(n1506), .Y(n1245) );
  OAI21X1 U180 ( .A(n32), .B(n758), .C(\mem<193> ), .Y(n1506) );
  OAI21X1 U181 ( .A(n706), .B(n759), .C(n1505), .Y(n1244) );
  OAI21X1 U182 ( .A(n30), .B(n758), .C(\mem<192> ), .Y(n1505) );
  OAI21X1 U185 ( .A(n262), .B(n757), .C(n1504), .Y(n1243) );
  OAI21X1 U186 ( .A(n69), .B(n755), .C(\mem<191> ), .Y(n1504) );
  OAI21X1 U187 ( .A(n244), .B(n757), .C(n1503), .Y(n1242) );
  OAI21X1 U188 ( .A(n66), .B(n755), .C(\mem<190> ), .Y(n1503) );
  OAI21X1 U189 ( .A(n720), .B(n757), .C(n1502), .Y(n1241) );
  OAI21X1 U190 ( .A(n63), .B(n755), .C(\mem<189> ), .Y(n1502) );
  OAI21X1 U191 ( .A(n719), .B(n757), .C(n1501), .Y(n1240) );
  OAI21X1 U192 ( .A(n60), .B(n755), .C(\mem<188> ), .Y(n1501) );
  OAI21X1 U193 ( .A(n241), .B(n757), .C(n1500), .Y(n1239) );
  OAI21X1 U194 ( .A(n57), .B(n755), .C(\mem<187> ), .Y(n1500) );
  OAI21X1 U195 ( .A(n223), .B(n757), .C(n1499), .Y(n1238) );
  OAI21X1 U196 ( .A(n54), .B(n755), .C(\mem<186> ), .Y(n1499) );
  OAI21X1 U197 ( .A(n205), .B(n757), .C(n1498), .Y(n1237) );
  OAI21X1 U198 ( .A(n51), .B(n755), .C(\mem<185> ), .Y(n1498) );
  OAI21X1 U199 ( .A(n187), .B(n757), .C(n1497), .Y(n1236) );
  OAI21X1 U200 ( .A(n48), .B(n755), .C(\mem<184> ), .Y(n1497) );
  OAI21X1 U201 ( .A(n718), .B(n756), .C(n1496), .Y(n1235) );
  OAI21X1 U202 ( .A(n45), .B(n754), .C(\mem<183> ), .Y(n1496) );
  OAI21X1 U203 ( .A(n717), .B(n756), .C(n1495), .Y(n1234) );
  OAI21X1 U204 ( .A(n43), .B(n754), .C(\mem<182> ), .Y(n1495) );
  OAI21X1 U205 ( .A(n716), .B(n756), .C(n1494), .Y(n1233) );
  OAI21X1 U206 ( .A(n40), .B(n754), .C(\mem<181> ), .Y(n1494) );
  OAI21X1 U207 ( .A(n715), .B(n756), .C(n1493), .Y(n1232) );
  OAI21X1 U208 ( .A(n38), .B(n754), .C(\mem<180> ), .Y(n1493) );
  OAI21X1 U209 ( .A(n714), .B(n756), .C(n1492), .Y(n1231) );
  OAI21X1 U210 ( .A(n36), .B(n754), .C(\mem<179> ), .Y(n1492) );
  OAI21X1 U211 ( .A(n713), .B(n756), .C(n1491), .Y(n1230) );
  OAI21X1 U212 ( .A(n34), .B(n754), .C(\mem<178> ), .Y(n1491) );
  OAI21X1 U213 ( .A(n712), .B(n756), .C(n1490), .Y(n1229) );
  OAI21X1 U214 ( .A(n32), .B(n754), .C(\mem<177> ), .Y(n1490) );
  OAI21X1 U215 ( .A(n706), .B(n756), .C(n1489), .Y(n1228) );
  OAI21X1 U216 ( .A(n30), .B(n754), .C(\mem<176> ), .Y(n1489) );
  OAI21X1 U219 ( .A(n262), .B(n753), .C(n1487), .Y(n1227) );
  OAI21X1 U220 ( .A(n69), .B(n751), .C(\mem<175> ), .Y(n1487) );
  OAI21X1 U221 ( .A(n244), .B(n753), .C(n1486), .Y(n1226) );
  OAI21X1 U222 ( .A(n66), .B(n751), .C(\mem<174> ), .Y(n1486) );
  OAI21X1 U223 ( .A(n720), .B(n753), .C(n1485), .Y(n1225) );
  OAI21X1 U224 ( .A(n63), .B(n751), .C(\mem<173> ), .Y(n1485) );
  OAI21X1 U225 ( .A(n719), .B(n753), .C(n1484), .Y(n1224) );
  OAI21X1 U226 ( .A(n60), .B(n751), .C(\mem<172> ), .Y(n1484) );
  OAI21X1 U227 ( .A(n241), .B(n753), .C(n1483), .Y(n1223) );
  OAI21X1 U228 ( .A(n57), .B(n751), .C(\mem<171> ), .Y(n1483) );
  OAI21X1 U229 ( .A(n223), .B(n753), .C(n1482), .Y(n1222) );
  OAI21X1 U230 ( .A(n54), .B(n751), .C(\mem<170> ), .Y(n1482) );
  OAI21X1 U231 ( .A(n205), .B(n753), .C(n1481), .Y(n1221) );
  OAI21X1 U232 ( .A(n51), .B(n751), .C(\mem<169> ), .Y(n1481) );
  OAI21X1 U233 ( .A(n187), .B(n753), .C(n1480), .Y(n1220) );
  OAI21X1 U234 ( .A(n48), .B(n751), .C(\mem<168> ), .Y(n1480) );
  OAI21X1 U235 ( .A(n718), .B(n752), .C(n1479), .Y(n1219) );
  OAI21X1 U236 ( .A(n45), .B(n750), .C(\mem<167> ), .Y(n1479) );
  OAI21X1 U237 ( .A(n717), .B(n752), .C(n1478), .Y(n1218) );
  OAI21X1 U238 ( .A(n43), .B(n750), .C(\mem<166> ), .Y(n1478) );
  OAI21X1 U239 ( .A(n716), .B(n752), .C(n1477), .Y(n1217) );
  OAI21X1 U240 ( .A(n40), .B(n750), .C(\mem<165> ), .Y(n1477) );
  OAI21X1 U241 ( .A(n715), .B(n752), .C(n1476), .Y(n1216) );
  OAI21X1 U242 ( .A(n38), .B(n750), .C(\mem<164> ), .Y(n1476) );
  OAI21X1 U243 ( .A(n714), .B(n752), .C(n1475), .Y(n1215) );
  OAI21X1 U244 ( .A(n36), .B(n750), .C(\mem<163> ), .Y(n1475) );
  OAI21X1 U245 ( .A(n713), .B(n752), .C(n1474), .Y(n1214) );
  OAI21X1 U246 ( .A(n34), .B(n750), .C(\mem<162> ), .Y(n1474) );
  OAI21X1 U247 ( .A(n712), .B(n752), .C(n1473), .Y(n1213) );
  OAI21X1 U248 ( .A(n32), .B(n750), .C(\mem<161> ), .Y(n1473) );
  OAI21X1 U249 ( .A(n706), .B(n752), .C(n1472), .Y(n1212) );
  OAI21X1 U250 ( .A(n30), .B(n750), .C(\mem<160> ), .Y(n1472) );
  OAI21X1 U253 ( .A(n262), .B(n749), .C(n1471), .Y(n1211) );
  OAI21X1 U254 ( .A(n69), .B(n747), .C(\mem<159> ), .Y(n1471) );
  OAI21X1 U255 ( .A(n244), .B(n749), .C(n1470), .Y(n1210) );
  OAI21X1 U256 ( .A(n66), .B(n747), .C(\mem<158> ), .Y(n1470) );
  OAI21X1 U257 ( .A(n720), .B(n749), .C(n1469), .Y(n1209) );
  OAI21X1 U258 ( .A(n63), .B(n747), .C(\mem<157> ), .Y(n1469) );
  OAI21X1 U259 ( .A(n719), .B(n749), .C(n1468), .Y(n1208) );
  OAI21X1 U260 ( .A(n60), .B(n747), .C(\mem<156> ), .Y(n1468) );
  OAI21X1 U261 ( .A(n241), .B(n749), .C(n1467), .Y(n1207) );
  OAI21X1 U262 ( .A(n57), .B(n747), .C(\mem<155> ), .Y(n1467) );
  OAI21X1 U263 ( .A(n223), .B(n749), .C(n1466), .Y(n1206) );
  OAI21X1 U264 ( .A(n54), .B(n747), .C(\mem<154> ), .Y(n1466) );
  OAI21X1 U265 ( .A(n205), .B(n749), .C(n1465), .Y(n1205) );
  OAI21X1 U266 ( .A(n51), .B(n747), .C(\mem<153> ), .Y(n1465) );
  OAI21X1 U267 ( .A(n187), .B(n749), .C(n1464), .Y(n1204) );
  OAI21X1 U268 ( .A(n48), .B(n747), .C(\mem<152> ), .Y(n1464) );
  OAI21X1 U269 ( .A(n718), .B(n748), .C(n1463), .Y(n1203) );
  OAI21X1 U270 ( .A(n45), .B(n746), .C(\mem<151> ), .Y(n1463) );
  OAI21X1 U271 ( .A(n717), .B(n748), .C(n1462), .Y(n1202) );
  OAI21X1 U272 ( .A(n43), .B(n746), .C(\mem<150> ), .Y(n1462) );
  OAI21X1 U273 ( .A(n716), .B(n748), .C(n1461), .Y(n1201) );
  OAI21X1 U274 ( .A(n40), .B(n746), .C(\mem<149> ), .Y(n1461) );
  OAI21X1 U275 ( .A(n715), .B(n748), .C(n1460), .Y(n1200) );
  OAI21X1 U276 ( .A(n38), .B(n746), .C(\mem<148> ), .Y(n1460) );
  OAI21X1 U277 ( .A(n714), .B(n748), .C(n1459), .Y(n1199) );
  OAI21X1 U278 ( .A(n36), .B(n746), .C(\mem<147> ), .Y(n1459) );
  OAI21X1 U279 ( .A(n713), .B(n748), .C(n1458), .Y(n1198) );
  OAI21X1 U280 ( .A(n34), .B(n746), .C(\mem<146> ), .Y(n1458) );
  OAI21X1 U281 ( .A(n712), .B(n748), .C(n1457), .Y(n1197) );
  OAI21X1 U282 ( .A(n32), .B(n746), .C(\mem<145> ), .Y(n1457) );
  OAI21X1 U283 ( .A(n706), .B(n748), .C(n1456), .Y(n1196) );
  OAI21X1 U284 ( .A(n30), .B(n746), .C(\mem<144> ), .Y(n1456) );
  OAI21X1 U287 ( .A(n262), .B(n745), .C(n1455), .Y(n1195) );
  OAI21X1 U288 ( .A(n69), .B(n743), .C(\mem<143> ), .Y(n1455) );
  OAI21X1 U289 ( .A(n244), .B(n745), .C(n1454), .Y(n1194) );
  OAI21X1 U290 ( .A(n66), .B(n743), .C(\mem<142> ), .Y(n1454) );
  OAI21X1 U291 ( .A(n720), .B(n745), .C(n1453), .Y(n1193) );
  OAI21X1 U292 ( .A(n63), .B(n743), .C(\mem<141> ), .Y(n1453) );
  OAI21X1 U293 ( .A(n719), .B(n745), .C(n1452), .Y(n1192) );
  OAI21X1 U294 ( .A(n60), .B(n743), .C(\mem<140> ), .Y(n1452) );
  OAI21X1 U295 ( .A(n241), .B(n745), .C(n1451), .Y(n1191) );
  OAI21X1 U296 ( .A(n57), .B(n743), .C(\mem<139> ), .Y(n1451) );
  OAI21X1 U297 ( .A(n223), .B(n745), .C(n1450), .Y(n1190) );
  OAI21X1 U298 ( .A(n54), .B(n743), .C(\mem<138> ), .Y(n1450) );
  OAI21X1 U299 ( .A(n205), .B(n745), .C(n1449), .Y(n1189) );
  OAI21X1 U300 ( .A(n51), .B(n743), .C(\mem<137> ), .Y(n1449) );
  OAI21X1 U301 ( .A(n187), .B(n745), .C(n1448), .Y(n1188) );
  OAI21X1 U302 ( .A(n48), .B(n743), .C(\mem<136> ), .Y(n1448) );
  OAI21X1 U303 ( .A(n718), .B(n744), .C(n1447), .Y(n1187) );
  OAI21X1 U304 ( .A(n45), .B(n742), .C(\mem<135> ), .Y(n1447) );
  OAI21X1 U305 ( .A(n717), .B(n744), .C(n1446), .Y(n1186) );
  OAI21X1 U306 ( .A(n43), .B(n742), .C(\mem<134> ), .Y(n1446) );
  OAI21X1 U307 ( .A(n716), .B(n744), .C(n1445), .Y(n1185) );
  OAI21X1 U308 ( .A(n40), .B(n742), .C(\mem<133> ), .Y(n1445) );
  OAI21X1 U309 ( .A(n715), .B(n744), .C(n1444), .Y(n1184) );
  OAI21X1 U310 ( .A(n38), .B(n742), .C(\mem<132> ), .Y(n1444) );
  OAI21X1 U311 ( .A(n714), .B(n744), .C(n1443), .Y(n1183) );
  OAI21X1 U312 ( .A(n36), .B(n742), .C(\mem<131> ), .Y(n1443) );
  OAI21X1 U313 ( .A(n713), .B(n744), .C(n1442), .Y(n1182) );
  OAI21X1 U314 ( .A(n34), .B(n742), .C(\mem<130> ), .Y(n1442) );
  OAI21X1 U315 ( .A(n712), .B(n744), .C(n1441), .Y(n1181) );
  OAI21X1 U316 ( .A(n32), .B(n742), .C(\mem<129> ), .Y(n1441) );
  OAI21X1 U317 ( .A(n706), .B(n744), .C(n1440), .Y(n1180) );
  OAI21X1 U318 ( .A(n30), .B(n742), .C(\mem<128> ), .Y(n1440) );
  OAI21X1 U321 ( .A(n262), .B(n741), .C(n1439), .Y(n1179) );
  OAI21X1 U322 ( .A(n69), .B(n739), .C(\mem<127> ), .Y(n1439) );
  OAI21X1 U323 ( .A(n244), .B(n741), .C(n1438), .Y(n1178) );
  OAI21X1 U324 ( .A(n66), .B(n739), .C(\mem<126> ), .Y(n1438) );
  OAI21X1 U325 ( .A(n720), .B(n741), .C(n1437), .Y(n1177) );
  OAI21X1 U326 ( .A(n63), .B(n739), .C(\mem<125> ), .Y(n1437) );
  OAI21X1 U327 ( .A(n719), .B(n741), .C(n1436), .Y(n1176) );
  OAI21X1 U328 ( .A(n60), .B(n739), .C(\mem<124> ), .Y(n1436) );
  OAI21X1 U329 ( .A(n241), .B(n741), .C(n1435), .Y(n1175) );
  OAI21X1 U330 ( .A(n57), .B(n739), .C(\mem<123> ), .Y(n1435) );
  OAI21X1 U331 ( .A(n223), .B(n741), .C(n1434), .Y(n1174) );
  OAI21X1 U332 ( .A(n54), .B(n739), .C(\mem<122> ), .Y(n1434) );
  OAI21X1 U333 ( .A(n205), .B(n741), .C(n1433), .Y(n1173) );
  OAI21X1 U334 ( .A(n51), .B(n739), .C(\mem<121> ), .Y(n1433) );
  OAI21X1 U335 ( .A(n187), .B(n741), .C(n1432), .Y(n1172) );
  OAI21X1 U336 ( .A(n48), .B(n739), .C(\mem<120> ), .Y(n1432) );
  OAI21X1 U337 ( .A(n718), .B(n740), .C(n1431), .Y(n1171) );
  OAI21X1 U338 ( .A(n45), .B(n739), .C(\mem<119> ), .Y(n1431) );
  OAI21X1 U339 ( .A(n717), .B(n740), .C(n1430), .Y(n1170) );
  OAI21X1 U340 ( .A(n43), .B(n739), .C(\mem<118> ), .Y(n1430) );
  OAI21X1 U341 ( .A(n716), .B(n740), .C(n1429), .Y(n1169) );
  OAI21X1 U342 ( .A(n40), .B(n739), .C(\mem<117> ), .Y(n1429) );
  OAI21X1 U343 ( .A(n715), .B(n740), .C(n1428), .Y(n1168) );
  OAI21X1 U344 ( .A(n38), .B(n739), .C(\mem<116> ), .Y(n1428) );
  OAI21X1 U345 ( .A(n714), .B(n740), .C(n1427), .Y(n1167) );
  OAI21X1 U346 ( .A(n36), .B(n739), .C(\mem<115> ), .Y(n1427) );
  OAI21X1 U347 ( .A(n713), .B(n740), .C(n1426), .Y(n1166) );
  OAI21X1 U348 ( .A(n34), .B(n739), .C(\mem<114> ), .Y(n1426) );
  OAI21X1 U349 ( .A(n712), .B(n740), .C(n1425), .Y(n1165) );
  OAI21X1 U350 ( .A(n32), .B(n739), .C(\mem<113> ), .Y(n1425) );
  OAI21X1 U351 ( .A(n706), .B(n740), .C(n1424), .Y(n1164) );
  OAI21X1 U352 ( .A(n30), .B(n739), .C(\mem<112> ), .Y(n1424) );
  OAI21X1 U355 ( .A(n262), .B(n738), .C(n1423), .Y(n1163) );
  OAI21X1 U356 ( .A(n69), .B(n736), .C(\mem<111> ), .Y(n1423) );
  OAI21X1 U357 ( .A(n244), .B(n738), .C(n1422), .Y(n1162) );
  OAI21X1 U358 ( .A(n66), .B(n736), .C(\mem<110> ), .Y(n1422) );
  OAI21X1 U359 ( .A(n720), .B(n738), .C(n1421), .Y(n1161) );
  OAI21X1 U360 ( .A(n63), .B(n736), .C(\mem<109> ), .Y(n1421) );
  OAI21X1 U361 ( .A(n719), .B(n738), .C(n1420), .Y(n1160) );
  OAI21X1 U362 ( .A(n60), .B(n736), .C(\mem<108> ), .Y(n1420) );
  OAI21X1 U363 ( .A(n241), .B(n738), .C(n1419), .Y(n1159) );
  OAI21X1 U364 ( .A(n57), .B(n736), .C(\mem<107> ), .Y(n1419) );
  OAI21X1 U365 ( .A(n223), .B(n738), .C(n1418), .Y(n1158) );
  OAI21X1 U366 ( .A(n54), .B(n736), .C(\mem<106> ), .Y(n1418) );
  OAI21X1 U367 ( .A(n205), .B(n738), .C(n1417), .Y(n1157) );
  OAI21X1 U368 ( .A(n51), .B(n736), .C(\mem<105> ), .Y(n1417) );
  OAI21X1 U369 ( .A(n187), .B(n738), .C(n1416), .Y(n1156) );
  OAI21X1 U370 ( .A(n48), .B(n736), .C(\mem<104> ), .Y(n1416) );
  OAI21X1 U371 ( .A(n718), .B(n737), .C(n1415), .Y(n1155) );
  OAI21X1 U372 ( .A(n45), .B(n736), .C(\mem<103> ), .Y(n1415) );
  OAI21X1 U373 ( .A(n717), .B(n737), .C(n1414), .Y(n1154) );
  OAI21X1 U374 ( .A(n43), .B(n736), .C(\mem<102> ), .Y(n1414) );
  OAI21X1 U375 ( .A(n716), .B(n737), .C(n1413), .Y(n1153) );
  OAI21X1 U376 ( .A(n40), .B(n736), .C(\mem<101> ), .Y(n1413) );
  OAI21X1 U377 ( .A(n715), .B(n737), .C(n1412), .Y(n1152) );
  OAI21X1 U378 ( .A(n38), .B(n736), .C(\mem<100> ), .Y(n1412) );
  OAI21X1 U379 ( .A(n714), .B(n737), .C(n1411), .Y(n1151) );
  OAI21X1 U380 ( .A(n36), .B(n736), .C(\mem<99> ), .Y(n1411) );
  OAI21X1 U381 ( .A(n713), .B(n737), .C(n1410), .Y(n1150) );
  OAI21X1 U382 ( .A(n34), .B(n736), .C(\mem<98> ), .Y(n1410) );
  OAI21X1 U383 ( .A(n712), .B(n737), .C(n1409), .Y(n1149) );
  OAI21X1 U384 ( .A(n32), .B(n736), .C(\mem<97> ), .Y(n1409) );
  OAI21X1 U385 ( .A(n706), .B(n737), .C(n1408), .Y(n1148) );
  OAI21X1 U386 ( .A(n30), .B(n736), .C(\mem<96> ), .Y(n1408) );
  OAI21X1 U389 ( .A(n262), .B(n735), .C(n1407), .Y(n1147) );
  OAI21X1 U390 ( .A(n69), .B(n733), .C(\mem<95> ), .Y(n1407) );
  OAI21X1 U391 ( .A(n244), .B(n735), .C(n1406), .Y(n1146) );
  OAI21X1 U392 ( .A(n66), .B(n733), .C(\mem<94> ), .Y(n1406) );
  OAI21X1 U393 ( .A(n720), .B(n735), .C(n1405), .Y(n1145) );
  OAI21X1 U394 ( .A(n63), .B(n733), .C(\mem<93> ), .Y(n1405) );
  OAI21X1 U395 ( .A(n719), .B(n735), .C(n1404), .Y(n1144) );
  OAI21X1 U396 ( .A(n60), .B(n733), .C(\mem<92> ), .Y(n1404) );
  OAI21X1 U397 ( .A(n241), .B(n735), .C(n1403), .Y(n1143) );
  OAI21X1 U398 ( .A(n57), .B(n733), .C(\mem<91> ), .Y(n1403) );
  OAI21X1 U399 ( .A(n223), .B(n735), .C(n1402), .Y(n1142) );
  OAI21X1 U400 ( .A(n54), .B(n733), .C(\mem<90> ), .Y(n1402) );
  OAI21X1 U401 ( .A(n205), .B(n735), .C(n1401), .Y(n1141) );
  OAI21X1 U402 ( .A(n51), .B(n733), .C(\mem<89> ), .Y(n1401) );
  OAI21X1 U403 ( .A(n187), .B(n735), .C(n1400), .Y(n1140) );
  OAI21X1 U404 ( .A(n48), .B(n733), .C(\mem<88> ), .Y(n1400) );
  OAI21X1 U405 ( .A(n718), .B(n734), .C(n1399), .Y(n1139) );
  OAI21X1 U406 ( .A(n45), .B(n733), .C(\mem<87> ), .Y(n1399) );
  OAI21X1 U407 ( .A(n717), .B(n734), .C(n1398), .Y(n1138) );
  OAI21X1 U408 ( .A(n43), .B(n733), .C(\mem<86> ), .Y(n1398) );
  OAI21X1 U409 ( .A(n716), .B(n734), .C(n1397), .Y(n1137) );
  OAI21X1 U410 ( .A(n40), .B(n733), .C(\mem<85> ), .Y(n1397) );
  OAI21X1 U411 ( .A(n715), .B(n734), .C(n1396), .Y(n1136) );
  OAI21X1 U412 ( .A(n38), .B(n733), .C(\mem<84> ), .Y(n1396) );
  OAI21X1 U413 ( .A(n714), .B(n734), .C(n1395), .Y(n1135) );
  OAI21X1 U414 ( .A(n36), .B(n733), .C(\mem<83> ), .Y(n1395) );
  OAI21X1 U415 ( .A(n713), .B(n734), .C(n1394), .Y(n1134) );
  OAI21X1 U416 ( .A(n34), .B(n733), .C(\mem<82> ), .Y(n1394) );
  OAI21X1 U417 ( .A(n712), .B(n734), .C(n1393), .Y(n1133) );
  OAI21X1 U418 ( .A(n32), .B(n733), .C(\mem<81> ), .Y(n1393) );
  OAI21X1 U419 ( .A(n706), .B(n734), .C(n1392), .Y(n1132) );
  OAI21X1 U420 ( .A(n30), .B(n733), .C(\mem<80> ), .Y(n1392) );
  OAI21X1 U423 ( .A(n262), .B(n732), .C(n1391), .Y(n1131) );
  OAI21X1 U424 ( .A(n69), .B(n730), .C(\mem<79> ), .Y(n1391) );
  OAI21X1 U425 ( .A(n244), .B(n732), .C(n1390), .Y(n1130) );
  OAI21X1 U426 ( .A(n66), .B(n730), .C(\mem<78> ), .Y(n1390) );
  OAI21X1 U427 ( .A(n720), .B(n732), .C(n1389), .Y(n1129) );
  OAI21X1 U428 ( .A(n63), .B(n730), .C(\mem<77> ), .Y(n1389) );
  OAI21X1 U429 ( .A(n719), .B(n732), .C(n1388), .Y(n1128) );
  OAI21X1 U430 ( .A(n60), .B(n730), .C(\mem<76> ), .Y(n1388) );
  OAI21X1 U431 ( .A(n241), .B(n732), .C(n1387), .Y(n1127) );
  OAI21X1 U432 ( .A(n57), .B(n730), .C(\mem<75> ), .Y(n1387) );
  OAI21X1 U433 ( .A(n223), .B(n732), .C(n1386), .Y(n1126) );
  OAI21X1 U434 ( .A(n54), .B(n730), .C(\mem<74> ), .Y(n1386) );
  OAI21X1 U435 ( .A(n205), .B(n732), .C(n1385), .Y(n1125) );
  OAI21X1 U436 ( .A(n51), .B(n730), .C(\mem<73> ), .Y(n1385) );
  OAI21X1 U437 ( .A(n187), .B(n732), .C(n1384), .Y(n1124) );
  OAI21X1 U438 ( .A(n48), .B(n730), .C(\mem<72> ), .Y(n1384) );
  OAI21X1 U439 ( .A(n718), .B(n731), .C(n1383), .Y(n1123) );
  OAI21X1 U440 ( .A(n45), .B(n730), .C(\mem<71> ), .Y(n1383) );
  OAI21X1 U441 ( .A(n717), .B(n731), .C(n1382), .Y(n1122) );
  OAI21X1 U442 ( .A(n43), .B(n730), .C(\mem<70> ), .Y(n1382) );
  OAI21X1 U443 ( .A(n716), .B(n731), .C(n1381), .Y(n1121) );
  OAI21X1 U444 ( .A(n40), .B(n730), .C(\mem<69> ), .Y(n1381) );
  OAI21X1 U445 ( .A(n715), .B(n731), .C(n1380), .Y(n1120) );
  OAI21X1 U446 ( .A(n38), .B(n730), .C(\mem<68> ), .Y(n1380) );
  OAI21X1 U447 ( .A(n714), .B(n731), .C(n1379), .Y(n1119) );
  OAI21X1 U448 ( .A(n36), .B(n730), .C(\mem<67> ), .Y(n1379) );
  OAI21X1 U449 ( .A(n713), .B(n731), .C(n1378), .Y(n1118) );
  OAI21X1 U450 ( .A(n34), .B(n730), .C(\mem<66> ), .Y(n1378) );
  OAI21X1 U451 ( .A(n712), .B(n731), .C(n1377), .Y(n1117) );
  OAI21X1 U452 ( .A(n32), .B(n730), .C(\mem<65> ), .Y(n1377) );
  OAI21X1 U453 ( .A(n706), .B(n731), .C(n1376), .Y(n1116) );
  OAI21X1 U454 ( .A(n30), .B(n730), .C(\mem<64> ), .Y(n1376) );
  OAI21X1 U458 ( .A(n262), .B(n729), .C(n1375), .Y(n1115) );
  OAI21X1 U459 ( .A(n69), .B(n727), .C(\mem<63> ), .Y(n1375) );
  OAI21X1 U460 ( .A(n244), .B(n729), .C(n1374), .Y(n1114) );
  OAI21X1 U461 ( .A(n66), .B(n727), .C(\mem<62> ), .Y(n1374) );
  OAI21X1 U462 ( .A(n720), .B(n729), .C(n1373), .Y(n1113) );
  OAI21X1 U463 ( .A(n63), .B(n727), .C(\mem<61> ), .Y(n1373) );
  OAI21X1 U464 ( .A(n719), .B(n729), .C(n1372), .Y(n1112) );
  OAI21X1 U465 ( .A(n60), .B(n727), .C(\mem<60> ), .Y(n1372) );
  OAI21X1 U466 ( .A(n241), .B(n729), .C(n1371), .Y(n1111) );
  OAI21X1 U467 ( .A(n57), .B(n727), .C(\mem<59> ), .Y(n1371) );
  OAI21X1 U468 ( .A(n223), .B(n729), .C(n1370), .Y(n1110) );
  OAI21X1 U469 ( .A(n54), .B(n727), .C(\mem<58> ), .Y(n1370) );
  OAI21X1 U470 ( .A(n205), .B(n729), .C(n1369), .Y(n1109) );
  OAI21X1 U471 ( .A(n51), .B(n727), .C(\mem<57> ), .Y(n1369) );
  OAI21X1 U472 ( .A(n187), .B(n729), .C(n1368), .Y(n1108) );
  OAI21X1 U473 ( .A(n48), .B(n727), .C(\mem<56> ), .Y(n1368) );
  OAI21X1 U474 ( .A(n718), .B(n728), .C(n1367), .Y(n1107) );
  OAI21X1 U475 ( .A(n45), .B(n727), .C(\mem<55> ), .Y(n1367) );
  OAI21X1 U476 ( .A(n717), .B(n728), .C(n1366), .Y(n1106) );
  OAI21X1 U477 ( .A(n43), .B(n727), .C(\mem<54> ), .Y(n1366) );
  OAI21X1 U478 ( .A(n716), .B(n728), .C(n1365), .Y(n1105) );
  OAI21X1 U479 ( .A(n40), .B(n727), .C(\mem<53> ), .Y(n1365) );
  OAI21X1 U480 ( .A(n715), .B(n728), .C(n1364), .Y(n1104) );
  OAI21X1 U481 ( .A(n38), .B(n727), .C(\mem<52> ), .Y(n1364) );
  OAI21X1 U482 ( .A(n714), .B(n728), .C(n1363), .Y(n1103) );
  OAI21X1 U483 ( .A(n36), .B(n727), .C(\mem<51> ), .Y(n1363) );
  OAI21X1 U484 ( .A(n713), .B(n728), .C(n1362), .Y(n1102) );
  OAI21X1 U485 ( .A(n34), .B(n727), .C(\mem<50> ), .Y(n1362) );
  OAI21X1 U486 ( .A(n712), .B(n728), .C(n1361), .Y(n1101) );
  OAI21X1 U487 ( .A(n32), .B(n727), .C(\mem<49> ), .Y(n1361) );
  OAI21X1 U488 ( .A(n706), .B(n728), .C(n1360), .Y(n1100) );
  OAI21X1 U489 ( .A(n30), .B(n727), .C(\mem<48> ), .Y(n1360) );
  OAI21X1 U492 ( .A(n262), .B(n726), .C(n1359), .Y(n1099) );
  OAI21X1 U493 ( .A(n69), .B(n724), .C(\mem<47> ), .Y(n1359) );
  OAI21X1 U494 ( .A(n244), .B(n726), .C(n1358), .Y(n1098) );
  OAI21X1 U495 ( .A(n66), .B(n724), .C(\mem<46> ), .Y(n1358) );
  OAI21X1 U496 ( .A(n720), .B(n726), .C(n1357), .Y(n1097) );
  OAI21X1 U497 ( .A(n63), .B(n724), .C(\mem<45> ), .Y(n1357) );
  OAI21X1 U498 ( .A(n719), .B(n726), .C(n1356), .Y(n1096) );
  OAI21X1 U499 ( .A(n60), .B(n724), .C(\mem<44> ), .Y(n1356) );
  OAI21X1 U500 ( .A(n241), .B(n726), .C(n1355), .Y(n1095) );
  OAI21X1 U501 ( .A(n57), .B(n724), .C(\mem<43> ), .Y(n1355) );
  OAI21X1 U502 ( .A(n223), .B(n726), .C(n1354), .Y(n1094) );
  OAI21X1 U503 ( .A(n54), .B(n724), .C(\mem<42> ), .Y(n1354) );
  OAI21X1 U504 ( .A(n205), .B(n726), .C(n1353), .Y(n1093) );
  OAI21X1 U505 ( .A(n51), .B(n724), .C(\mem<41> ), .Y(n1353) );
  OAI21X1 U506 ( .A(n187), .B(n726), .C(n1352), .Y(n1092) );
  OAI21X1 U507 ( .A(n48), .B(n724), .C(\mem<40> ), .Y(n1352) );
  OAI21X1 U508 ( .A(n718), .B(n725), .C(n1351), .Y(n1091) );
  OAI21X1 U509 ( .A(n45), .B(n724), .C(\mem<39> ), .Y(n1351) );
  OAI21X1 U510 ( .A(n717), .B(n725), .C(n1350), .Y(n1090) );
  OAI21X1 U511 ( .A(n43), .B(n724), .C(\mem<38> ), .Y(n1350) );
  OAI21X1 U512 ( .A(n716), .B(n725), .C(n1349), .Y(n1089) );
  OAI21X1 U513 ( .A(n40), .B(n724), .C(\mem<37> ), .Y(n1349) );
  OAI21X1 U514 ( .A(n715), .B(n725), .C(n1348), .Y(n1088) );
  OAI21X1 U515 ( .A(n38), .B(n724), .C(\mem<36> ), .Y(n1348) );
  OAI21X1 U516 ( .A(n714), .B(n725), .C(n1347), .Y(n1087) );
  OAI21X1 U517 ( .A(n36), .B(n724), .C(\mem<35> ), .Y(n1347) );
  OAI21X1 U518 ( .A(n713), .B(n725), .C(n1346), .Y(n1086) );
  OAI21X1 U519 ( .A(n34), .B(n724), .C(\mem<34> ), .Y(n1346) );
  OAI21X1 U520 ( .A(n712), .B(n725), .C(n1345), .Y(n1085) );
  OAI21X1 U521 ( .A(n32), .B(n724), .C(\mem<33> ), .Y(n1345) );
  OAI21X1 U522 ( .A(n706), .B(n725), .C(n1344), .Y(n1084) );
  OAI21X1 U523 ( .A(n30), .B(n724), .C(\mem<32> ), .Y(n1344) );
  OAI21X1 U526 ( .A(n262), .B(n723), .C(n1343), .Y(n1083) );
  OAI21X1 U527 ( .A(n69), .B(n721), .C(\mem<31> ), .Y(n1343) );
  OAI21X1 U528 ( .A(n244), .B(n723), .C(n1342), .Y(n1082) );
  OAI21X1 U529 ( .A(n66), .B(n721), .C(\mem<30> ), .Y(n1342) );
  OAI21X1 U530 ( .A(n720), .B(n723), .C(n1341), .Y(n1081) );
  OAI21X1 U531 ( .A(n63), .B(n721), .C(\mem<29> ), .Y(n1341) );
  OAI21X1 U532 ( .A(n719), .B(n723), .C(n1340), .Y(n1080) );
  OAI21X1 U533 ( .A(n60), .B(n721), .C(\mem<28> ), .Y(n1340) );
  OAI21X1 U534 ( .A(n241), .B(n723), .C(n1339), .Y(n1079) );
  OAI21X1 U535 ( .A(n57), .B(n721), .C(\mem<27> ), .Y(n1339) );
  OAI21X1 U536 ( .A(n223), .B(n723), .C(n1338), .Y(n1078) );
  OAI21X1 U537 ( .A(n54), .B(n721), .C(\mem<26> ), .Y(n1338) );
  OAI21X1 U538 ( .A(n205), .B(n723), .C(n1337), .Y(n1077) );
  OAI21X1 U539 ( .A(n51), .B(n721), .C(\mem<25> ), .Y(n1337) );
  OAI21X1 U540 ( .A(n187), .B(n723), .C(n1336), .Y(n1076) );
  OAI21X1 U541 ( .A(n48), .B(n721), .C(\mem<24> ), .Y(n1336) );
  OAI21X1 U542 ( .A(n718), .B(n722), .C(n1335), .Y(n1075) );
  OAI21X1 U543 ( .A(n45), .B(n721), .C(\mem<23> ), .Y(n1335) );
  OAI21X1 U544 ( .A(n717), .B(n722), .C(n1334), .Y(n1074) );
  OAI21X1 U545 ( .A(n43), .B(n721), .C(\mem<22> ), .Y(n1334) );
  OAI21X1 U546 ( .A(n716), .B(n722), .C(n1333), .Y(n1073) );
  OAI21X1 U547 ( .A(n40), .B(n721), .C(\mem<21> ), .Y(n1333) );
  OAI21X1 U548 ( .A(n715), .B(n722), .C(n1332), .Y(n1072) );
  OAI21X1 U549 ( .A(n38), .B(n721), .C(\mem<20> ), .Y(n1332) );
  OAI21X1 U550 ( .A(n714), .B(n722), .C(n1331), .Y(n1071) );
  OAI21X1 U551 ( .A(n36), .B(n721), .C(\mem<19> ), .Y(n1331) );
  OAI21X1 U552 ( .A(n713), .B(n722), .C(n1330), .Y(n1070) );
  OAI21X1 U553 ( .A(n34), .B(n721), .C(\mem<18> ), .Y(n1330) );
  OAI21X1 U554 ( .A(n712), .B(n722), .C(n1329), .Y(n1069) );
  OAI21X1 U555 ( .A(n32), .B(n721), .C(\mem<17> ), .Y(n1329) );
  OAI21X1 U556 ( .A(n706), .B(n722), .C(n1328), .Y(n1068) );
  OAI21X1 U557 ( .A(n30), .B(n721), .C(\mem<16> ), .Y(n1328) );
  OAI21X1 U561 ( .A(n262), .B(n711), .C(n1327), .Y(n1067) );
  OAI21X1 U562 ( .A(n69), .B(n707), .C(\mem<15> ), .Y(n1327) );
  OAI21X1 U565 ( .A(n244), .B(n711), .C(n1324), .Y(n1066) );
  OAI21X1 U566 ( .A(n66), .B(n707), .C(\mem<14> ), .Y(n1324) );
  OAI21X1 U569 ( .A(n720), .B(n711), .C(n1322), .Y(n1065) );
  OAI21X1 U570 ( .A(n63), .B(n707), .C(\mem<13> ), .Y(n1322) );
  OAI21X1 U573 ( .A(n719), .B(n711), .C(n1321), .Y(n1064) );
  OAI21X1 U574 ( .A(n60), .B(n707), .C(\mem<12> ), .Y(n1321) );
  OAI21X1 U577 ( .A(n241), .B(n711), .C(n1320), .Y(n1063) );
  OAI21X1 U578 ( .A(n57), .B(n707), .C(\mem<11> ), .Y(n1320) );
  OAI21X1 U581 ( .A(n223), .B(n711), .C(n1318), .Y(n1062) );
  OAI21X1 U582 ( .A(n54), .B(n707), .C(\mem<10> ), .Y(n1318) );
  OAI21X1 U585 ( .A(n205), .B(n711), .C(n1317), .Y(n1061) );
  OAI21X1 U586 ( .A(n51), .B(n707), .C(\mem<9> ), .Y(n1317) );
  OAI21X1 U589 ( .A(n187), .B(n711), .C(n1316), .Y(n1060) );
  OAI21X1 U590 ( .A(n48), .B(n707), .C(\mem<8> ), .Y(n1316) );
  OAI21X1 U593 ( .A(n718), .B(n710), .C(n1315), .Y(n1059) );
  OAI21X1 U594 ( .A(n45), .B(n707), .C(\mem<7> ), .Y(n1315) );
  OAI21X1 U597 ( .A(n717), .B(n710), .C(n1314), .Y(n1058) );
  OAI21X1 U598 ( .A(n43), .B(n707), .C(\mem<6> ), .Y(n1314) );
  OAI21X1 U601 ( .A(n716), .B(n710), .C(n1313), .Y(n1057) );
  OAI21X1 U602 ( .A(n40), .B(n707), .C(\mem<5> ), .Y(n1313) );
  OAI21X1 U605 ( .A(n715), .B(n710), .C(n1312), .Y(n1056) );
  OAI21X1 U606 ( .A(n38), .B(n707), .C(\mem<4> ), .Y(n1312) );
  OAI21X1 U610 ( .A(n714), .B(n710), .C(n1311), .Y(n1055) );
  OAI21X1 U611 ( .A(n36), .B(n707), .C(\mem<3> ), .Y(n1311) );
  OAI21X1 U614 ( .A(n713), .B(n710), .C(n1310), .Y(n1054) );
  OAI21X1 U615 ( .A(n34), .B(n707), .C(\mem<2> ), .Y(n1310) );
  OAI21X1 U618 ( .A(n712), .B(n710), .C(n1309), .Y(n1053) );
  OAI21X1 U619 ( .A(n32), .B(n707), .C(\mem<1> ), .Y(n1309) );
  OAI21X1 U623 ( .A(n706), .B(n710), .C(n1308), .Y(n1052) );
  OAI21X1 U624 ( .A(n30), .B(n707), .C(\mem<0> ), .Y(n1308) );
  INVX1 U2 ( .A(n694), .Y(n1) );
  BUFX4 U3 ( .A(n775), .Y(n694) );
  INVX1 U4 ( .A(n783), .Y(n682) );
  INVX2 U5 ( .A(n783), .Y(n683) );
  INVX8 U10 ( .A(n783), .Y(n777) );
  INVX8 U11 ( .A(n783), .Y(n781) );
  AND2X2 U12 ( .A(n863), .B(n785), .Y(n13) );
  AND2X2 U13 ( .A(n921), .B(n704), .Y(n9) );
  INVX2 U14 ( .A(n774), .Y(n698) );
  AND2X1 U15 ( .A(n983), .B(N23), .Y(n27) );
  INVX1 U16 ( .A(\mem<113> ), .Y(n703) );
  INVX1 U17 ( .A(\mem<112> ), .Y(n702) );
  INVX1 U18 ( .A(n786), .Y(n679) );
  INVX1 U19 ( .A(n701), .Y(n905) );
  AND2X1 U20 ( .A(N25), .B(n800), .Y(n1488) );
  AND2X1 U21 ( .A(data_in), .B(n709), .Y(n1556) );
  AND2X1 U22 ( .A(N25), .B(N24), .Y(n1555) );
  BUFX2 U23 ( .A(n1556), .Y(n773) );
  AND2X1 U24 ( .A(N23), .B(N22), .Y(n1554) );
  AND2X1 U25 ( .A(N23), .B(n799), .Y(n1537) );
  BUFX2 U26 ( .A(n1556), .Y(n772) );
  BUFX2 U27 ( .A(n150), .Y(n709) );
  BUFX2 U28 ( .A(n150), .Y(n708) );
  BUFX2 U29 ( .A(n659), .Y(n771) );
  BUFX2 U30 ( .A(n657), .Y(n768) );
  BUFX2 U31 ( .A(n659), .Y(n770) );
  BUFX2 U32 ( .A(n655), .Y(n767) );
  BUFX2 U33 ( .A(n653), .Y(n764) );
  BUFX2 U34 ( .A(n655), .Y(n766) );
  BUFX2 U35 ( .A(n651), .Y(n763) );
  BUFX2 U36 ( .A(n651), .Y(n762) );
  BUFX2 U37 ( .A(n649), .Y(n760) );
  BUFX2 U38 ( .A(n649), .Y(n759) );
  BUFX2 U39 ( .A(n647), .Y(n757) );
  BUFX2 U40 ( .A(n645), .Y(n754) );
  BUFX2 U41 ( .A(n647), .Y(n756) );
  BUFX2 U42 ( .A(n643), .Y(n753) );
  BUFX2 U43 ( .A(n641), .Y(n750) );
  BUFX2 U44 ( .A(n643), .Y(n752) );
  BUFX2 U45 ( .A(n639), .Y(n749) );
  BUFX2 U46 ( .A(n637), .Y(n746) );
  BUFX2 U47 ( .A(n639), .Y(n748) );
  BUFX2 U48 ( .A(n635), .Y(n745) );
  BUFX2 U81 ( .A(n374), .Y(n742) );
  BUFX2 U82 ( .A(n635), .Y(n744) );
  BUFX2 U115 ( .A(n362), .Y(n741) );
  BUFX2 U116 ( .A(n362), .Y(n740) );
  BUFX2 U149 ( .A(n354), .Y(n738) );
  BUFX2 U150 ( .A(n354), .Y(n737) );
  BUFX2 U183 ( .A(n351), .Y(n735) );
  BUFX2 U184 ( .A(n351), .Y(n734) );
  BUFX2 U217 ( .A(n333), .Y(n732) );
  BUFX2 U218 ( .A(n333), .Y(n731) );
  BUFX2 U251 ( .A(n315), .Y(n729) );
  BUFX2 U252 ( .A(n315), .Y(n728) );
  BUFX2 U285 ( .A(n298), .Y(n726) );
  BUFX2 U286 ( .A(n298), .Y(n725) );
  BUFX2 U319 ( .A(n280), .Y(n723) );
  BUFX2 U320 ( .A(n280), .Y(n722) );
  BUFX2 U353 ( .A(n169), .Y(n711) );
  BUFX2 U354 ( .A(n169), .Y(n710) );
  INVX1 U387 ( .A(n792), .Y(n676) );
  INVX1 U388 ( .A(n692), .Y(n690) );
  INVX1 U421 ( .A(n72), .Y(n707) );
  INVX1 U422 ( .A(n87), .Y(n721) );
  INVX1 U455 ( .A(n95), .Y(n730) );
  INVX1 U456 ( .A(n112), .Y(n733) );
  INVX1 U457 ( .A(n131), .Y(n758) );
  INVX1 U490 ( .A(n133), .Y(n761) );
  INVX1 U491 ( .A(n84), .Y(n719) );
  INVX1 U524 ( .A(n86), .Y(n720) );
  INVX1 U525 ( .A(n89), .Y(n724) );
  INVX1 U558 ( .A(n114), .Y(n736) );
  INVX1 U559 ( .A(n93), .Y(n727) );
  INVX1 U560 ( .A(n130), .Y(n739) );
  BUFX2 U563 ( .A(n374), .Y(n743) );
  BUFX2 U564 ( .A(n637), .Y(n747) );
  BUFX2 U567 ( .A(n641), .Y(n751) );
  BUFX2 U568 ( .A(n645), .Y(n755) );
  BUFX2 U571 ( .A(n653), .Y(n765) );
  BUFX2 U572 ( .A(n657), .Y(n769) );
  INVX1 U575 ( .A(n71), .Y(n706) );
  INVX1 U576 ( .A(n74), .Y(n712) );
  INVX1 U579 ( .A(n75), .Y(n713) );
  INVX1 U580 ( .A(n77), .Y(n714) );
  INVX1 U583 ( .A(n78), .Y(n715) );
  INVX1 U584 ( .A(n80), .Y(n716) );
  INVX1 U587 ( .A(n81), .Y(n717) );
  INVX1 U588 ( .A(n83), .Y(n718) );
  INVX4 U591 ( .A(N18), .Y(n775) );
  AND2X2 U592 ( .A(n16), .B(n26), .Y(n2) );
  AND2X2 U595 ( .A(N21), .B(n856), .Y(n3) );
  INVX1 U596 ( .A(n3), .Y(n4) );
  AND2X2 U599 ( .A(n18), .B(n4), .Y(n5) );
  AND2X2 U600 ( .A(n28), .B(n20), .Y(n6) );
  AND2X2 U603 ( .A(n10), .B(n22), .Y(n7) );
  AND2X2 U604 ( .A(n12), .B(n14), .Y(n8) );
  INVX1 U607 ( .A(n9), .Y(n10) );
  AND2X2 U608 ( .A(n864), .B(n705), .Y(n11) );
  INVX1 U609 ( .A(n11), .Y(n12) );
  INVX1 U612 ( .A(n13), .Y(n14) );
  AND2X2 U613 ( .A(n818), .B(n691), .Y(n15) );
  INVX1 U616 ( .A(n15), .Y(n16) );
  AND2X1 U617 ( .A(n857), .B(n700), .Y(n17) );
  INVX1 U620 ( .A(n17), .Y(n18) );
  AND2X1 U621 ( .A(n984), .B(n704), .Y(n19) );
  INVX1 U622 ( .A(n19), .Y(n20) );
  AND2X1 U625 ( .A(n920), .B(N23), .Y(n21) );
  INVX1 U626 ( .A(n21), .Y(n22) );
  OR2X1 U627 ( .A(rst), .B(write), .Y(n23) );
  INVX1 U628 ( .A(n23), .Y(n24) );
  AND2X1 U629 ( .A(n817), .B(n784), .Y(n25) );
  INVX1 U630 ( .A(n25), .Y(n26) );
  INVX1 U631 ( .A(n27), .Y(n28) );
  AND2X1 U632 ( .A(n71), .B(n708), .Y(n29) );
  INVX1 U633 ( .A(n29), .Y(n30) );
  AND2X1 U634 ( .A(n74), .B(n708), .Y(n31) );
  INVX1 U635 ( .A(n31), .Y(n32) );
  AND2X1 U636 ( .A(n75), .B(n708), .Y(n33) );
  INVX1 U637 ( .A(n33), .Y(n34) );
  AND2X1 U638 ( .A(n77), .B(n708), .Y(n35) );
  INVX1 U639 ( .A(n35), .Y(n36) );
  AND2X1 U640 ( .A(n78), .B(n708), .Y(n37) );
  INVX1 U641 ( .A(n37), .Y(n38) );
  AND2X1 U642 ( .A(n80), .B(n708), .Y(n39) );
  INVX1 U643 ( .A(n39), .Y(n40) );
  AND2X1 U644 ( .A(n81), .B(n708), .Y(n41) );
  INVX1 U645 ( .A(n41), .Y(n43) );
  AND2X1 U646 ( .A(n83), .B(n708), .Y(n44) );
  INVX1 U647 ( .A(n44), .Y(n45) );
  AND2X1 U648 ( .A(n171), .B(n709), .Y(n47) );
  INVX1 U649 ( .A(n47), .Y(n48) );
  AND2X1 U650 ( .A(n189), .B(n709), .Y(n50) );
  INVX1 U651 ( .A(n50), .Y(n51) );
  AND2X1 U652 ( .A(n207), .B(n709), .Y(n53) );
  INVX1 U653 ( .A(n53), .Y(n54) );
  AND2X1 U654 ( .A(n225), .B(n709), .Y(n56) );
  INVX1 U655 ( .A(n56), .Y(n57) );
  AND2X1 U656 ( .A(n84), .B(n709), .Y(n59) );
  INVX1 U657 ( .A(n59), .Y(n60) );
  AND2X1 U658 ( .A(n86), .B(n709), .Y(n62) );
  INVX1 U659 ( .A(n62), .Y(n63) );
  AND2X1 U660 ( .A(n242), .B(n709), .Y(n65) );
  INVX1 U661 ( .A(n65), .Y(n66) );
  AND2X1 U662 ( .A(n260), .B(n709), .Y(n68) );
  INVX1 U663 ( .A(n68), .Y(n69) );
  AND2X1 U664 ( .A(n669), .B(n661), .Y(n71) );
  AND2X1 U665 ( .A(n671), .B(n663), .Y(n72) );
  AND2X1 U666 ( .A(n669), .B(n665), .Y(n74) );
  AND2X1 U667 ( .A(n669), .B(n1323), .Y(n75) );
  AND2X1 U668 ( .A(n669), .B(n1325), .Y(n77) );
  AND2X1 U669 ( .A(n673), .B(n661), .Y(n78) );
  AND2X1 U670 ( .A(n673), .B(n665), .Y(n80) );
  AND2X1 U671 ( .A(n673), .B(n1323), .Y(n81) );
  AND2X1 U672 ( .A(n673), .B(n1325), .Y(n83) );
  AND2X1 U673 ( .A(n661), .B(n1326), .Y(n84) );
  AND2X1 U674 ( .A(n665), .B(n1326), .Y(n86) );
  AND2X1 U675 ( .A(n671), .B(n667), .Y(n87) );
  AND2X1 U676 ( .A(n671), .B(n1537), .Y(n89) );
  AND2X1 U677 ( .A(n671), .B(n1554), .Y(n93) );
  AND2X1 U678 ( .A(n675), .B(n663), .Y(n95) );
  AND2X1 U679 ( .A(n675), .B(n667), .Y(n112) );
  AND2X1 U680 ( .A(n675), .B(n1537), .Y(n114) );
  AND2X1 U681 ( .A(n675), .B(n1554), .Y(n130) );
  AND2X1 U682 ( .A(n663), .B(n1555), .Y(n131) );
  AND2X1 U683 ( .A(n667), .B(n1555), .Y(n133) );
  OR2X1 U684 ( .A(n1051), .B(rst), .Y(n149) );
  INVX1 U685 ( .A(n149), .Y(n150) );
  AND2X1 U686 ( .A(n72), .B(n772), .Y(n152) );
  INVX1 U687 ( .A(n152), .Y(n169) );
  AND2X1 U688 ( .A(n1319), .B(n661), .Y(n171) );
  INVX1 U689 ( .A(n171), .Y(n187) );
  AND2X1 U690 ( .A(n1319), .B(n665), .Y(n189) );
  INVX1 U691 ( .A(n189), .Y(n205) );
  AND2X1 U692 ( .A(n1319), .B(n1323), .Y(n207) );
  INVX1 U693 ( .A(n207), .Y(n223) );
  AND2X1 U694 ( .A(n1319), .B(n1325), .Y(n225) );
  INVX1 U695 ( .A(n225), .Y(n241) );
  AND2X1 U696 ( .A(n1323), .B(n1326), .Y(n242) );
  INVX1 U697 ( .A(n242), .Y(n244) );
  AND2X1 U698 ( .A(n1326), .B(n1325), .Y(n260) );
  INVX1 U699 ( .A(n260), .Y(n262) );
  AND2X1 U700 ( .A(n87), .B(n772), .Y(n278) );
  INVX1 U701 ( .A(n278), .Y(n280) );
  AND2X1 U702 ( .A(n89), .B(n772), .Y(n296) );
  INVX1 U703 ( .A(n296), .Y(n298) );
  AND2X1 U704 ( .A(n93), .B(n772), .Y(n314) );
  INVX1 U705 ( .A(n314), .Y(n315) );
  AND2X1 U706 ( .A(n95), .B(n772), .Y(n317) );
  INVX1 U707 ( .A(n317), .Y(n333) );
  AND2X1 U708 ( .A(n112), .B(n772), .Y(n335) );
  INVX1 U709 ( .A(n335), .Y(n351) );
  AND2X1 U710 ( .A(n114), .B(n772), .Y(n353) );
  INVX1 U711 ( .A(n353), .Y(n354) );
  AND2X1 U712 ( .A(n130), .B(n773), .Y(n360) );
  INVX1 U713 ( .A(n360), .Y(n362) );
  AND2X1 U714 ( .A(n1488), .B(n663), .Y(n369) );
  INVX1 U715 ( .A(n369), .Y(n374) );
  AND2X1 U716 ( .A(n369), .B(n773), .Y(n634) );
  INVX1 U717 ( .A(n634), .Y(n635) );
  AND2X1 U718 ( .A(n1488), .B(n667), .Y(n636) );
  INVX1 U719 ( .A(n636), .Y(n637) );
  AND2X1 U720 ( .A(n636), .B(n773), .Y(n638) );
  INVX1 U721 ( .A(n638), .Y(n639) );
  AND2X1 U722 ( .A(n1488), .B(n1537), .Y(n640) );
  INVX1 U723 ( .A(n640), .Y(n641) );
  AND2X1 U724 ( .A(n640), .B(n773), .Y(n642) );
  INVX1 U725 ( .A(n642), .Y(n643) );
  AND2X1 U726 ( .A(n1488), .B(n1554), .Y(n644) );
  INVX1 U727 ( .A(n644), .Y(n645) );
  AND2X1 U728 ( .A(n644), .B(n773), .Y(n646) );
  INVX1 U729 ( .A(n646), .Y(n647) );
  AND2X1 U730 ( .A(n131), .B(n773), .Y(n648) );
  INVX1 U731 ( .A(n648), .Y(n649) );
  AND2X1 U732 ( .A(n133), .B(n773), .Y(n650) );
  INVX1 U733 ( .A(n650), .Y(n651) );
  AND2X1 U734 ( .A(n1537), .B(n1555), .Y(n652) );
  INVX1 U735 ( .A(n652), .Y(n653) );
  AND2X1 U736 ( .A(n652), .B(n773), .Y(n654) );
  INVX1 U737 ( .A(n654), .Y(n655) );
  AND2X1 U738 ( .A(n1555), .B(n1554), .Y(n656) );
  INVX1 U739 ( .A(n656), .Y(n657) );
  AND2X1 U740 ( .A(n772), .B(n656), .Y(n658) );
  INVX1 U741 ( .A(n658), .Y(n659) );
  OR2X1 U742 ( .A(n778), .B(n789), .Y(n660) );
  INVX1 U743 ( .A(n660), .Y(n661) );
  OR2X1 U744 ( .A(N22), .B(N23), .Y(n662) );
  INVX1 U745 ( .A(n662), .Y(n663) );
  OR2X1 U746 ( .A(n688), .B(n789), .Y(n664) );
  INVX1 U747 ( .A(n664), .Y(n665) );
  OR2X1 U748 ( .A(n799), .B(N23), .Y(n666) );
  INVX1 U749 ( .A(n666), .Y(n667) );
  OR2X1 U750 ( .A(n794), .B(n797), .Y(n668) );
  INVX1 U751 ( .A(n668), .Y(n669) );
  OR2X1 U752 ( .A(N24), .B(N25), .Y(n670) );
  INVX1 U753 ( .A(n670), .Y(n671) );
  OR2X1 U754 ( .A(n795), .B(n797), .Y(n672) );
  INVX1 U755 ( .A(n672), .Y(n673) );
  OR2X1 U756 ( .A(n800), .B(N25), .Y(n674) );
  INVX1 U757 ( .A(n674), .Y(n675) );
  MUX2X1 U758 ( .B(n1033), .A(n1034), .S(n676), .Y(n1042) );
  MUX2X1 U759 ( .B(\mem<201> ), .A(\mem<200> ), .S(n688), .Y(n992) );
  INVX1 U760 ( .A(n685), .Y(n677) );
  MUX2X1 U761 ( .B(n1019), .A(n1020), .S(n676), .Y(n1028) );
  MUX2X1 U762 ( .B(n995), .A(n996), .S(n796), .Y(n997) );
  MUX2X1 U763 ( .B(n993), .A(n994), .S(n697), .Y(n995) );
  INVX2 U764 ( .A(n790), .Y(n788) );
  INVX1 U765 ( .A(n787), .Y(n697) );
  MUX2X1 U766 ( .B(n999), .A(n1000), .S(n684), .Y(n1004) );
  INVX1 U767 ( .A(n787), .Y(n684) );
  MUX2X1 U768 ( .B(\mem<153> ), .A(\mem<152> ), .S(n678), .Y(n944) );
  INVX1 U769 ( .A(n774), .Y(n678) );
  MUX2X1 U770 ( .B(\mem<65> ), .A(\mem<64> ), .S(n782), .Y(n862) );
  MUX2X1 U771 ( .B(n1043), .A(n1044), .S(n799), .Y(n1045) );
  MUX2X1 U772 ( .B(n1031), .A(n1032), .S(n691), .Y(n1033) );
  INVX2 U773 ( .A(n790), .Y(n789) );
  MUX2X1 U774 ( .B(\mem<212> ), .A(\mem<213> ), .S(n686), .Y(n1002) );
  INVX8 U775 ( .A(n782), .Y(n779) );
  MUX2X1 U776 ( .B(n896), .A(n897), .S(n679), .Y(n901) );
  INVX1 U777 ( .A(n782), .Y(n680) );
  INVX1 U778 ( .A(write), .Y(n1051) );
  INVX1 U779 ( .A(n678), .Y(n681) );
  MUX2X1 U780 ( .B(n939), .A(n940), .S(n684), .Y(n941) );
  MUX2X1 U781 ( .B(n943), .A(n944), .S(n790), .Y(n948) );
  MUX2X1 U782 ( .B(\mem<19> ), .A(\mem<18> ), .S(n698), .Y(n815) );
  BUFX2 U783 ( .A(n774), .Y(n685) );
  INVX1 U784 ( .A(n698), .Y(n686) );
  MUX2X1 U785 ( .B(\mem<35> ), .A(\mem<34> ), .S(n677), .Y(n830) );
  BUFX4 U786 ( .A(n694), .Y(n687) );
  MUX2X1 U787 ( .B(n815), .A(n816), .S(n791), .Y(n819) );
  INVX1 U788 ( .A(n689), .Y(n688) );
  INVX1 U789 ( .A(n678), .Y(n689) );
  MUX2X1 U790 ( .B(n801), .A(n802), .S(n791), .Y(n806) );
  MUX2X1 U791 ( .B(\mem<197> ), .A(\mem<196> ), .S(n698), .Y(n988) );
  MUX2X1 U792 ( .B(\mem<105> ), .A(\mem<104> ), .S(n696), .Y(n897) );
  INVX1 U793 ( .A(n784), .Y(n691) );
  INVX4 U794 ( .A(N19), .Y(n791) );
  INVX4 U795 ( .A(N19), .Y(n790) );
  INVX1 U796 ( .A(n774), .Y(n692) );
  INVX1 U797 ( .A(n695), .Y(n693) );
  MUX2X1 U798 ( .B(n1009), .A(n1010), .S(n795), .Y(n1011) );
  MUX2X1 U799 ( .B(\mem<157> ), .A(\mem<156> ), .S(n687), .Y(n946) );
  INVX1 U800 ( .A(n692), .Y(n695) );
  INVX1 U801 ( .A(n695), .Y(n696) );
  MUX2X1 U802 ( .B(n985), .A(n986), .S(n790), .Y(n990) );
  MUX2X1 U803 ( .B(n989), .A(n990), .S(n795), .Y(n998) );
  INVX2 U804 ( .A(n795), .Y(n792) );
  MUX2X1 U805 ( .B(n1011), .A(n1012), .S(n798), .Y(n1013) );
  INVX1 U806 ( .A(n798), .Y(n797) );
  MUX2X1 U807 ( .B(\mem<51> ), .A(\mem<50> ), .S(n698), .Y(n844) );
  MUX2X1 U808 ( .B(n945), .A(n946), .S(n697), .Y(n947) );
  MUX2X1 U809 ( .B(\mem<37> ), .A(\mem<36> ), .S(n782), .Y(n833) );
  INVX1 U810 ( .A(n692), .Y(n699) );
  MUX2X1 U811 ( .B(\mem<33> ), .A(\mem<32> ), .S(n693), .Y(n831) );
  MUX2X1 U812 ( .B(n834), .A(n835), .S(n796), .Y(n843) );
  INVX2 U813 ( .A(n796), .Y(n794) );
  MUX2X1 U814 ( .B(n902), .A(n903), .S(n798), .Y(n919) );
  INVX1 U815 ( .A(N21), .Y(n700) );
  MUX2X1 U816 ( .B(n879), .A(n878), .S(N20), .Y(n887) );
  MUX2X1 U817 ( .B(n703), .A(n702), .S(n775), .Y(n701) );
  MUX2X1 U818 ( .B(n908), .A(n909), .S(n796), .Y(n917) );
  INVX2 U819 ( .A(n796), .Y(n793) );
  MUX2X1 U820 ( .B(n919), .A(n918), .S(N22), .Y(n920) );
  INVX1 U821 ( .A(N22), .Y(n799) );
  MUX2X1 U822 ( .B(\mem<155> ), .A(\mem<154> ), .S(n687), .Y(n943) );
  MUX2X1 U823 ( .B(n951), .A(n952), .S(n799), .Y(n984) );
  MUX2X1 U824 ( .B(\mem<69> ), .A(\mem<68> ), .S(n698), .Y(n864) );
  MUX2X1 U825 ( .B(n950), .A(n949), .S(N21), .Y(n951) );
  INVX1 U826 ( .A(N21), .Y(n798) );
  MUX2X1 U827 ( .B(n1047), .A(n6), .S(n800), .Y(n1048) );
  MUX2X1 U828 ( .B(n859), .A(n860), .S(n704), .Y(n922) );
  MUX2X1 U829 ( .B(n922), .A(n7), .S(N24), .Y(n1049) );
  INVX1 U830 ( .A(N24), .Y(n800) );
  INVX1 U831 ( .A(N23), .Y(n704) );
  INVX1 U832 ( .A(n785), .Y(n705) );
  MUX2X1 U833 ( .B(n888), .A(n889), .S(n799), .Y(n921) );
  INVX8 U834 ( .A(n775), .Y(n774) );
  INVX8 U835 ( .A(n782), .Y(n776) );
  INVX8 U836 ( .A(n694), .Y(n778) );
  INVX8 U837 ( .A(n782), .Y(n780) );
  INVX8 U838 ( .A(n774), .Y(n782) );
  INVX8 U839 ( .A(n774), .Y(n783) );
  INVX8 U840 ( .A(n791), .Y(n784) );
  INVX8 U841 ( .A(n791), .Y(n785) );
  INVX8 U842 ( .A(n791), .Y(n786) );
  INVX8 U843 ( .A(n790), .Y(n787) );
  INVX4 U844 ( .A(N20), .Y(n795) );
  INVX4 U845 ( .A(N20), .Y(n796) );
  MUX2X1 U846 ( .B(\mem<0> ), .A(\mem<1> ), .S(n776), .Y(n802) );
  MUX2X1 U847 ( .B(\mem<2> ), .A(\mem<3> ), .S(n778), .Y(n801) );
  MUX2X1 U848 ( .B(\mem<4> ), .A(\mem<5> ), .S(n699), .Y(n804) );
  MUX2X1 U849 ( .B(\mem<6> ), .A(\mem<7> ), .S(n781), .Y(n803) );
  MUX2X1 U850 ( .B(n804), .A(n803), .S(n784), .Y(n805) );
  MUX2X1 U851 ( .B(n806), .A(n805), .S(n792), .Y(n814) );
  MUX2X1 U852 ( .B(\mem<8> ), .A(\mem<9> ), .S(n781), .Y(n808) );
  MUX2X1 U853 ( .B(\mem<10> ), .A(\mem<11> ), .S(n777), .Y(n807) );
  MUX2X1 U854 ( .B(n808), .A(n807), .S(n784), .Y(n812) );
  MUX2X1 U855 ( .B(\mem<12> ), .A(\mem<13> ), .S(n778), .Y(n810) );
  MUX2X1 U856 ( .B(\mem<14> ), .A(\mem<15> ), .S(n778), .Y(n809) );
  MUX2X1 U857 ( .B(n810), .A(n809), .S(n784), .Y(n811) );
  MUX2X1 U858 ( .B(n812), .A(n811), .S(n794), .Y(n813) );
  MUX2X1 U859 ( .B(n814), .A(n813), .S(N21), .Y(n829) );
  MUX2X1 U860 ( .B(\mem<16> ), .A(\mem<17> ), .S(n777), .Y(n816) );
  MUX2X1 U861 ( .B(\mem<20> ), .A(\mem<21> ), .S(n781), .Y(n818) );
  MUX2X1 U862 ( .B(\mem<22> ), .A(\mem<23> ), .S(n682), .Y(n817) );
  MUX2X1 U863 ( .B(n819), .A(n2), .S(n794), .Y(n827) );
  MUX2X1 U864 ( .B(\mem<24> ), .A(\mem<25> ), .S(n781), .Y(n821) );
  MUX2X1 U865 ( .B(\mem<26> ), .A(\mem<27> ), .S(n777), .Y(n820) );
  MUX2X1 U866 ( .B(n821), .A(n820), .S(n784), .Y(n825) );
  MUX2X1 U867 ( .B(\mem<28> ), .A(\mem<29> ), .S(n777), .Y(n823) );
  MUX2X1 U868 ( .B(\mem<30> ), .A(\mem<31> ), .S(n777), .Y(n822) );
  MUX2X1 U869 ( .B(n823), .A(n822), .S(n784), .Y(n824) );
  MUX2X1 U870 ( .B(n825), .A(n824), .S(n794), .Y(n826) );
  MUX2X1 U871 ( .B(n827), .A(n826), .S(N21), .Y(n828) );
  MUX2X1 U872 ( .B(n829), .A(n828), .S(N22), .Y(n860) );
  MUX2X1 U873 ( .B(n831), .A(n830), .S(n784), .Y(n835) );
  MUX2X1 U874 ( .B(\mem<38> ), .A(\mem<39> ), .S(n680), .Y(n832) );
  MUX2X1 U875 ( .B(n833), .A(n832), .S(n784), .Y(n834) );
  MUX2X1 U876 ( .B(\mem<40> ), .A(\mem<41> ), .S(n780), .Y(n837) );
  MUX2X1 U877 ( .B(\mem<42> ), .A(\mem<43> ), .S(n777), .Y(n836) );
  MUX2X1 U878 ( .B(n837), .A(n836), .S(n784), .Y(n841) );
  MUX2X1 U879 ( .B(\mem<44> ), .A(\mem<45> ), .S(n780), .Y(n839) );
  MUX2X1 U880 ( .B(\mem<46> ), .A(\mem<47> ), .S(n780), .Y(n838) );
  MUX2X1 U881 ( .B(n839), .A(n838), .S(n784), .Y(n840) );
  MUX2X1 U882 ( .B(n841), .A(n840), .S(n794), .Y(n842) );
  MUX2X1 U883 ( .B(n843), .A(n842), .S(N21), .Y(n858) );
  MUX2X1 U884 ( .B(\mem<48> ), .A(\mem<49> ), .S(n780), .Y(n845) );
  MUX2X1 U885 ( .B(n845), .A(n844), .S(n784), .Y(n849) );
  MUX2X1 U886 ( .B(\mem<52> ), .A(\mem<53> ), .S(n780), .Y(n847) );
  MUX2X1 U887 ( .B(\mem<54> ), .A(\mem<55> ), .S(n780), .Y(n846) );
  MUX2X1 U888 ( .B(n847), .A(n846), .S(n785), .Y(n848) );
  MUX2X1 U889 ( .B(n849), .A(n848), .S(n794), .Y(n857) );
  MUX2X1 U890 ( .B(\mem<56> ), .A(\mem<57> ), .S(n777), .Y(n851) );
  MUX2X1 U891 ( .B(\mem<58> ), .A(\mem<59> ), .S(n780), .Y(n850) );
  MUX2X1 U892 ( .B(n851), .A(n850), .S(n785), .Y(n855) );
  MUX2X1 U893 ( .B(\mem<60> ), .A(\mem<61> ), .S(n780), .Y(n853) );
  MUX2X1 U894 ( .B(\mem<62> ), .A(\mem<63> ), .S(n781), .Y(n852) );
  MUX2X1 U895 ( .B(n853), .A(n852), .S(n785), .Y(n854) );
  MUX2X1 U896 ( .B(n855), .A(n854), .S(n794), .Y(n856) );
  MUX2X1 U897 ( .B(n858), .A(n5), .S(N22), .Y(n859) );
  MUX2X1 U898 ( .B(\mem<66> ), .A(\mem<67> ), .S(n777), .Y(n861) );
  MUX2X1 U899 ( .B(n862), .A(n861), .S(n785), .Y(n865) );
  MUX2X1 U900 ( .B(\mem<70> ), .A(\mem<71> ), .S(n1), .Y(n863) );
  MUX2X1 U901 ( .B(n865), .A(n8), .S(n794), .Y(n873) );
  MUX2X1 U902 ( .B(\mem<72> ), .A(\mem<73> ), .S(n781), .Y(n867) );
  MUX2X1 U903 ( .B(\mem<74> ), .A(\mem<75> ), .S(n778), .Y(n866) );
  MUX2X1 U904 ( .B(n867), .A(n866), .S(n785), .Y(n871) );
  MUX2X1 U905 ( .B(\mem<76> ), .A(\mem<77> ), .S(n683), .Y(n869) );
  MUX2X1 U906 ( .B(\mem<78> ), .A(\mem<79> ), .S(n779), .Y(n868) );
  MUX2X1 U907 ( .B(n869), .A(n868), .S(n785), .Y(n870) );
  MUX2X1 U908 ( .B(n871), .A(n870), .S(n793), .Y(n872) );
  MUX2X1 U909 ( .B(n873), .A(n872), .S(N21), .Y(n889) );
  MUX2X1 U910 ( .B(\mem<80> ), .A(\mem<81> ), .S(n699), .Y(n875) );
  MUX2X1 U911 ( .B(\mem<82> ), .A(\mem<83> ), .S(n681), .Y(n874) );
  MUX2X1 U912 ( .B(n875), .A(n874), .S(n785), .Y(n879) );
  MUX2X1 U913 ( .B(\mem<84> ), .A(\mem<85> ), .S(n690), .Y(n877) );
  MUX2X1 U914 ( .B(\mem<86> ), .A(\mem<87> ), .S(n778), .Y(n876) );
  MUX2X1 U915 ( .B(n877), .A(n876), .S(n785), .Y(n878) );
  MUX2X1 U916 ( .B(\mem<88> ), .A(\mem<89> ), .S(n781), .Y(n881) );
  MUX2X1 U917 ( .B(\mem<90> ), .A(\mem<91> ), .S(n781), .Y(n880) );
  MUX2X1 U918 ( .B(n881), .A(n880), .S(n785), .Y(n885) );
  MUX2X1 U919 ( .B(\mem<92> ), .A(\mem<93> ), .S(n781), .Y(n883) );
  MUX2X1 U920 ( .B(\mem<94> ), .A(\mem<95> ), .S(n781), .Y(n882) );
  MUX2X1 U921 ( .B(n883), .A(n882), .S(n785), .Y(n884) );
  MUX2X1 U922 ( .B(n885), .A(n884), .S(n793), .Y(n886) );
  MUX2X1 U923 ( .B(n887), .A(n886), .S(N21), .Y(n888) );
  MUX2X1 U924 ( .B(\mem<96> ), .A(\mem<97> ), .S(n689), .Y(n891) );
  MUX2X1 U925 ( .B(\mem<98> ), .A(\mem<99> ), .S(n690), .Y(n890) );
  MUX2X1 U926 ( .B(n891), .A(n890), .S(n785), .Y(n895) );
  MUX2X1 U927 ( .B(\mem<100> ), .A(\mem<101> ), .S(n777), .Y(n893) );
  MUX2X1 U928 ( .B(\mem<102> ), .A(\mem<103> ), .S(n781), .Y(n892) );
  MUX2X1 U929 ( .B(n893), .A(n892), .S(n786), .Y(n894) );
  MUX2X1 U930 ( .B(n895), .A(n894), .S(n793), .Y(n903) );
  MUX2X1 U931 ( .B(\mem<106> ), .A(\mem<107> ), .S(n780), .Y(n896) );
  MUX2X1 U932 ( .B(\mem<108> ), .A(\mem<109> ), .S(n779), .Y(n899) );
  MUX2X1 U933 ( .B(\mem<110> ), .A(\mem<111> ), .S(n781), .Y(n898) );
  MUX2X1 U934 ( .B(n899), .A(n898), .S(n786), .Y(n900) );
  MUX2X1 U935 ( .B(n901), .A(n900), .S(n793), .Y(n902) );
  MUX2X1 U936 ( .B(\mem<114> ), .A(\mem<115> ), .S(n776), .Y(n904) );
  MUX2X1 U937 ( .B(n905), .A(n904), .S(n786), .Y(n909) );
  MUX2X1 U938 ( .B(\mem<116> ), .A(\mem<117> ), .S(n779), .Y(n907) );
  MUX2X1 U939 ( .B(\mem<118> ), .A(\mem<119> ), .S(n777), .Y(n906) );
  MUX2X1 U940 ( .B(n907), .A(n906), .S(n786), .Y(n908) );
  MUX2X1 U941 ( .B(\mem<120> ), .A(\mem<121> ), .S(n680), .Y(n911) );
  MUX2X1 U942 ( .B(\mem<122> ), .A(\mem<123> ), .S(n681), .Y(n910) );
  MUX2X1 U943 ( .B(n911), .A(n910), .S(n786), .Y(n915) );
  MUX2X1 U944 ( .B(\mem<124> ), .A(\mem<125> ), .S(n776), .Y(n913) );
  MUX2X1 U945 ( .B(\mem<126> ), .A(\mem<127> ), .S(n689), .Y(n912) );
  MUX2X1 U946 ( .B(n913), .A(n912), .S(n786), .Y(n914) );
  MUX2X1 U947 ( .B(n915), .A(n914), .S(n793), .Y(n916) );
  MUX2X1 U948 ( .B(n917), .A(n916), .S(N21), .Y(n918) );
  MUX2X1 U949 ( .B(\mem<128> ), .A(\mem<129> ), .S(n686), .Y(n924) );
  MUX2X1 U950 ( .B(\mem<130> ), .A(\mem<131> ), .S(n779), .Y(n923) );
  MUX2X1 U951 ( .B(n924), .A(n923), .S(n786), .Y(n928) );
  MUX2X1 U952 ( .B(\mem<132> ), .A(\mem<133> ), .S(n681), .Y(n926) );
  MUX2X1 U953 ( .B(\mem<134> ), .A(\mem<135> ), .S(n690), .Y(n925) );
  MUX2X1 U954 ( .B(n926), .A(n925), .S(n786), .Y(n927) );
  MUX2X1 U955 ( .B(n928), .A(n927), .S(n793), .Y(n936) );
  MUX2X1 U956 ( .B(\mem<136> ), .A(\mem<137> ), .S(n778), .Y(n930) );
  MUX2X1 U957 ( .B(\mem<138> ), .A(\mem<139> ), .S(n780), .Y(n929) );
  MUX2X1 U958 ( .B(n930), .A(n929), .S(n786), .Y(n934) );
  MUX2X1 U959 ( .B(\mem<140> ), .A(\mem<141> ), .S(n778), .Y(n932) );
  MUX2X1 U960 ( .B(\mem<142> ), .A(\mem<143> ), .S(n778), .Y(n931) );
  MUX2X1 U961 ( .B(n932), .A(n931), .S(n786), .Y(n933) );
  MUX2X1 U962 ( .B(n934), .A(n933), .S(n793), .Y(n935) );
  MUX2X1 U963 ( .B(n936), .A(n935), .S(N21), .Y(n952) );
  MUX2X1 U964 ( .B(\mem<144> ), .A(\mem<145> ), .S(n685), .Y(n938) );
  MUX2X1 U965 ( .B(\mem<146> ), .A(\mem<147> ), .S(n685), .Y(n937) );
  MUX2X1 U966 ( .B(n938), .A(n937), .S(n787), .Y(n942) );
  MUX2X1 U967 ( .B(\mem<148> ), .A(\mem<149> ), .S(n778), .Y(n940) );
  MUX2X1 U968 ( .B(\mem<150> ), .A(\mem<151> ), .S(n779), .Y(n939) );
  MUX2X1 U969 ( .B(n942), .A(n941), .S(n793), .Y(n950) );
  MUX2X1 U970 ( .B(\mem<158> ), .A(\mem<159> ), .S(n777), .Y(n945) );
  MUX2X1 U971 ( .B(n948), .A(n947), .S(n793), .Y(n949) );
  MUX2X1 U972 ( .B(\mem<160> ), .A(\mem<161> ), .S(n781), .Y(n954) );
  MUX2X1 U973 ( .B(\mem<162> ), .A(\mem<163> ), .S(n695), .Y(n953) );
  MUX2X1 U974 ( .B(n954), .A(n953), .S(n787), .Y(n958) );
  MUX2X1 U975 ( .B(\mem<164> ), .A(\mem<165> ), .S(n685), .Y(n956) );
  MUX2X1 U976 ( .B(\mem<166> ), .A(\mem<167> ), .S(n777), .Y(n955) );
  MUX2X1 U977 ( .B(n956), .A(n955), .S(n787), .Y(n957) );
  MUX2X1 U978 ( .B(n958), .A(n957), .S(n792), .Y(n966) );
  MUX2X1 U979 ( .B(\mem<168> ), .A(\mem<169> ), .S(n778), .Y(n960) );
  MUX2X1 U980 ( .B(\mem<170> ), .A(\mem<171> ), .S(n695), .Y(n959) );
  MUX2X1 U981 ( .B(n960), .A(n959), .S(n787), .Y(n964) );
  MUX2X1 U982 ( .B(\mem<172> ), .A(\mem<173> ), .S(n781), .Y(n962) );
  MUX2X1 U983 ( .B(\mem<174> ), .A(\mem<175> ), .S(n777), .Y(n961) );
  MUX2X1 U984 ( .B(n962), .A(n961), .S(n787), .Y(n963) );
  MUX2X1 U985 ( .B(n964), .A(n963), .S(n792), .Y(n965) );
  MUX2X1 U986 ( .B(n966), .A(n965), .S(N21), .Y(n982) );
  MUX2X1 U987 ( .B(\mem<176> ), .A(\mem<177> ), .S(n778), .Y(n968) );
  MUX2X1 U988 ( .B(\mem<178> ), .A(\mem<179> ), .S(n778), .Y(n967) );
  MUX2X1 U989 ( .B(n968), .A(n967), .S(n787), .Y(n972) );
  MUX2X1 U990 ( .B(\mem<180> ), .A(\mem<181> ), .S(n699), .Y(n970) );
  MUX2X1 U991 ( .B(\mem<182> ), .A(\mem<183> ), .S(n777), .Y(n969) );
  MUX2X1 U992 ( .B(n970), .A(n969), .S(n787), .Y(n971) );
  MUX2X1 U993 ( .B(n972), .A(n971), .S(n792), .Y(n980) );
  MUX2X1 U994 ( .B(\mem<184> ), .A(\mem<185> ), .S(n683), .Y(n974) );
  MUX2X1 U995 ( .B(\mem<186> ), .A(\mem<187> ), .S(n777), .Y(n973) );
  MUX2X1 U996 ( .B(n974), .A(n973), .S(n787), .Y(n978) );
  MUX2X1 U997 ( .B(\mem<188> ), .A(\mem<189> ), .S(n777), .Y(n976) );
  MUX2X1 U998 ( .B(\mem<190> ), .A(\mem<191> ), .S(n777), .Y(n975) );
  MUX2X1 U999 ( .B(n976), .A(n975), .S(n787), .Y(n977) );
  MUX2X1 U1000 ( .B(n978), .A(n977), .S(n792), .Y(n979) );
  MUX2X1 U1001 ( .B(n980), .A(n979), .S(N21), .Y(n981) );
  MUX2X1 U1002 ( .B(n982), .A(n981), .S(N22), .Y(n983) );
  MUX2X1 U1003 ( .B(\mem<192> ), .A(\mem<193> ), .S(n777), .Y(n986) );
  MUX2X1 U1004 ( .B(\mem<194> ), .A(\mem<195> ), .S(n779), .Y(n985) );
  MUX2X1 U1005 ( .B(\mem<198> ), .A(\mem<199> ), .S(n779), .Y(n987) );
  MUX2X1 U1006 ( .B(n988), .A(n987), .S(n788), .Y(n989) );
  MUX2X1 U1007 ( .B(\mem<202> ), .A(\mem<203> ), .S(n779), .Y(n991) );
  MUX2X1 U1008 ( .B(n992), .A(n991), .S(n788), .Y(n996) );
  MUX2X1 U1009 ( .B(\mem<204> ), .A(\mem<205> ), .S(n683), .Y(n994) );
  MUX2X1 U1010 ( .B(\mem<206> ), .A(\mem<207> ), .S(n777), .Y(n993) );
  MUX2X1 U1011 ( .B(n998), .A(n997), .S(n797), .Y(n1014) );
  MUX2X1 U1012 ( .B(\mem<208> ), .A(\mem<209> ), .S(n781), .Y(n1000) );
  MUX2X1 U1013 ( .B(\mem<210> ), .A(\mem<211> ), .S(n683), .Y(n999) );
  MUX2X1 U1014 ( .B(\mem<214> ), .A(\mem<215> ), .S(n781), .Y(n1001) );
  MUX2X1 U1015 ( .B(n1002), .A(n1001), .S(n788), .Y(n1003) );
  MUX2X1 U1016 ( .B(n1004), .A(n1003), .S(n792), .Y(n1012) );
  MUX2X1 U1017 ( .B(\mem<216> ), .A(\mem<217> ), .S(n690), .Y(n1006) );
  MUX2X1 U1018 ( .B(\mem<218> ), .A(\mem<219> ), .S(n781), .Y(n1005) );
  MUX2X1 U1019 ( .B(n1006), .A(n1005), .S(n788), .Y(n1010) );
  MUX2X1 U1020 ( .B(\mem<220> ), .A(\mem<221> ), .S(n779), .Y(n1008) );
  MUX2X1 U1021 ( .B(\mem<222> ), .A(\mem<223> ), .S(n781), .Y(n1007) );
  MUX2X1 U1022 ( .B(n1008), .A(n1007), .S(n788), .Y(n1009) );
  MUX2X1 U1023 ( .B(n1014), .A(n1013), .S(N22), .Y(n1046) );
  MUX2X1 U1024 ( .B(\mem<224> ), .A(\mem<225> ), .S(n777), .Y(n1016) );
  MUX2X1 U1025 ( .B(\mem<226> ), .A(\mem<227> ), .S(n781), .Y(n1015) );
  MUX2X1 U1026 ( .B(n1016), .A(n1015), .S(n788), .Y(n1020) );
  MUX2X1 U1027 ( .B(\mem<228> ), .A(\mem<229> ), .S(n781), .Y(n1018) );
  MUX2X1 U1028 ( .B(\mem<230> ), .A(\mem<231> ), .S(n777), .Y(n1017) );
  MUX2X1 U1029 ( .B(n1018), .A(n1017), .S(n788), .Y(n1019) );
  MUX2X1 U1030 ( .B(\mem<232> ), .A(\mem<233> ), .S(n781), .Y(n1022) );
  MUX2X1 U1031 ( .B(\mem<234> ), .A(\mem<235> ), .S(n776), .Y(n1021) );
  MUX2X1 U1032 ( .B(n1022), .A(n1021), .S(n788), .Y(n1026) );
  MUX2X1 U1033 ( .B(\mem<236> ), .A(\mem<237> ), .S(n776), .Y(n1024) );
  MUX2X1 U1034 ( .B(\mem<238> ), .A(\mem<239> ), .S(n776), .Y(n1023) );
  MUX2X1 U1035 ( .B(n1024), .A(n1023), .S(n788), .Y(n1025) );
  MUX2X1 U1036 ( .B(n1026), .A(n1025), .S(n792), .Y(n1027) );
  MUX2X1 U1037 ( .B(n1028), .A(n1027), .S(n797), .Y(n1044) );
  MUX2X1 U1038 ( .B(\mem<240> ), .A(\mem<241> ), .S(n776), .Y(n1030) );
  MUX2X1 U1039 ( .B(\mem<242> ), .A(\mem<243> ), .S(n776), .Y(n1029) );
  MUX2X1 U1040 ( .B(n1030), .A(n1029), .S(n789), .Y(n1034) );
  MUX2X1 U1041 ( .B(\mem<244> ), .A(\mem<245> ), .S(n776), .Y(n1032) );
  MUX2X1 U1042 ( .B(\mem<246> ), .A(\mem<247> ), .S(n776), .Y(n1031) );
  MUX2X1 U1043 ( .B(\mem<248> ), .A(\mem<249> ), .S(n776), .Y(n1036) );
  MUX2X1 U1044 ( .B(\mem<250> ), .A(\mem<251> ), .S(n776), .Y(n1035) );
  MUX2X1 U1045 ( .B(n1036), .A(n1035), .S(n789), .Y(n1040) );
  MUX2X1 U1046 ( .B(\mem<252> ), .A(\mem<253> ), .S(n776), .Y(n1038) );
  MUX2X1 U1047 ( .B(\mem<254> ), .A(\mem<255> ), .S(n776), .Y(n1037) );
  MUX2X1 U1048 ( .B(n1038), .A(n1037), .S(n789), .Y(n1039) );
  MUX2X1 U1049 ( .B(n1040), .A(n1039), .S(n792), .Y(n1041) );
  MUX2X1 U1050 ( .B(n1042), .A(n1041), .S(n797), .Y(n1043) );
  MUX2X1 U1051 ( .B(n1046), .A(n1045), .S(N23), .Y(n1047) );
  MUX2X1 U1052 ( .B(n1049), .A(n1048), .S(N25), .Y(n1050) );
  AND2X2 U1053 ( .A(n1050), .B(n24), .Y(data_out) );
endmodule


module final_memory_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1046, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n373, n374, n375, n376, n377, n378, n380,
         n382, n383, n384, n385, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n584, n585, n586, n587,
         n588, n589, n590, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n50, n150, n189, n289, n348, n372, n379, n381, n386, n387,
         n401, n402, n409, n421, n422, n434, n435, n447, n448, n460, n461,
         n473, n474, n486, n487, n507, n508, n522, n523, n537, n538, n552,
         n553, n567, n568, n582, n583, n591, n592, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n870), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n869), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n868), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n867), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n866), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n865), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n864), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n863), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n862), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n861), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n860), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n859), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n858), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n857), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n856), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n855), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n854), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n853), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n852), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n851), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n850), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n849), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n848), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n847), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n846), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n845), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n844), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n843), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n842), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n841), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n840), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n839), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n838), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n837), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n836), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n835), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n834), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n833), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n832), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n831), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n830), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n829), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n828), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n827), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n826), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n825), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n824), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n823), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n822), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n821), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n820), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n819), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n818), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n817), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n816), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n815), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n814), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n813), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n812), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n811), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n810), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n809), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n808), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n807), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n806), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n805), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n804), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n803), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n802), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n801), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n800), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n799), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n798), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n797), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n796), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n795), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n794), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n793), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n792), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n791), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n790), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n789), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n788), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n787), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n786), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n785), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n784), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n783), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n782), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n781), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n780), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n779), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n778), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n777), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n776), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n775), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n774), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n773), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n772), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n771), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n770), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n769), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n768), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n767), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n766), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n765), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n764), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n763), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n762), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n761), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n760), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n759), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n758), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n757), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n756), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n755), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n754), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n753), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n752), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n751), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n750), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n749), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n748), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n747), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n746), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n745), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n744), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n743), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n742), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n741), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n740), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n739), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n738), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n737), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n736), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n735), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n734), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n733), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n732), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n731), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n730), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n729), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n728), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n727), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n726), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n725), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n724), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n723), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n722), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n721), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n720), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n719), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n718), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n717), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n716), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n715), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n714), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n713), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n712), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n711), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n710), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n709), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n708), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n707), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n706), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n705), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n704), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n703), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n702), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n701), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n700), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n699), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n698), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n697), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n696), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n695), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n694), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n693), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n692), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n691), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n690), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n689), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n688), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n687), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n686), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n685), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n684), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n683), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n682), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n681), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n680), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n679), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n678), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n677), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n676), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n675), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n674), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n673), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n672), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n671), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n670), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n669), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n668), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n667), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n666), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n665), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n664), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n663), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n662), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n661), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n660), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n659), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n658), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n657), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n656), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n655), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n654), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n653), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n652), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n651), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n650), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n649), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n648), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n647), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n646), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n645), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n644), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n643), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n642), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n641), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n640), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n639), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n638), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n637), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n636), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n635), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n634), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n633), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n632), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n631), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n630), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n629), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n628), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n627), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n626), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n625), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n624), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n623), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n622), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n621), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n620), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n619), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n618), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n617), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n616), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n615), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n614), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n613), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n612), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n611), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n610), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n609), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n608), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n607), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U4 ( .A(wr1), .B(n1013), .Y(n48) );
  AND2X2 U9 ( .A(n413), .B(n414), .Y(n412) );
  AND2X2 U10 ( .A(n418), .B(n419), .Y(n417) );
  AND2X2 U11 ( .A(n426), .B(n427), .Y(n425) );
  AND2X2 U12 ( .A(n431), .B(n432), .Y(n430) );
  AND2X2 U13 ( .A(n439), .B(n440), .Y(n438) );
  AND2X2 U14 ( .A(n444), .B(n445), .Y(n443) );
  AND2X2 U15 ( .A(n452), .B(n453), .Y(n451) );
  AND2X2 U16 ( .A(n457), .B(n458), .Y(n456) );
  AND2X2 U17 ( .A(n465), .B(n466), .Y(n464) );
  AND2X2 U18 ( .A(n470), .B(n471), .Y(n469) );
  AND2X2 U19 ( .A(n478), .B(n479), .Y(n477) );
  AND2X2 U20 ( .A(n483), .B(n484), .Y(n482) );
  AND2X2 U21 ( .A(n491), .B(n492), .Y(n490) );
  AND2X2 U22 ( .A(n496), .B(n497), .Y(n495) );
  AND2X2 U30 ( .A(n588), .B(n1026), .Y(n248) );
  AND2X2 U31 ( .A(n589), .B(n1026), .Y(n91) );
  AND2X2 U32 ( .A(n588), .B(\addr_1c<0> ), .Y(n228) );
  AND2X2 U33 ( .A(n589), .B(\addr_1c<0> ), .Y(n71) );
  AND2X2 U34 ( .A(n596), .B(n597), .Y(n595) );
  AND2X2 U45 ( .A(n603), .B(n604), .Y(n602) );
  NOR3X1 U94 ( .A(n1015), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1014), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n40), .Y(n607) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n40) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n41), .Y(n608) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n41) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n42), .Y(n609) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n42) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n43), .Y(n610) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n43) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n44), .Y(n611) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n44) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n45), .Y(n612) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n45) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n46), .Y(n613) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n46) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n47), .Y(n614) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n47) );
  NAND3X1 U112 ( .A(n48), .B(n49), .C(n964), .Y(n39) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n51), .Y(n615) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n51) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n52), .Y(n616) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n52) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n53), .Y(n617) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n53) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n54), .Y(n618) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n54) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n55), .Y(n619) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n55) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n56), .Y(n620) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n56) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n57), .Y(n621) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n57) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n58), .Y(n622) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n58) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n62), .Y(n623) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n62) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n63), .Y(n624) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n63) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n64), .Y(n625) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n64) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n65), .Y(n626) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n65) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n66), .Y(n627) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n66) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n67), .Y(n628) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n67) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n68), .Y(n629) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n68) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n69), .Y(n630) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n69) );
  NAND3X1 U146 ( .A(n70), .B(n48), .C(n71), .Y(n61) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n73), .Y(n631) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n73) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n74), .Y(n632) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n74) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n75), .Y(n633) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n75) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n76), .Y(n634) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n76) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n77), .Y(n635) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n77) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n78), .Y(n636) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n78) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n79), .Y(n637) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n79) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n80), .Y(n638) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n80) );
  NAND3X1 U163 ( .A(n973), .B(n48), .C(n81), .Y(n72) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n83), .Y(n639) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n83) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n84), .Y(n640) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n84) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n85), .Y(n641) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n85) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n86), .Y(n642) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n86) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n87), .Y(n643) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n87) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n88), .Y(n644) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n88) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n89), .Y(n645) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n89) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n90), .Y(n646) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n90) );
  NAND3X1 U180 ( .A(n70), .B(n48), .C(n91), .Y(n82) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n93), .Y(n647) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n93) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n94), .Y(n648) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n94) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n95), .Y(n649) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n95) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n96), .Y(n650) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n96) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n97), .Y(n651) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n97) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n98), .Y(n652) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n98) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n99), .Y(n653) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n99) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n100), .Y(n654) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n100) );
  NAND3X1 U197 ( .A(n973), .B(n48), .C(n101), .Y(n92) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n103), .Y(n655) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n103) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n104), .Y(n656) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n104) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n105), .Y(n657) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n105) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n106), .Y(n658) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n106) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n107), .Y(n659) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n107) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n108), .Y(n660) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n108) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n109), .Y(n661) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n109) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n110), .Y(n662) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n110) );
  NAND3X1 U214 ( .A(n71), .B(n48), .C(n111), .Y(n102) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n113), .Y(n663) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n113) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n114), .Y(n664) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n114) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n115), .Y(n665) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n115) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n116), .Y(n666) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n116) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n117), .Y(n667) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n117) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n118), .Y(n668) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n118) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n119), .Y(n669) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n119) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n120), .Y(n670) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n120) );
  NAND3X1 U231 ( .A(n973), .B(n48), .C(n121), .Y(n112) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n123), .Y(n671) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n123) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n124), .Y(n672) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n124) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n125), .Y(n673) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n125) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n126), .Y(n674) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n126) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n127), .Y(n675) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n127) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n128), .Y(n676) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n128) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n129), .Y(n677) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n129) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n130), .Y(n678) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n130) );
  NAND3X1 U248 ( .A(n91), .B(n48), .C(n111), .Y(n122) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n132), .Y(n679) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n132) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n133), .Y(n680) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n133) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n134), .Y(n681) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n134) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n135), .Y(n682) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n135) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n136), .Y(n683) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n136) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n137), .Y(n684) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n137) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n138), .Y(n685) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n138) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n139), .Y(n686) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n139) );
  NAND3X1 U265 ( .A(n973), .B(n48), .C(n140), .Y(n131) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n142), .Y(n687) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n142) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n143), .Y(n688) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n143) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n144), .Y(n689) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n144) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n145), .Y(n690) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n145) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n146), .Y(n691) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n146) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n147), .Y(n692) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n147) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n148), .Y(n693) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n148) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n149), .Y(n694) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n149) );
  NAND3X1 U282 ( .A(n71), .B(n48), .C(n969), .Y(n141) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n152), .Y(n695) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n152) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n153), .Y(n696) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n153) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n154), .Y(n697) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n154) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n155), .Y(n698) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n155) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n156), .Y(n699) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n156) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n157), .Y(n700) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n157) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n158), .Y(n701) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n158) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n159), .Y(n702) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n159) );
  NAND3X1 U299 ( .A(n973), .B(n48), .C(n160), .Y(n151) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n162), .Y(n703) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n162) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n163), .Y(n704) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n163) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n164), .Y(n705) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n164) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n165), .Y(n706) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n165) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n166), .Y(n707) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n166) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n167), .Y(n708) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n167) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n168), .Y(n709) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n168) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n169), .Y(n710) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n169) );
  NAND3X1 U316 ( .A(n91), .B(n48), .C(n969), .Y(n161) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n171), .Y(n711) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n171) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n172), .Y(n712) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n172) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n173), .Y(n713) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n173) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n174), .Y(n714) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n174) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n175), .Y(n715) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n175) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n176), .Y(n716) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n176) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n177), .Y(n717) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n177) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n178), .Y(n718) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n178) );
  NAND3X1 U333 ( .A(n973), .B(n48), .C(n179), .Y(n170) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n181), .Y(n719) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n181) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n182), .Y(n720) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n182) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n183), .Y(n721) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n183) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n184), .Y(n722) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n184) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n185), .Y(n723) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n185) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n186), .Y(n724) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n186) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n187), .Y(n725) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n187) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n188), .Y(n726) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n188) );
  NAND3X1 U350 ( .A(n71), .B(n48), .C(n967), .Y(n180) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n191), .Y(n727) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n191) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n192), .Y(n728) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n192) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n193), .Y(n729) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n193) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n194), .Y(n730) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n194) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n195), .Y(n731) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n195) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n196), .Y(n732) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n196) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n197), .Y(n733) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n197) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n198), .Y(n734) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n198) );
  NAND3X1 U367 ( .A(n973), .B(n48), .C(n199), .Y(n190) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n201), .Y(n735) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n201) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n202), .Y(n736) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n202) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n203), .Y(n737) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n203) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n204), .Y(n738) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n204) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n205), .Y(n739) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n205) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n206), .Y(n740) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n206) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n207), .Y(n741) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n207) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n208), .Y(n742) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n208) );
  NAND3X1 U384 ( .A(n91), .B(n48), .C(n967), .Y(n200) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n210), .Y(n743) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n210) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n211), .Y(n744) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n211) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n212), .Y(n745) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n212) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n213), .Y(n746) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n213) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n214), .Y(n747) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n214) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n215), .Y(n748) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n215) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n216), .Y(n749) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n216) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n217), .Y(n750) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n217) );
  NAND3X1 U401 ( .A(n973), .B(n48), .C(n218), .Y(n209) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n220), .Y(n751) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n220) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n221), .Y(n752) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n221) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n222), .Y(n753) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n222) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n223), .Y(n754) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n223) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n224), .Y(n755) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n224) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n225), .Y(n756) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n225) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n226), .Y(n757) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n226) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n227), .Y(n758) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n227) );
  NAND3X1 U418 ( .A(n70), .B(n48), .C(n228), .Y(n219) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n230), .Y(n759) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n230) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n231), .Y(n760) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n231) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n232), .Y(n761) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n232) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n233), .Y(n762) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n233) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n234), .Y(n763) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n234) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n235), .Y(n764) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n235) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n236), .Y(n765) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n236) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n237), .Y(n766) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n237) );
  NAND3X1 U435 ( .A(n973), .B(n48), .C(n238), .Y(n229) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n240), .Y(n767) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n240) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n241), .Y(n768) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n241) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n242), .Y(n769) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n242) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n243), .Y(n770) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n243) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n244), .Y(n771) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n244) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n245), .Y(n772) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n245) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n246), .Y(n773) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n246) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n247), .Y(n774) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n247) );
  NAND3X1 U452 ( .A(n70), .B(n48), .C(n248), .Y(n239) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n251), .Y(n775) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n251) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n252), .Y(n776) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n252) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n253), .Y(n777) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n253) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n254), .Y(n778) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n254) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n255), .Y(n779) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n255) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n256), .Y(n780) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n256) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n257), .Y(n781) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n257) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n258), .Y(n782) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n258) );
  NAND3X1 U469 ( .A(n973), .B(n48), .C(n259), .Y(n250) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n261), .Y(n783) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n261) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n262), .Y(n784) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n262) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n263), .Y(n785) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n263) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n264), .Y(n786) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n264) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n265), .Y(n787) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n265) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n266), .Y(n788) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n266) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n267), .Y(n789) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n267) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n268), .Y(n790) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n268) );
  NAND3X1 U486 ( .A(n111), .B(n48), .C(n228), .Y(n260) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n270), .Y(n791) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n270) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n271), .Y(n792) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n271) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n272), .Y(n793) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n272) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n273), .Y(n794) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n273) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n274), .Y(n795) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n274) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n275), .Y(n796) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n275) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n276), .Y(n797) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n276) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n277), .Y(n798) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n277) );
  NAND3X1 U503 ( .A(n973), .B(n48), .C(n278), .Y(n269) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n280), .Y(n799) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n280) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n281), .Y(n800) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n281) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n282), .Y(n801) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n282) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n283), .Y(n802) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n283) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n284), .Y(n803) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n284) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n285), .Y(n804) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n285) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n286), .Y(n805) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n286) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n287), .Y(n806) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n287) );
  NAND3X1 U520 ( .A(n111), .B(n48), .C(n248), .Y(n279) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n291), .Y(n807) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n291) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n292), .Y(n808) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n292) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n293), .Y(n809) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n293) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n294), .Y(n810) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n294) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n295), .Y(n811) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n295) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n296), .Y(n812) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n296) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n297), .Y(n813) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n297) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n298), .Y(n814) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n298) );
  NAND3X1 U537 ( .A(n973), .B(n48), .C(n299), .Y(n290) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n301), .Y(n815) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n301) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n302), .Y(n816) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n302) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n303), .Y(n817) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n303) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n304), .Y(n818) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n304) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n305), .Y(n819) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n305) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n306), .Y(n820) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n306) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n307), .Y(n821) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n307) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n308), .Y(n822) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n308) );
  NAND3X1 U554 ( .A(n969), .B(n48), .C(n228), .Y(n300) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n310), .Y(n823) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n310) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n311), .Y(n824) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n311) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n312), .Y(n825) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n312) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n313), .Y(n826) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n313) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n314), .Y(n827) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n314) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n315), .Y(n828) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n315) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n316), .Y(n829) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n316) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n317), .Y(n830) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n317) );
  NAND3X1 U571 ( .A(n973), .B(n48), .C(n318), .Y(n309) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n320), .Y(n831) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n320) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n321), .Y(n832) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n321) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n322), .Y(n833) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n322) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n323), .Y(n834) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n323) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n324), .Y(n835) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n324) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n325), .Y(n836) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n325) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n326), .Y(n837) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n326) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n327), .Y(n838) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n327) );
  NAND3X1 U588 ( .A(n969), .B(n48), .C(n248), .Y(n319) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n330), .Y(n839) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n330) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n331), .Y(n840) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n331) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n332), .Y(n841) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n332) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n333), .Y(n842) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n333) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n334), .Y(n843) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n334) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n335), .Y(n844) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n335) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n336), .Y(n845) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n336) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n337), .Y(n846) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n337) );
  NAND3X1 U606 ( .A(n973), .B(n48), .C(n338), .Y(n329) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n340), .Y(n847) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n340) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n341), .Y(n848) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n341) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n342), .Y(n849) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n342) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n343), .Y(n850) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n343) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n344), .Y(n851) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n344) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n345), .Y(n852) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n345) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n346), .Y(n853) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n346) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n347), .Y(n854) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n347) );
  NAND3X1 U623 ( .A(n967), .B(n48), .C(n228), .Y(n339) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n349), .Y(n855) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n349) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n350), .Y(n856) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n350) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n351), .Y(n857) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n351) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n352), .Y(n858) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n352) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n353), .Y(n859) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n353) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n354), .Y(n860) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n354) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n355), .Y(n861) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n355) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n356), .Y(n862) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n356) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n59) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n359), .Y(n863) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n359) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n360), .Y(n864) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n360) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n361), .Y(n865) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n361) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n362), .Y(n866) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n362) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n363), .Y(n867) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n363) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n364), .Y(n868) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n364) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n365), .Y(n869) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n365) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n366), .Y(n870) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n366) );
  NAND3X1 U658 ( .A(n967), .B(n48), .C(n248), .Y(n358) );
  NOR3X1 U661 ( .A(n370), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n369) );
  NOR3X1 U662 ( .A(n371), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n368) );
  AOI21X1 U663 ( .A(n473), .B(n373), .C(n963), .Y(n1046) );
  OAI21X1 U665 ( .A(rd), .B(n374), .C(wr), .Y(n373) );
  NAND3X1 U667 ( .A(n375), .B(n1025), .C(n376), .Y(n374) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n376) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n375) );
  AOI21X1 U670 ( .A(n460), .B(n378), .C(n1016), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n380), .C(n4), .Y(n378) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n91), .C(\mem<0><1> ), .D(n248), .Y(n383) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n71), .C(\mem<2><1> ), .D(n228), .Y(n382) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n91), .C(\mem<4><1> ), .D(n248), .Y(n385) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n71), .C(\mem<6><1> ), .D(n228), .Y(n384) );
  AOI22X1 U678 ( .A(n288), .B(n893), .C(n249), .D(n933), .Y(n377) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n91), .C(\mem<12><1> ), .D(n248), .Y(
        n389) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n71), .C(\mem<14><1> ), .D(n228), .Y(
        n388) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n91), .C(\mem<8><1> ), .D(n248), .Y(n391) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n71), .C(\mem<10><1> ), .D(n228), .Y(
        n390) );
  AOI21X1 U685 ( .A(n448), .B(n393), .C(n1016), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n940), .B(n395), .C(n950), .Y(n393) );
  AOI21X1 U687 ( .A(n397), .B(n398), .C(n971), .Y(n396) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n91), .C(\mem<0><0> ), .D(n248), .Y(n398) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n71), .C(\mem<2><0> ), .D(n228), .Y(n397) );
  AOI21X1 U690 ( .A(n399), .B(n400), .C(n970), .Y(n394) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n91), .C(\mem<4><0> ), .D(n248), .Y(n400) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n71), .C(\mem<6><0> ), .D(n228), .Y(n399) );
  AOI22X1 U693 ( .A(n288), .B(n891), .C(n249), .D(n931), .Y(n392) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n91), .C(\mem<12><0> ), .D(n248), .Y(
        n404) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n71), .C(\mem<14><0> ), .D(n228), .Y(
        n403) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n91), .C(\mem<8><0> ), .D(n248), .Y(n406) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n71), .C(\mem<10><0> ), .D(n228), .Y(
        n405) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n407) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n199), .C(\mem<19><7> ), .D(n179), .Y(
        n414) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n160), .C(\mem<23><7> ), .D(n140), .Y(
        n413) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n121), .C(\mem<27><7> ), .D(n101), .Y(
        n411) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n81), .C(\mem<31><7> ), .D(n60), .Y(n410) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n357), .C(\mem<3><7> ), .D(n338), .Y(n419) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n318), .C(\mem<7><7> ), .D(n299), .Y(n418) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n278), .C(\mem<11><7> ), .D(n259), .Y(
        n416) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n238), .C(\mem<15><7> ), .D(n218), .Y(
        n415) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n420) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n199), .C(\mem<19><6> ), .D(n179), .Y(
        n427) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n160), .C(\mem<23><6> ), .D(n140), .Y(
        n426) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n121), .C(\mem<27><6> ), .D(n101), .Y(
        n424) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n81), .C(\mem<31><6> ), .D(n60), .Y(n423) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n357), .C(\mem<3><6> ), .D(n338), .Y(n432) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n318), .C(\mem<7><6> ), .D(n299), .Y(n431) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n278), .C(\mem<11><6> ), .D(n259), .Y(
        n429) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n238), .C(\mem<15><6> ), .D(n218), .Y(
        n428) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n433) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n199), .C(\mem<19><5> ), .D(n179), .Y(
        n440) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n160), .C(\mem<23><5> ), .D(n140), .Y(
        n439) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n121), .C(\mem<27><5> ), .D(n101), .Y(
        n437) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n81), .C(\mem<31><5> ), .D(n60), .Y(n436) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n357), .C(\mem<3><5> ), .D(n338), .Y(n445) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n318), .C(\mem<7><5> ), .D(n299), .Y(n444) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n278), .C(\mem<11><5> ), .D(n259), .Y(
        n442) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n238), .C(\mem<15><5> ), .D(n218), .Y(
        n441) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n446) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n199), .C(\mem<19><4> ), .D(n179), .Y(
        n453) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n160), .C(\mem<23><4> ), .D(n140), .Y(
        n452) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n121), .C(\mem<27><4> ), .D(n101), .Y(
        n450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n81), .C(\mem<31><4> ), .D(n60), .Y(n449) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n357), .C(\mem<3><4> ), .D(n338), .Y(n458) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n318), .C(\mem<7><4> ), .D(n299), .Y(n457) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n278), .C(\mem<11><4> ), .D(n259), .Y(
        n455) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n238), .C(\mem<15><4> ), .D(n218), .Y(
        n454) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n459) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n199), .C(\mem<19><3> ), .D(n179), .Y(
        n466) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n160), .C(\mem<23><3> ), .D(n140), .Y(
        n465) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n121), .C(\mem<27><3> ), .D(n101), .Y(
        n463) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n81), .C(\mem<31><3> ), .D(n60), .Y(n462) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n357), .C(\mem<3><3> ), .D(n338), .Y(n471) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n318), .C(\mem<7><3> ), .D(n299), .Y(n470) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n278), .C(\mem<11><3> ), .D(n259), .Y(
        n468) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n238), .C(\mem<15><3> ), .D(n218), .Y(
        n467) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n472) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n199), .C(\mem<19><2> ), .D(n179), .Y(
        n479) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n160), .C(\mem<23><2> ), .D(n140), .Y(
        n478) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n121), .C(\mem<27><2> ), .D(n101), .Y(
        n476) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n81), .C(\mem<31><2> ), .D(n60), .Y(n475) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n357), .C(\mem<3><2> ), .D(n338), .Y(n484) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n318), .C(\mem<7><2> ), .D(n299), .Y(n483) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n278), .C(\mem<11><2> ), .D(n259), .Y(
        n481) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n238), .C(\mem<15><2> ), .D(n218), .Y(
        n480) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n485) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n199), .C(\mem<19><1> ), .D(n179), .Y(
        n492) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n160), .C(\mem<23><1> ), .D(n140), .Y(
        n491) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n121), .C(\mem<27><1> ), .D(n101), .Y(
        n489) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n81), .C(\mem<31><1> ), .D(n60), .Y(n488) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n357), .C(\mem<3><1> ), .D(n338), .Y(n497) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n318), .C(\mem<7><1> ), .D(n299), .Y(n496) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n278), .C(\mem<11><1> ), .D(n259), .Y(
        n494) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n238), .C(\mem<15><1> ), .D(n218), .Y(
        n493) );
  AOI21X1 U777 ( .A(n447), .B(n499), .C(n1016), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n939), .B(n501), .C(n949), .Y(n499) );
  AOI21X1 U779 ( .A(n503), .B(n504), .C(n971), .Y(n502) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n91), .C(\mem<0><7> ), .D(n248), .Y(n504) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n71), .C(\mem<2><7> ), .D(n228), .Y(n503) );
  AOI21X1 U782 ( .A(n505), .B(n506), .C(n970), .Y(n500) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n91), .C(\mem<4><7> ), .D(n248), .Y(n506) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n71), .C(\mem<6><7> ), .D(n228), .Y(n505) );
  AOI22X1 U785 ( .A(n288), .B(n889), .C(n249), .D(n929), .Y(n498) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n91), .C(\mem<12><7> ), .D(n248), .Y(
        n510) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n71), .C(\mem<14><7> ), .D(n228), .Y(
        n509) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n91), .C(\mem<8><7> ), .D(n248), .Y(n512) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n71), .C(\mem<10><7> ), .D(n228), .Y(
        n511) );
  AOI21X1 U792 ( .A(n435), .B(n514), .C(n1016), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n938), .B(n516), .C(n948), .Y(n514) );
  AOI21X1 U794 ( .A(n518), .B(n519), .C(n971), .Y(n517) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n91), .C(\mem<0><6> ), .D(n248), .Y(n519) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n71), .C(\mem<2><6> ), .D(n228), .Y(n518) );
  AOI21X1 U797 ( .A(n520), .B(n521), .C(n970), .Y(n515) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n91), .C(\mem<4><6> ), .D(n248), .Y(n521) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n71), .C(\mem<6><6> ), .D(n228), .Y(n520) );
  AOI22X1 U800 ( .A(n288), .B(n887), .C(n249), .D(n927), .Y(n513) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n91), .C(\mem<12><6> ), .D(n248), .Y(
        n525) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n71), .C(\mem<14><6> ), .D(n228), .Y(
        n524) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n91), .C(\mem<8><6> ), .D(n248), .Y(n527) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n71), .C(\mem<10><6> ), .D(n228), .Y(
        n526) );
  AOI21X1 U807 ( .A(n434), .B(n529), .C(n1016), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n937), .B(n531), .C(n947), .Y(n529) );
  AOI21X1 U809 ( .A(n533), .B(n534), .C(n971), .Y(n532) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n91), .C(\mem<0><5> ), .D(n248), .Y(n534) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n71), .C(\mem<2><5> ), .D(n228), .Y(n533) );
  AOI21X1 U812 ( .A(n535), .B(n536), .C(n970), .Y(n530) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n91), .C(\mem<4><5> ), .D(n248), .Y(n536) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n71), .C(\mem<6><5> ), .D(n228), .Y(n535) );
  AOI22X1 U815 ( .A(n288), .B(n885), .C(n249), .D(n925), .Y(n528) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n91), .C(\mem<12><5> ), .D(n248), .Y(
        n540) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n71), .C(\mem<14><5> ), .D(n228), .Y(
        n539) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n91), .C(\mem<8><5> ), .D(n248), .Y(n542) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n71), .C(\mem<10><5> ), .D(n228), .Y(
        n541) );
  AOI21X1 U822 ( .A(n422), .B(n544), .C(n1016), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n936), .B(n546), .C(n946), .Y(n544) );
  AOI21X1 U824 ( .A(n548), .B(n549), .C(n971), .Y(n547) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n91), .C(\mem<0><4> ), .D(n248), .Y(n549) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n71), .C(\mem<2><4> ), .D(n228), .Y(n548) );
  AOI21X1 U827 ( .A(n550), .B(n551), .C(n970), .Y(n545) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n91), .C(\mem<4><4> ), .D(n248), .Y(n551) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n71), .C(\mem<6><4> ), .D(n228), .Y(n550) );
  AOI22X1 U830 ( .A(n288), .B(n883), .C(n249), .D(n923), .Y(n543) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n91), .C(\mem<12><4> ), .D(n248), .Y(
        n555) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n71), .C(\mem<14><4> ), .D(n228), .Y(
        n554) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n91), .C(\mem<8><4> ), .D(n248), .Y(n557) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n71), .C(\mem<10><4> ), .D(n228), .Y(
        n556) );
  AOI21X1 U837 ( .A(n421), .B(n559), .C(n1016), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n935), .B(n561), .C(n945), .Y(n559) );
  AOI21X1 U839 ( .A(n563), .B(n564), .C(n971), .Y(n562) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n91), .C(\mem<0><3> ), .D(n248), .Y(n564) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n71), .C(\mem<2><3> ), .D(n228), .Y(n563) );
  AOI21X1 U842 ( .A(n565), .B(n566), .C(n970), .Y(n560) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n91), .C(\mem<4><3> ), .D(n248), .Y(n566) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n71), .C(\mem<6><3> ), .D(n228), .Y(n565) );
  AOI22X1 U845 ( .A(n288), .B(n881), .C(n249), .D(n921), .Y(n558) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n91), .C(\mem<12><3> ), .D(n248), .Y(
        n570) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n71), .C(\mem<14><3> ), .D(n228), .Y(
        n569) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n91), .C(\mem<8><3> ), .D(n248), .Y(n572) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n71), .C(\mem<10><3> ), .D(n228), .Y(
        n571) );
  AOI21X1 U852 ( .A(n409), .B(n574), .C(n1016), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n934), .B(n576), .C(n944), .Y(n574) );
  AOI21X1 U854 ( .A(n578), .B(n579), .C(n971), .Y(n577) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n91), .C(\mem<0><2> ), .D(n248), .Y(n579) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n71), .C(\mem<2><2> ), .D(n228), .Y(n578) );
  AOI21X1 U857 ( .A(n580), .B(n581), .C(n970), .Y(n575) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n91), .C(\mem<4><2> ), .D(n248), .Y(n581) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n71), .C(\mem<6><2> ), .D(n228), .Y(n580) );
  AOI22X1 U860 ( .A(n288), .B(n879), .C(n249), .D(n919), .Y(n573) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n91), .C(\mem<12><2> ), .D(n248), .Y(
        n585) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n71), .C(\mem<14><2> ), .D(n228), .Y(
        n584) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n91), .C(\mem<8><2> ), .D(n248), .Y(n587) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n71), .C(\mem<10><2> ), .D(n228), .Y(
        n586) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n588) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n589) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n590) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n199), .C(\mem<19><0> ), .D(n179), .Y(
        n597) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n160), .C(\mem<23><0> ), .D(n140), .Y(
        n596) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n121), .C(\mem<27><0> ), .D(n101), .Y(
        n594) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n81), .C(\mem<31><0> ), .D(n60), .Y(n593) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n357), .C(\mem<3><0> ), .D(n338), .Y(n604) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n367) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n318), .C(\mem<7><0> ), .D(n299), .Y(n603) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n328) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n278), .C(\mem<11><0> ), .D(n259), .Y(
        n601) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n238), .C(\mem<15><0> ), .D(n218), .Y(
        n600) );
  dff_203 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_202 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_185 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_186 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_187 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_188 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_189 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_190 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_191 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_192 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_193 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_194 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_195 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_196 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_197 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_169 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_170 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_171 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_172 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_173 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_174 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_175 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_176 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_177 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_178 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_179 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_180 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_181 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_182 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_183 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_184 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_153 \reg2[0]  ( .q(\data_out<0> ), .d(n1024), .clk(clk), .rst(n1012) );
  dff_154 \reg2[1]  ( .q(\data_out<1> ), .d(n1023), .clk(clk), .rst(n1012) );
  dff_155 \reg2[2]  ( .q(\data_out<2> ), .d(n1022), .clk(clk), .rst(n1012) );
  dff_156 \reg2[3]  ( .q(\data_out<3> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_157 \reg2[4]  ( .q(\data_out<4> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_158 \reg2[5]  ( .q(\data_out<5> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_159 \reg2[6]  ( .q(\data_out<6> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_160 \reg2[7]  ( .q(\data_out<7> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_161 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_162 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_163 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_164 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_165 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_166 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_167 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_168 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_201 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_200 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_199 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_198 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(wr1), .Y(n1025) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n357), .Y(n49) );
  OR2X1 U5 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n371) );
  INVX1 U6 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U7 ( .A(\addr_1c<2> ), .Y(n1028) );
  INVX1 U8 ( .A(\addr_1c<1> ), .Y(n1027) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n370) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n598) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(n1026), .Y(n599) );
  AND2X1 U26 ( .A(n249), .B(n964), .Y(n70) );
  AND2X1 U27 ( .A(n288), .B(n964), .Y(n111) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1029), .Y(n605) );
  AND2X1 U29 ( .A(n1026), .B(n1029), .Y(n606) );
  INVX1 U35 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U36 ( .A(\addr_1c<2> ), .B(n1027), .Y(n288) );
  AND2X1 U37 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n249) );
  AND2X1 U38 ( .A(n599), .B(n249), .Y(n81) );
  AND2X1 U39 ( .A(n288), .B(n598), .Y(n101) );
  AND2X1 U40 ( .A(n288), .B(n599), .Y(n121) );
  AND2X1 U41 ( .A(n941), .B(n598), .Y(n140) );
  AND2X1 U42 ( .A(n941), .B(n599), .Y(n160) );
  AND2X1 U43 ( .A(n598), .B(n951), .Y(n179) );
  AND2X1 U44 ( .A(n599), .B(n951), .Y(n199) );
  AND2X1 U46 ( .A(n605), .B(n249), .Y(n218) );
  AND2X1 U47 ( .A(n249), .B(n606), .Y(n238) );
  AND2X1 U48 ( .A(n605), .B(n288), .Y(n259) );
  AND2X1 U49 ( .A(n288), .B(n606), .Y(n278) );
  AND2X1 U50 ( .A(n605), .B(n941), .Y(n299) );
  AND2X1 U51 ( .A(n941), .B(n606), .Y(n318) );
  OR2X1 U52 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U53 ( .A(n605), .B(n951), .Y(n338) );
  OR2X1 U54 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U55 ( .A(n49), .B(\mem<32><0> ), .Y(n395) );
  AND2X1 U56 ( .A(n49), .B(\mem<32><1> ), .Y(n380) );
  AND2X1 U57 ( .A(n49), .B(\mem<32><2> ), .Y(n576) );
  AND2X1 U58 ( .A(n49), .B(\mem<32><3> ), .Y(n561) );
  AND2X1 U59 ( .A(n49), .B(\mem<32><4> ), .Y(n546) );
  AND2X1 U60 ( .A(n49), .B(\mem<32><5> ), .Y(n531) );
  AND2X1 U61 ( .A(n49), .B(\mem<32><6> ), .Y(n516) );
  AND2X1 U62 ( .A(n49), .B(\mem<32><7> ), .Y(n501) );
  INVX1 U63 ( .A(rd1), .Y(n1016) );
  BUFX2 U64 ( .A(n961), .Y(n1010) );
  BUFX2 U65 ( .A(n961), .Y(n1009) );
  BUFX2 U66 ( .A(n960), .Y(n1007) );
  BUFX2 U67 ( .A(n960), .Y(n1006) );
  BUFX2 U68 ( .A(n959), .Y(n1004) );
  BUFX2 U69 ( .A(n959), .Y(n1003) );
  BUFX2 U70 ( .A(n958), .Y(n1001) );
  BUFX2 U71 ( .A(n958), .Y(n1000) );
  BUFX2 U72 ( .A(n957), .Y(n990) );
  BUFX2 U73 ( .A(n957), .Y(n989) );
  BUFX2 U74 ( .A(n956), .Y(n987) );
  BUFX2 U75 ( .A(n956), .Y(n986) );
  BUFX2 U76 ( .A(n955), .Y(n984) );
  BUFX2 U77 ( .A(n955), .Y(n983) );
  BUFX2 U78 ( .A(n954), .Y(n981) );
  BUFX2 U79 ( .A(n954), .Y(n980) );
  INVX1 U80 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U81 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U82 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U83 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U84 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U85 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U86 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U87 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U88 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U89 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U90 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U91 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U92 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U93 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U129 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U589 ( .A(\data_in_1c<15> ), .Y(n1045) );
  INVX1 U640 ( .A(n590), .Y(n1024) );
  INVX1 U659 ( .A(n485), .Y(n1023) );
  INVX1 U660 ( .A(n472), .Y(n1022) );
  INVX1 U664 ( .A(n459), .Y(n1021) );
  INVX1 U666 ( .A(n446), .Y(n1020) );
  INVX1 U672 ( .A(n433), .Y(n1019) );
  INVX1 U675 ( .A(n420), .Y(n1018) );
  INVX1 U679 ( .A(n407), .Y(n1017) );
  INVX1 U682 ( .A(rst), .Y(n1013) );
  INVX2 U694 ( .A(n1013), .Y(n1012) );
  INVX1 U697 ( .A(wr), .Y(n1015) );
  INVX1 U701 ( .A(rd), .Y(n1014) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n60), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n487), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n474), .B(n486), .Y(n10) );
  OR2X1 U761 ( .A(n522), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n507), .B(n508), .Y(n12) );
  OR2X1 U772 ( .A(n538), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n523), .B(n537), .Y(n14) );
  OR2X1 U789 ( .A(n567), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n552), .B(n553), .Y(n16) );
  OR2X1 U804 ( .A(n583), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n568), .B(n582), .Y(n18) );
  OR2X1 U819 ( .A(n871), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n591), .B(n592), .Y(n20) );
  OR2X1 U834 ( .A(n874), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n872), .B(n873), .Y(n22) );
  OR2X1 U849 ( .A(n877), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n875), .B(n876), .Y(n24) );
  OR2X1 U864 ( .A(n896), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n894), .B(n895), .Y(n26) );
  OR2X1 U875 ( .A(n899), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n897), .B(n898), .Y(n28) );
  OR2X1 U883 ( .A(n902), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n900), .B(n901), .Y(n30) );
  OR2X1 U885 ( .A(n905), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n903), .B(n904), .Y(n32) );
  OR2X1 U887 ( .A(n908), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n906), .B(n907), .Y(n34) );
  OR2X1 U889 ( .A(n911), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n909), .B(n910), .Y(n36) );
  OR2X1 U891 ( .A(n914), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n912), .B(n913), .Y(n38) );
  OR2X1 U893 ( .A(n917), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n915), .B(n916), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n48), .Y(n189) );
  AND2X1 U896 ( .A(n48), .B(n357), .Y(n289) );
  AND2X1 U897 ( .A(n941), .B(n943), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n941), .B(n942), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1046), .Y(err) );
  BUFX2 U906 ( .A(n573), .Y(n409) );
  BUFX2 U907 ( .A(n558), .Y(n421) );
  BUFX2 U908 ( .A(n543), .Y(n422) );
  BUFX2 U909 ( .A(n528), .Y(n434) );
  BUFX2 U910 ( .A(n513), .Y(n435) );
  BUFX2 U911 ( .A(n498), .Y(n447) );
  BUFX2 U912 ( .A(n392), .Y(n448) );
  BUFX2 U913 ( .A(n377), .Y(n460) );
  AND2X2 U914 ( .A(rd), .B(n374), .Y(n461) );
  INVX1 U915 ( .A(n461), .Y(n473) );
  INVX1 U916 ( .A(n602), .Y(n474) );
  INVX1 U917 ( .A(n601), .Y(n486) );
  INVX1 U918 ( .A(n600), .Y(n487) );
  INVX1 U919 ( .A(n495), .Y(n507) );
  INVX1 U920 ( .A(n494), .Y(n508) );
  INVX1 U921 ( .A(n493), .Y(n522) );
  INVX1 U922 ( .A(n482), .Y(n523) );
  INVX1 U923 ( .A(n481), .Y(n537) );
  INVX1 U924 ( .A(n480), .Y(n538) );
  INVX1 U925 ( .A(n469), .Y(n552) );
  INVX1 U926 ( .A(n468), .Y(n553) );
  INVX1 U927 ( .A(n467), .Y(n567) );
  INVX1 U928 ( .A(n456), .Y(n568) );
  INVX1 U929 ( .A(n455), .Y(n582) );
  INVX1 U930 ( .A(n454), .Y(n583) );
  INVX1 U931 ( .A(n443), .Y(n591) );
  INVX1 U932 ( .A(n442), .Y(n592) );
  INVX1 U933 ( .A(n441), .Y(n871) );
  INVX1 U934 ( .A(n430), .Y(n872) );
  INVX1 U935 ( .A(n429), .Y(n873) );
  INVX1 U936 ( .A(n428), .Y(n874) );
  INVX1 U937 ( .A(n417), .Y(n875) );
  INVX1 U938 ( .A(n416), .Y(n876) );
  INVX1 U939 ( .A(n415), .Y(n877) );
  AND2X2 U940 ( .A(n586), .B(n587), .Y(n878) );
  INVX1 U941 ( .A(n878), .Y(n879) );
  AND2X2 U942 ( .A(n571), .B(n572), .Y(n880) );
  INVX1 U943 ( .A(n880), .Y(n881) );
  AND2X2 U944 ( .A(n556), .B(n557), .Y(n882) );
  INVX1 U945 ( .A(n882), .Y(n883) );
  AND2X2 U946 ( .A(n541), .B(n542), .Y(n884) );
  INVX1 U947 ( .A(n884), .Y(n885) );
  AND2X2 U948 ( .A(n526), .B(n527), .Y(n886) );
  INVX1 U949 ( .A(n886), .Y(n887) );
  AND2X2 U950 ( .A(n511), .B(n512), .Y(n888) );
  INVX1 U951 ( .A(n888), .Y(n889) );
  AND2X2 U952 ( .A(n405), .B(n406), .Y(n890) );
  INVX1 U953 ( .A(n890), .Y(n891) );
  AND2X2 U954 ( .A(n390), .B(n391), .Y(n892) );
  INVX1 U955 ( .A(n892), .Y(n893) );
  INVX1 U956 ( .A(n595), .Y(n894) );
  INVX1 U957 ( .A(n594), .Y(n895) );
  INVX1 U958 ( .A(n593), .Y(n896) );
  INVX1 U959 ( .A(n490), .Y(n897) );
  INVX1 U960 ( .A(n489), .Y(n898) );
  INVX1 U961 ( .A(n488), .Y(n899) );
  INVX1 U962 ( .A(n477), .Y(n900) );
  INVX1 U963 ( .A(n476), .Y(n901) );
  INVX1 U964 ( .A(n475), .Y(n902) );
  INVX1 U965 ( .A(n464), .Y(n903) );
  INVX1 U966 ( .A(n463), .Y(n904) );
  INVX1 U967 ( .A(n462), .Y(n905) );
  INVX1 U968 ( .A(n451), .Y(n906) );
  INVX1 U969 ( .A(n450), .Y(n907) );
  INVX1 U970 ( .A(n449), .Y(n908) );
  INVX1 U971 ( .A(n438), .Y(n909) );
  INVX1 U972 ( .A(n437), .Y(n910) );
  INVX1 U973 ( .A(n436), .Y(n911) );
  INVX1 U974 ( .A(n425), .Y(n912) );
  INVX1 U975 ( .A(n424), .Y(n913) );
  INVX1 U976 ( .A(n423), .Y(n914) );
  INVX1 U977 ( .A(n412), .Y(n915) );
  INVX1 U978 ( .A(n411), .Y(n916) );
  INVX1 U979 ( .A(n410), .Y(n917) );
  AND2X2 U980 ( .A(n584), .B(n585), .Y(n918) );
  INVX1 U981 ( .A(n918), .Y(n919) );
  AND2X2 U982 ( .A(n569), .B(n570), .Y(n920) );
  INVX1 U983 ( .A(n920), .Y(n921) );
  AND2X2 U984 ( .A(n554), .B(n555), .Y(n922) );
  INVX1 U985 ( .A(n922), .Y(n923) );
  AND2X2 U986 ( .A(n539), .B(n540), .Y(n924) );
  INVX1 U987 ( .A(n924), .Y(n925) );
  AND2X2 U988 ( .A(n524), .B(n525), .Y(n926) );
  INVX1 U989 ( .A(n926), .Y(n927) );
  AND2X2 U990 ( .A(n509), .B(n510), .Y(n928) );
  INVX1 U991 ( .A(n928), .Y(n929) );
  AND2X2 U992 ( .A(n403), .B(n404), .Y(n930) );
  INVX1 U993 ( .A(n930), .Y(n931) );
  AND2X2 U994 ( .A(n388), .B(n389), .Y(n932) );
  INVX1 U995 ( .A(n932), .Y(n933) );
  BUFX2 U996 ( .A(n575), .Y(n934) );
  BUFX2 U997 ( .A(n560), .Y(n935) );
  BUFX2 U998 ( .A(n545), .Y(n936) );
  BUFX2 U999 ( .A(n530), .Y(n937) );
  BUFX2 U1000 ( .A(n515), .Y(n938) );
  BUFX2 U1001 ( .A(n500), .Y(n939) );
  BUFX2 U1002 ( .A(n394), .Y(n940) );
  INVX1 U1003 ( .A(n970), .Y(n941) );
  INVX1 U1004 ( .A(n385), .Y(n942) );
  INVX1 U1005 ( .A(n384), .Y(n943) );
  BUFX2 U1006 ( .A(n328), .Y(n970) );
  BUFX2 U1007 ( .A(n577), .Y(n944) );
  BUFX2 U1008 ( .A(n562), .Y(n945) );
  BUFX2 U1009 ( .A(n547), .Y(n946) );
  BUFX2 U1010 ( .A(n532), .Y(n947) );
  BUFX2 U1011 ( .A(n517), .Y(n948) );
  BUFX2 U1012 ( .A(n502), .Y(n949) );
  BUFX2 U1013 ( .A(n396), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n383), .Y(n952) );
  INVX1 U1016 ( .A(n382), .Y(n953) );
  BUFX2 U1017 ( .A(n367), .Y(n971) );
  BUFX2 U1018 ( .A(n358), .Y(n972) );
  BUFX2 U1019 ( .A(n339), .Y(n974) );
  BUFX2 U1020 ( .A(n329), .Y(n975) );
  BUFX2 U1021 ( .A(n319), .Y(n976) );
  BUFX2 U1022 ( .A(n309), .Y(n977) );
  BUFX2 U1023 ( .A(n300), .Y(n978) );
  BUFX2 U1024 ( .A(n290), .Y(n979) );
  BUFX2 U1025 ( .A(n269), .Y(n982) );
  BUFX2 U1026 ( .A(n250), .Y(n985) );
  BUFX2 U1027 ( .A(n229), .Y(n988) );
  BUFX2 U1028 ( .A(n209), .Y(n991) );
  BUFX2 U1029 ( .A(n200), .Y(n992) );
  BUFX2 U1030 ( .A(n190), .Y(n993) );
  BUFX2 U1031 ( .A(n180), .Y(n994) );
  BUFX2 U1032 ( .A(n170), .Y(n995) );
  BUFX2 U1033 ( .A(n161), .Y(n996) );
  BUFX2 U1034 ( .A(n151), .Y(n997) );
  BUFX2 U1035 ( .A(n141), .Y(n998) );
  BUFX2 U1036 ( .A(n131), .Y(n999) );
  BUFX2 U1037 ( .A(n112), .Y(n1002) );
  BUFX2 U1038 ( .A(n92), .Y(n1005) );
  BUFX2 U1039 ( .A(n72), .Y(n1008) );
  BUFX2 U1040 ( .A(n59), .Y(n973) );
  AND2X1 U1041 ( .A(n249), .B(n598), .Y(n60) );
  BUFX2 U1042 ( .A(n39), .Y(n1011) );
  BUFX2 U1043 ( .A(n279), .Y(n954) );
  BUFX2 U1044 ( .A(n260), .Y(n955) );
  BUFX2 U1045 ( .A(n239), .Y(n956) );
  BUFX2 U1046 ( .A(n219), .Y(n957) );
  BUFX2 U1047 ( .A(n122), .Y(n958) );
  BUFX2 U1048 ( .A(n102), .Y(n959) );
  BUFX2 U1049 ( .A(n82), .Y(n960) );
  BUFX2 U1050 ( .A(n61), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n368), .B(n369), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n606), .Y(n357) );
endmodule


module final_memory_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U4 ( .A(wr1), .B(n1013), .Y(n1828) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1026), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1026), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1023), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1022), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n964), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1025), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1024), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1024), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n950), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1024), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n949), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1024), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n948), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1024), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n947), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1024), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n946), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1024), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n945), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1024), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n944), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_152 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_151 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_150 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_149 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_148 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_147 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_146 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_145 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_144 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_143 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_142 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_141 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_140 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_139 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_138 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_137 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_136 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_135 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_134 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_133 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_132 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_131 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_130 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_129 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_128 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_127 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_126 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_125 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_124 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_123 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_122 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_121 \reg2[0]  ( .q(\data_out<0> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_120 \reg2[1]  ( .q(\data_out<1> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_119 \reg2[2]  ( .q(\data_out<2> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_118 \reg2[3]  ( .q(\data_out<3> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_117 \reg2[4]  ( .q(\data_out<4> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_116 \reg2[5]  ( .q(\data_out<5> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_115 \reg2[6]  ( .q(\data_out<6> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_114 \reg2[7]  ( .q(\data_out<7> ), .d(n1014), .clk(clk), .rst(n1012) );
  dff_113 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_112 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_111 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_110 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_109 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_108 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_107 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_106 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_105 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_104 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_103 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_102 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  OR2X1 U2 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  INVX1 U7 ( .A(wr1), .Y(n1025) );
  OR2X1 U8 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U23 ( .A(n1630), .B(n964), .Y(n1807) );
  AND2X1 U24 ( .A(n1591), .B(n964), .Y(n1766) );
  INVX1 U25 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U26 ( .A(n1026), .B(n1029), .Y(n1310) );
  AND2X1 U27 ( .A(\addr_1c<0> ), .B(n1029), .Y(n1311) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U29 ( .A(\addr_1c<3> ), .B(n1026), .Y(n1317) );
  INVX1 U35 ( .A(\addr_1c<1> ), .Y(n1027) );
  AND2X1 U36 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U37 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U38 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U39 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U40 ( .A(n1318), .B(n951), .Y(n1699) );
  AND2X1 U41 ( .A(n1317), .B(n951), .Y(n1680) );
  AND2X1 U42 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U43 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U44 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U46 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U47 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U48 ( .A(n1311), .B(n951), .Y(n1542) );
  OR2X1 U49 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U50 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U51 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U52 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U53 ( .A(\addr_1c<2> ), .B(n1027), .Y(n1591) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  BUFX2 U55 ( .A(n961), .Y(n1010) );
  BUFX2 U56 ( .A(n961), .Y(n1009) );
  BUFX2 U57 ( .A(n960), .Y(n1007) );
  BUFX2 U58 ( .A(n960), .Y(n1006) );
  BUFX2 U59 ( .A(n959), .Y(n1004) );
  BUFX2 U60 ( .A(n959), .Y(n1003) );
  BUFX2 U61 ( .A(n958), .Y(n1001) );
  BUFX2 U62 ( .A(n958), .Y(n1000) );
  BUFX2 U63 ( .A(n957), .Y(n990) );
  BUFX2 U64 ( .A(n957), .Y(n989) );
  BUFX2 U65 ( .A(n956), .Y(n987) );
  BUFX2 U66 ( .A(n956), .Y(n986) );
  BUFX2 U67 ( .A(n955), .Y(n984) );
  BUFX2 U68 ( .A(n955), .Y(n983) );
  BUFX2 U69 ( .A(n954), .Y(n981) );
  BUFX2 U70 ( .A(n954), .Y(n980) );
  INVX1 U71 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U72 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U73 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U74 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U75 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U76 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U77 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U78 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U79 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U80 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U81 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U82 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U83 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U84 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U85 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U86 ( .A(\data_in_1c<15> ), .Y(n1045) );
  AND2X1 U87 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U88 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U89 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U90 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U91 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U92 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U93 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U129 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U589 ( .A(rd1), .Y(n1024) );
  INVX1 U640 ( .A(n1324), .Y(n1021) );
  INVX1 U659 ( .A(n1415), .Y(n1020) );
  INVX1 U660 ( .A(n1426), .Y(n1019) );
  INVX1 U664 ( .A(n1437), .Y(n1018) );
  INVX1 U666 ( .A(n1448), .Y(n1017) );
  INVX1 U672 ( .A(n1459), .Y(n1016) );
  INVX1 U675 ( .A(n1470), .Y(n1015) );
  INVX1 U679 ( .A(n1481), .Y(n1014) );
  INVX1 U682 ( .A(rst), .Y(n1013) );
  INVX2 U694 ( .A(n1013), .Y(n1012) );
  INVX1 U697 ( .A(wr), .Y(n1023) );
  INVX1 U701 ( .A(rd), .Y(n1022) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1838), .Y(err) );
  BUFX2 U1007 ( .A(n1335), .Y(n944) );
  BUFX2 U1008 ( .A(n1348), .Y(n945) );
  BUFX2 U1009 ( .A(n1361), .Y(n946) );
  BUFX2 U1010 ( .A(n1374), .Y(n947) );
  BUFX2 U1011 ( .A(n1387), .Y(n948) );
  BUFX2 U1012 ( .A(n1400), .Y(n949) );
  BUFX2 U1013 ( .A(n1490), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n1501), .Y(n952) );
  INVX1 U1016 ( .A(n1502), .Y(n953) );
  BUFX2 U1017 ( .A(n1514), .Y(n971) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n1513), .B(n1512), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n1310), .Y(n1524) );
endmodule


module final_memory_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U4 ( .A(wr1), .B(n1013), .Y(n1828) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1026), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1026), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1023), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1022), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n964), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1025), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1024), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1024), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n949), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1024), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n948), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1024), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n947), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1024), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n946), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1024), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n945), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1024), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n944), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1024), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n943), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_101 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_100 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_99 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_98 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_97 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_96 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_95 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_94 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_93 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_92 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_91 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_90 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_89 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1012) );
  dff_88 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1012) );
  dff_87 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1012) );
  dff_86 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_85 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_84 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_83 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_82 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_81 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_80 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_79 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_78 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_77 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_76 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_75 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_74 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_73 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_72 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_71 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_70 \reg2[0]  ( .q(\data_out<0> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_69 \reg2[1]  ( .q(\data_out<1> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_68 \reg2[2]  ( .q(\data_out<2> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_67 \reg2[3]  ( .q(\data_out<3> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_66 \reg2[4]  ( .q(\data_out<4> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_65 \reg2[5]  ( .q(\data_out<5> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_64 \reg2[6]  ( .q(\data_out<6> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_63 \reg2[7]  ( .q(\data_out<7> ), .d(n1014), .clk(clk), .rst(n1012) );
  dff_62 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1012) );
  dff_61 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1012) );
  dff_60 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_59 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_58 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_57 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_56 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_55 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_54 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_53 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_52 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_51 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  OR2X1 U2 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  INVX1 U7 ( .A(wr1), .Y(n1025) );
  OR2X1 U8 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U23 ( .A(n1630), .B(n964), .Y(n1807) );
  AND2X1 U24 ( .A(n1591), .B(n964), .Y(n1766) );
  INVX1 U25 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U26 ( .A(n1026), .B(n1029), .Y(n1310) );
  AND2X1 U27 ( .A(\addr_1c<0> ), .B(n1029), .Y(n1311) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U29 ( .A(\addr_1c<3> ), .B(n1026), .Y(n1317) );
  INVX1 U35 ( .A(\addr_1c<1> ), .Y(n1027) );
  AND2X1 U36 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U37 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U38 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U39 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U40 ( .A(n1318), .B(n950), .Y(n1699) );
  AND2X1 U41 ( .A(n1317), .B(n950), .Y(n1680) );
  AND2X1 U42 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U43 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U44 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U46 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U47 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U48 ( .A(n1311), .B(n950), .Y(n1542) );
  OR2X1 U49 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U50 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U51 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U52 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U53 ( .A(\addr_1c<2> ), .B(n1027), .Y(n1591) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  BUFX2 U55 ( .A(n961), .Y(n1010) );
  BUFX2 U56 ( .A(n961), .Y(n1009) );
  BUFX2 U57 ( .A(n960), .Y(n1007) );
  BUFX2 U58 ( .A(n960), .Y(n1006) );
  BUFX2 U59 ( .A(n959), .Y(n1004) );
  BUFX2 U60 ( .A(n959), .Y(n1003) );
  BUFX2 U61 ( .A(n958), .Y(n1001) );
  BUFX2 U62 ( .A(n958), .Y(n1000) );
  BUFX2 U63 ( .A(n957), .Y(n990) );
  BUFX2 U64 ( .A(n957), .Y(n989) );
  BUFX2 U65 ( .A(n956), .Y(n987) );
  BUFX2 U66 ( .A(n956), .Y(n986) );
  BUFX2 U67 ( .A(n955), .Y(n984) );
  BUFX2 U68 ( .A(n955), .Y(n983) );
  BUFX2 U69 ( .A(n954), .Y(n981) );
  BUFX2 U70 ( .A(n954), .Y(n980) );
  INVX1 U71 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U72 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U73 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U74 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U75 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U76 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U77 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U78 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U79 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U80 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U81 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U82 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U83 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U84 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U85 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U86 ( .A(\data_in_1c<15> ), .Y(n1045) );
  AND2X1 U87 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U88 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U89 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U90 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U91 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U92 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U93 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U129 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U589 ( .A(rd1), .Y(n1024) );
  INVX1 U640 ( .A(n1324), .Y(n1021) );
  INVX1 U659 ( .A(n1415), .Y(n1020) );
  INVX1 U660 ( .A(n1426), .Y(n1019) );
  INVX1 U664 ( .A(n1437), .Y(n1018) );
  INVX1 U666 ( .A(n1448), .Y(n1017) );
  INVX1 U672 ( .A(n1459), .Y(n1016) );
  INVX1 U675 ( .A(n1470), .Y(n1015) );
  INVX1 U679 ( .A(n1481), .Y(n1014) );
  INVX1 U682 ( .A(rst), .Y(n1013) );
  INVX2 U694 ( .A(n1013), .Y(n1012) );
  INVX1 U697 ( .A(wr), .Y(n1023) );
  INVX1 U701 ( .A(rd), .Y(n1022) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n950), .B(n952), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n950), .B(n951), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1335), .Y(n943) );
  BUFX2 U1007 ( .A(n1348), .Y(n944) );
  BUFX2 U1008 ( .A(n1361), .Y(n945) );
  BUFX2 U1009 ( .A(n1374), .Y(n946) );
  BUFX2 U1010 ( .A(n1387), .Y(n947) );
  BUFX2 U1011 ( .A(n1400), .Y(n948) );
  BUFX2 U1012 ( .A(n1490), .Y(n949) );
  INVX1 U1013 ( .A(n971), .Y(n950) );
  INVX1 U1014 ( .A(n1501), .Y(n951) );
  INVX1 U1015 ( .A(n1502), .Y(n952) );
  BUFX2 U1016 ( .A(n1514), .Y(n971) );
  BUFX2 U1017 ( .A(n1838), .Y(err) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n1513), .B(n1512), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n950), .B(n1310), .Y(n1524) );
endmodule


module final_memory_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U4 ( .A(wr1), .B(n1013), .Y(n1828) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1026), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1026), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1023), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1022), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n964), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1025), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1024), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1024), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n950), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1024), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n949), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1024), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n948), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1024), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n947), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1024), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n946), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1024), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n945), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1024), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n944), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_50 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_49 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_48 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_47 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_46 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_45 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_44 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_43 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_42 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_41 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_40 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_39 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_38 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1012) );
  dff_37 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1012) );
  dff_36 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1012) );
  dff_35 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_34 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_33 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_32 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_31 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_30 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_29 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_28 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_27 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_26 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_25 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_24 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_23 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_22 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_21 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_20 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_19 \reg2[0]  ( .q(\data_out<0> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_18 \reg2[1]  ( .q(\data_out<1> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_17 \reg2[2]  ( .q(\data_out<2> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_16 \reg2[3]  ( .q(\data_out<3> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_15 \reg2[4]  ( .q(\data_out<4> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_14 \reg2[5]  ( .q(\data_out<5> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_13 \reg2[6]  ( .q(\data_out<6> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_12 \reg2[7]  ( .q(\data_out<7> ), .d(n1014), .clk(clk), .rst(n1012) );
  dff_11 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1012) );
  dff_10 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1012) );
  dff_9 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_8 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_7 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_6 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_5 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_4 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_3 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_2 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_1 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_0 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  OR2X1 U2 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  INVX1 U7 ( .A(wr1), .Y(n1025) );
  OR2X1 U8 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U23 ( .A(n1630), .B(n964), .Y(n1807) );
  AND2X1 U24 ( .A(n1591), .B(n964), .Y(n1766) );
  INVX1 U25 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U26 ( .A(n1026), .B(n1029), .Y(n1310) );
  AND2X1 U27 ( .A(\addr_1c<0> ), .B(n1029), .Y(n1311) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U29 ( .A(\addr_1c<3> ), .B(n1026), .Y(n1317) );
  INVX1 U35 ( .A(\addr_1c<1> ), .Y(n1027) );
  AND2X1 U36 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U37 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U38 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U39 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U40 ( .A(n1318), .B(n951), .Y(n1699) );
  AND2X1 U41 ( .A(n1317), .B(n951), .Y(n1680) );
  AND2X1 U42 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U43 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U44 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U46 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U47 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U48 ( .A(n1311), .B(n951), .Y(n1542) );
  OR2X1 U49 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U50 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U51 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U52 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U53 ( .A(\addr_1c<2> ), .B(n1027), .Y(n1591) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  BUFX2 U55 ( .A(n961), .Y(n1010) );
  BUFX2 U56 ( .A(n961), .Y(n1009) );
  BUFX2 U57 ( .A(n960), .Y(n1007) );
  BUFX2 U58 ( .A(n960), .Y(n1006) );
  BUFX2 U59 ( .A(n959), .Y(n1004) );
  BUFX2 U60 ( .A(n959), .Y(n1003) );
  BUFX2 U61 ( .A(n958), .Y(n1001) );
  BUFX2 U62 ( .A(n958), .Y(n1000) );
  BUFX2 U63 ( .A(n957), .Y(n990) );
  BUFX2 U64 ( .A(n957), .Y(n989) );
  BUFX2 U65 ( .A(n956), .Y(n987) );
  BUFX2 U66 ( .A(n956), .Y(n986) );
  BUFX2 U67 ( .A(n955), .Y(n984) );
  BUFX2 U68 ( .A(n955), .Y(n983) );
  BUFX2 U69 ( .A(n954), .Y(n981) );
  BUFX2 U70 ( .A(n954), .Y(n980) );
  INVX1 U71 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U72 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U73 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U74 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U75 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U76 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U77 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U78 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U79 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U80 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U81 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U82 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U83 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U84 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U85 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U86 ( .A(\data_in_1c<15> ), .Y(n1045) );
  AND2X1 U87 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U88 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U89 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U90 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U91 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U92 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U93 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U129 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U589 ( .A(rd1), .Y(n1024) );
  INVX1 U640 ( .A(n1324), .Y(n1021) );
  INVX1 U659 ( .A(n1415), .Y(n1020) );
  INVX1 U660 ( .A(n1426), .Y(n1019) );
  INVX1 U664 ( .A(n1437), .Y(n1018) );
  INVX1 U666 ( .A(n1448), .Y(n1017) );
  INVX1 U672 ( .A(n1459), .Y(n1016) );
  INVX1 U675 ( .A(n1470), .Y(n1015) );
  INVX1 U679 ( .A(n1481), .Y(n1014) );
  INVX1 U682 ( .A(rst), .Y(n1013) );
  INVX2 U694 ( .A(n1013), .Y(n1012) );
  INVX1 U697 ( .A(wr), .Y(n1023) );
  INVX1 U701 ( .A(rd), .Y(n1022) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1838), .Y(err) );
  BUFX2 U1007 ( .A(n1335), .Y(n944) );
  BUFX2 U1008 ( .A(n1348), .Y(n945) );
  BUFX2 U1009 ( .A(n1361), .Y(n946) );
  BUFX2 U1010 ( .A(n1374), .Y(n947) );
  BUFX2 U1011 ( .A(n1387), .Y(n948) );
  BUFX2 U1012 ( .A(n1400), .Y(n949) );
  BUFX2 U1013 ( .A(n1490), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n1501), .Y(n952) );
  INVX1 U1016 ( .A(n1502), .Y(n953) );
  BUFX2 U1017 ( .A(n1514), .Y(n971) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n1513), .B(n1512), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n1310), .Y(n1524) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module cache_cache_id1 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n151, n152, n153, n154, n155, wr_word0, wr_word1, wr_word2, wr_word3,
         \w0<15> , \w0<14> , \w0<13> , \w0<12> , \w0<11> , \w0<10> , \w0<9> ,
         \w0<8> , \w0<7> , \w0<6> , \w0<5> , \w0<4> , \w0<3> , \w0<2> ,
         \w0<1> , \w0<0> , \w1<15> , \w1<14> , \w1<13> , \w1<12> , \w1<11> ,
         \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , \w1<4> ,
         \w1<3> , \w1<2> , \w1<1> , \w1<0> , \w2<15> , \w2<14> , \w2<13> ,
         \w2<12> , \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> ,
         \w2<5> , \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> , \w3<15> ,
         \w3<14> , \w3<13> , \w3<12> , \w3<11> , \w3<10> , \w3<9> , \w3<8> ,
         \w3<7> , \w3<6> , \w3<5> , \w3<4> , \w3<3> , \w3<2> , \w3<1> ,
         \w3<0> , dirtybit, validbit, net58822, net58824, net58855, net58857,
         net58858, net58859, net58860, net58863, net58867, net58875, net62346,
         net65749, net65770, net65818, net65825, net65831, net65893, net72484,
         net73228, net78407, net78431, net81395, net86922, net86921, net96813,
         net97027, net100784, net100783, net101245, net101736, net96812,
         net96811, net58877, net100792, net100786, net97026, net58845,
         net100182, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81,
         n83, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n97, n98, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149;
  assign \tag_out<2>  = net65749;
  assign \tag_out<3>  = net65818;
  assign \tag_out<1>  = net65825;
  assign \tag_out<0>  = net65831;
  assign \tag_out<4>  = net72484;
  assign \data_out<4>  = net97027;

  memc_Size16_7 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({n112, n110, n108, 
        n106, n104, n102, n100, n97}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word0), .clk(clk), .rst(n114), .createdump(createdump), 
        .file_id({1'b0, 1'b1, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_6 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({n112, n110, n108, 
        n106, n104, n102, n100, n97}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word1), .clk(clk), .rst(n114), .createdump(createdump), 
        .file_id({1'b0, 1'b1, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_5 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({n112, n110, n108, 
        n106, n104, n102, n100, n97}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word2), .clk(clk), .rst(n114), .createdump(createdump), 
        .file_id({1'b0, 1'b1, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_4 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({n112, n110, n108, 
        n106, n104, n102, n100, n97}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word3), .clk(clk), .rst(n114), .createdump(createdump), 
        .file_id({1'b0, 1'b1, 1'b0, 1'b1, 1'b1}) );
  memc_Size5_1 mem_tg ( .data_out({n151, n152, n153, n154, n155}), .addr({n112, 
        n110, n108, n106, n104, n102, n100, \index<0> }), .data_in({
        \tag_in<4> , \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), 
        .write(net101245), .clk(clk), .rst(n114), .createdump(createdump), 
        .file_id({1'b0, 1'b1, 1'b1, 1'b0, 1'b0}) );
  memc_Size1_1 mem_dr ( .data_out(dirtybit), .addr({n112, n110, n108, n106, 
        n104, n102, n100, n97}), .data_in(comp), .write(n23), .clk(clk), .rst(
        n114), .createdump(createdump), .file_id({1'b0, 1'b1, 1'b1, 1'b0, 1'b1}) );
  memv_1 mem_vl ( .data_out(validbit), .addr({n112, n110, n108, n106, n104, 
        n102, n100, n22}), .data_in(valid_in), .write(net100784), .clk(clk), 
        .rst(n114), .createdump(createdump), .file_id({1'b0, 1'b1, 1'b0, 1'b0, 
        1'b0}) );
  OR2X1 U3 ( .A(\offset<1> ), .B(net58858), .Y(n88) );
  INVX1 U4 ( .A(\tag_in<0> ), .Y(n7) );
  INVX1 U5 ( .A(\tag_in<3> ), .Y(n9) );
  AND2X1 U6 ( .A(\offset<2> ), .B(\offset<1> ), .Y(net81395) );
  OR2X1 U7 ( .A(\offset<1> ), .B(\offset<2> ), .Y(n90) );
  BUFX2 U8 ( .A(net58822), .Y(net62346) );
  INVX1 U9 ( .A(net78431), .Y(net58824) );
  INVX1 U10 ( .A(\tag_in<1> ), .Y(n6) );
  INVX1 U11 ( .A(\tag_in<2> ), .Y(n8) );
  INVX1 U12 ( .A(n111), .Y(n110) );
  INVX1 U13 ( .A(\index<6> ), .Y(n111) );
  INVX1 U14 ( .A(n113), .Y(n112) );
  INVX1 U15 ( .A(\index<7> ), .Y(n113) );
  INVX1 U16 ( .A(n109), .Y(n108) );
  INVX1 U17 ( .A(\index<5> ), .Y(n109) );
  AND2X1 U18 ( .A(dirtybit), .B(net58867), .Y(n94) );
  BUFX2 U19 ( .A(n2), .Y(n1) );
  AOI22X1 U20 ( .A(net86922), .B(\w1<4> ), .C(\w0<4> ), .D(net62346), .Y(n2)
         );
  INVX1 U21 ( .A(net86921), .Y(net86922) );
  AND2X2 U22 ( .A(net100182), .B(n1), .Y(net97026) );
  INVX1 U23 ( .A(net97026), .Y(net97027) );
  BUFX2 U24 ( .A(net58845), .Y(net100182) );
  AOI22X1 U25 ( .A(net78407), .B(\w3<4> ), .C(\w2<4> ), .D(net58824), .Y(
        net58845) );
  AND2X1 U26 ( .A(net81395), .B(net58857), .Y(net78407) );
  OR2X2 U27 ( .A(n4), .B(n3), .Y(n5) );
  OR2X2 U28 ( .A(n13), .B(n12), .Y(n4) );
  XNOR2X1 U29 ( .A(n152), .B(n9), .Y(n13) );
  XNOR2X1 U30 ( .A(n153), .B(n8), .Y(n12) );
  OR2X2 U31 ( .A(n11), .B(n10), .Y(n3) );
  XNOR2X1 U32 ( .A(n155), .B(n7), .Y(n11) );
  XNOR2X1 U33 ( .A(n154), .B(n6), .Y(n10) );
  OR2X2 U34 ( .A(net100786), .B(n5), .Y(net100792) );
  AND2X2 U35 ( .A(net58867), .B(net58877), .Y(net96811) );
  INVX1 U36 ( .A(net58863), .Y(net58867) );
  INVX1 U37 ( .A(net100792), .Y(net58877) );
  INVX1 U38 ( .A(net96811), .Y(net101736) );
  INVX1 U39 ( .A(net96811), .Y(net96812) );
  INVX1 U40 ( .A(net96811), .Y(net96813) );
  AND2X2 U41 ( .A(n17), .B(n15), .Y(net100786) );
  INVX1 U42 ( .A(n16), .Y(n17) );
  AND2X2 U43 ( .A(\tag_in<4> ), .B(n151), .Y(n16) );
  NAND2X1 U44 ( .A(n14), .B(net65893), .Y(n15) );
  INVX1 U45 ( .A(\tag_in<4> ), .Y(n14) );
  INVX1 U46 ( .A(n151), .Y(net65893) );
  BUFX2 U47 ( .A(net100792), .Y(net65770) );
  AND2X2 U48 ( .A(n20), .B(n18), .Y(wr_word1) );
  INVX1 U49 ( .A(n19), .Y(n20) );
  OR2X1 U50 ( .A(net58860), .B(\offset<2> ), .Y(n19) );
  INVX1 U51 ( .A(\offset<1> ), .Y(net58860) );
  OAI21X1 U52 ( .A(net58875), .B(net96812), .C(net73228), .Y(n18) );
  INVX1 U53 ( .A(write), .Y(net58875) );
  INVX1 U54 ( .A(net100784), .Y(net73228) );
  OAI21X1 U55 ( .A(net58875), .B(net101736), .C(net73228), .Y(n21) );
  INVX1 U56 ( .A(rst), .Y(n115) );
  BUFX2 U57 ( .A(\index<0> ), .Y(n22) );
  OAI21X1 U58 ( .A(net101736), .B(net58875), .C(net73228), .Y(n23) );
  OAI21X1 U59 ( .A(net58875), .B(net96813), .C(net73228), .Y(n24) );
  INVX1 U60 ( .A(comp), .Y(n116) );
  INVX1 U61 ( .A(net100783), .Y(net101245) );
  OR2X2 U62 ( .A(n117), .B(net58863), .Y(net100783) );
  INVX1 U63 ( .A(net100783), .Y(net100784) );
  BUFX2 U64 ( .A(n119), .Y(n25) );
  BUFX2 U65 ( .A(n122), .Y(n26) );
  BUFX2 U66 ( .A(n124), .Y(n27) );
  BUFX2 U67 ( .A(n126), .Y(n28) );
  BUFX2 U68 ( .A(n128), .Y(n29) );
  BUFX2 U69 ( .A(n130), .Y(n30) );
  BUFX2 U70 ( .A(n132), .Y(n31) );
  BUFX2 U71 ( .A(n134), .Y(n32) );
  BUFX2 U72 ( .A(n136), .Y(n33) );
  BUFX2 U73 ( .A(n138), .Y(n34) );
  BUFX2 U74 ( .A(n140), .Y(n35) );
  BUFX2 U75 ( .A(n141), .Y(n36) );
  BUFX2 U76 ( .A(n143), .Y(n37) );
  BUFX2 U77 ( .A(n146), .Y(n38) );
  BUFX2 U78 ( .A(n147), .Y(n39) );
  BUFX2 U79 ( .A(n120), .Y(n40) );
  BUFX2 U80 ( .A(n121), .Y(n41) );
  BUFX2 U81 ( .A(n123), .Y(n42) );
  BUFX2 U82 ( .A(n125), .Y(n43) );
  BUFX2 U83 ( .A(n127), .Y(n44) );
  BUFX2 U84 ( .A(n129), .Y(n45) );
  BUFX2 U85 ( .A(n131), .Y(n46) );
  BUFX2 U86 ( .A(n133), .Y(n47) );
  BUFX2 U87 ( .A(n135), .Y(n48) );
  BUFX2 U88 ( .A(n137), .Y(n49) );
  BUFX2 U89 ( .A(n139), .Y(n50) );
  BUFX2 U90 ( .A(n142), .Y(n51) );
  BUFX2 U91 ( .A(n144), .Y(n52) );
  BUFX2 U92 ( .A(n145), .Y(n53) );
  BUFX2 U93 ( .A(n148), .Y(n54) );
  AND2X2 U94 ( .A(comp), .B(net65770), .Y(n55) );
  INVX1 U95 ( .A(n55), .Y(n56) );
  AND2X2 U96 ( .A(n25), .B(n40), .Y(n57) );
  INVX1 U97 ( .A(n57), .Y(\data_out<0> ) );
  AND2X2 U98 ( .A(n41), .B(n26), .Y(n59) );
  INVX1 U99 ( .A(n59), .Y(\data_out<1> ) );
  AND2X2 U100 ( .A(n27), .B(n42), .Y(n61) );
  INVX1 U101 ( .A(n61), .Y(\data_out<2> ) );
  AND2X2 U102 ( .A(n28), .B(n43), .Y(n63) );
  INVX1 U103 ( .A(n63), .Y(\data_out<3> ) );
  AND2X2 U104 ( .A(n44), .B(n29), .Y(n65) );
  INVX1 U105 ( .A(n65), .Y(\data_out<5> ) );
  AND2X2 U106 ( .A(n30), .B(n45), .Y(n67) );
  INVX1 U107 ( .A(n67), .Y(\data_out<6> ) );
  AND2X2 U108 ( .A(n31), .B(n46), .Y(n69) );
  INVX1 U109 ( .A(n69), .Y(\data_out<7> ) );
  AND2X2 U110 ( .A(n32), .B(n47), .Y(n71) );
  INVX1 U111 ( .A(n71), .Y(\data_out<8> ) );
  AND2X2 U112 ( .A(n33), .B(n48), .Y(n73) );
  INVX1 U113 ( .A(n73), .Y(\data_out<9> ) );
  AND2X2 U114 ( .A(n34), .B(n49), .Y(n75) );
  INVX1 U115 ( .A(n75), .Y(\data_out<10> ) );
  AND2X2 U116 ( .A(n35), .B(n50), .Y(n77) );
  INVX1 U117 ( .A(n77), .Y(\data_out<11> ) );
  AND2X2 U118 ( .A(n51), .B(n36), .Y(n79) );
  INVX1 U119 ( .A(n79), .Y(\data_out<12> ) );
  AND2X2 U120 ( .A(n37), .B(n52), .Y(n81) );
  INVX1 U121 ( .A(n81), .Y(\data_out<13> ) );
  AND2X2 U122 ( .A(n53), .B(n38), .Y(n83) );
  INVX1 U123 ( .A(n83), .Y(\data_out<14> ) );
  AND2X2 U124 ( .A(n54), .B(n39), .Y(n85) );
  INVX1 U125 ( .A(n85), .Y(\data_out<15> ) );
  OR2X1 U126 ( .A(net58860), .B(n87), .Y(net86921) );
  OR2X1 U127 ( .A(\offset<2> ), .B(net58855), .Y(n87) );
  INVX1 U128 ( .A(n88), .Y(n89) );
  INVX1 U129 ( .A(n90), .Y(n91) );
  OR2X2 U130 ( .A(n118), .B(net58863), .Y(n92) );
  INVX1 U131 ( .A(n92), .Y(n93) );
  INVX1 U132 ( .A(n94), .Y(n95) );
  BUFX2 U133 ( .A(n149), .Y(dirty) );
  BUFX2 U134 ( .A(net58859), .Y(net78431) );
  INVX1 U135 ( .A(net58855), .Y(net58857) );
  INVX1 U136 ( .A(\offset<2> ), .Y(net58858) );
  INVX1 U137 ( .A(net65893), .Y(net72484) );
  BUFX2 U138 ( .A(n22), .Y(n97) );
  INVX1 U139 ( .A(n98), .Y(err) );
  INVX1 U140 ( .A(\offset<0> ), .Y(n98) );
  INVX1 U141 ( .A(n117), .Y(n118) );
  BUFX2 U142 ( .A(n155), .Y(net65831) );
  BUFX2 U143 ( .A(n154), .Y(net65825) );
  BUFX2 U144 ( .A(n152), .Y(net65818) );
  BUFX2 U145 ( .A(n153), .Y(net65749) );
  INVX1 U146 ( .A(net101736), .Y(hit) );
  INVX8 U147 ( .A(n101), .Y(n100) );
  INVX8 U148 ( .A(\index<1> ), .Y(n101) );
  INVX8 U149 ( .A(n103), .Y(n102) );
  INVX8 U150 ( .A(\index<2> ), .Y(n103) );
  INVX8 U151 ( .A(n105), .Y(n104) );
  INVX8 U152 ( .A(\index<3> ), .Y(n105) );
  INVX8 U153 ( .A(n107), .Y(n106) );
  INVX8 U154 ( .A(\index<4> ), .Y(n107) );
  INVX8 U155 ( .A(n115), .Y(n114) );
  NAND2X1 U156 ( .A(enable), .B(n115), .Y(net58863) );
  NAND2X1 U157 ( .A(write), .B(n116), .Y(n117) );
  AND2X2 U158 ( .A(net81395), .B(n24), .Y(wr_word3) );
  AND2X2 U159 ( .A(n24), .B(n89), .Y(wr_word2) );
  AND2X2 U160 ( .A(n91), .B(n21), .Y(wr_word0) );
  AND2X2 U161 ( .A(validbit), .B(n93), .Y(valid) );
  AOI21X1 U162 ( .A(write), .B(n56), .C(n95), .Y(n149) );
  OR2X2 U163 ( .A(write), .B(net58863), .Y(net58855) );
  NAND3X1 U164 ( .A(\offset<2> ), .B(net58857), .C(net58860), .Y(net58859) );
  AOI22X1 U165 ( .A(net78407), .B(\w3<0> ), .C(\w2<0> ), .D(net58824), .Y(n120) );
  NOR3X1 U166 ( .A(\offset<2> ), .B(net58855), .C(\offset<1> ), .Y(net58822)
         );
  AOI22X1 U167 ( .A(net86922), .B(\w1<0> ), .C(net62346), .D(\w0<0> ), .Y(n119) );
  AOI22X1 U168 ( .A(net78407), .B(\w3<1> ), .C(net58824), .D(\w2<1> ), .Y(n122) );
  AOI22X1 U169 ( .A(net86922), .B(\w1<1> ), .C(net62346), .D(\w0<1> ), .Y(n121) );
  AOI22X1 U170 ( .A(net78407), .B(\w3<2> ), .C(net58824), .D(\w2<2> ), .Y(n124) );
  AOI22X1 U171 ( .A(net86922), .B(\w1<2> ), .C(\w0<2> ), .D(net62346), .Y(n123) );
  AOI22X1 U172 ( .A(net78407), .B(\w3<3> ), .C(net58824), .D(\w2<3> ), .Y(n126) );
  AOI22X1 U173 ( .A(net86922), .B(\w1<3> ), .C(net62346), .D(\w0<3> ), .Y(n125) );
  AOI22X1 U174 ( .A(\w3<5> ), .B(net78407), .C(\w2<5> ), .D(net58824), .Y(n128) );
  AOI22X1 U175 ( .A(net86922), .B(\w1<5> ), .C(\w0<5> ), .D(net62346), .Y(n127) );
  AOI22X1 U176 ( .A(net78407), .B(\w3<6> ), .C(net58824), .D(\w2<6> ), .Y(n130) );
  AOI22X1 U177 ( .A(net86922), .B(\w1<6> ), .C(net62346), .D(\w0<6> ), .Y(n129) );
  AOI22X1 U178 ( .A(\w3<7> ), .B(net78407), .C(\w2<7> ), .D(net58824), .Y(n132) );
  AOI22X1 U179 ( .A(net86922), .B(\w1<7> ), .C(\w0<7> ), .D(net62346), .Y(n131) );
  AOI22X1 U180 ( .A(net78407), .B(\w3<8> ), .C(\w2<8> ), .D(net58824), .Y(n134) );
  AOI22X1 U181 ( .A(net86922), .B(\w1<8> ), .C(\w0<8> ), .D(net62346), .Y(n133) );
  AOI22X1 U182 ( .A(net78407), .B(\w3<9> ), .C(net58824), .D(\w2<9> ), .Y(n136) );
  AOI22X1 U183 ( .A(net86922), .B(\w1<9> ), .C(net62346), .D(\w0<9> ), .Y(n135) );
  AOI22X1 U184 ( .A(\w3<10> ), .B(net78407), .C(net58824), .D(\w2<10> ), .Y(
        n138) );
  AOI22X1 U185 ( .A(net86922), .B(\w1<10> ), .C(\w0<10> ), .D(net62346), .Y(
        n137) );
  AOI22X1 U186 ( .A(net78407), .B(\w3<11> ), .C(\w2<11> ), .D(net58824), .Y(
        n140) );
  AOI22X1 U187 ( .A(net86922), .B(\w1<11> ), .C(\w0<11> ), .D(net62346), .Y(
        n139) );
  AOI22X1 U188 ( .A(net78407), .B(\w3<12> ), .C(net58824), .D(\w2<12> ), .Y(
        n142) );
  AOI22X1 U189 ( .A(net86922), .B(\w1<12> ), .C(\w0<12> ), .D(net62346), .Y(
        n141) );
  AOI22X1 U190 ( .A(net78407), .B(\w3<13> ), .C(net58824), .D(\w2<13> ), .Y(
        n144) );
  AOI22X1 U191 ( .A(net86922), .B(\w1<13> ), .C(net62346), .D(\w0<13> ), .Y(
        n143) );
  AOI22X1 U192 ( .A(net78407), .B(\w3<14> ), .C(net58824), .D(\w2<14> ), .Y(
        n146) );
  AOI22X1 U193 ( .A(net86922), .B(\w1<14> ), .C(net62346), .D(\w0<14> ), .Y(
        n145) );
  AOI22X1 U194 ( .A(\w3<15> ), .B(net78407), .C(\w2<15> ), .D(net58824), .Y(
        n148) );
  AOI22X1 U195 ( .A(net86922), .B(\w1<15> ), .C(\w0<15> ), .D(net62346), .Y(
        n147) );
endmodule


module cache_cache_id3 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n195, n196, n197, n198, n199, wr_word0, wr_word1, wr_word2, wr_word3,
         \w0<15> , \w0<14> , \w0<13> , \w0<12> , \w0<11> , \w0<10> , \w0<9> ,
         \w0<8> , \w0<7> , \w0<6> , \w0<5> , \w0<4> , \w0<3> , \w0<2> ,
         \w0<1> , \w0<0> , \w1<15> , \w1<14> , \w1<13> , \w1<12> , \w1<11> ,
         \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , \w1<4> ,
         \w1<3> , \w1<2> , \w1<1> , \w1<0> , \w2<15> , \w2<14> , \w2<13> ,
         \w2<12> , \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> ,
         \w2<5> , \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> , \w3<15> ,
         \w3<14> , \w3<13> , \w3<12> , \w3<11> , \w3<10> , \w3<9> , \w3<8> ,
         \w3<7> , \w3<6> , \w3<5> , \w3<4> , \w3<3> , \w3<2> , \w3<1> ,
         \w3<0> , dirtybit, validbit, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n54,
         n56, n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82,
         n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n116, n120, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n194;

  memc_Size16_3 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({n139, n137, n135, 
        n133, n131, n3, n127, n116}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word0), .clk(clk), .rst(n141), .createdump(createdump), 
        .file_id({1'b1, 1'b1, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_2 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({n139, n137, n135, 
        n133, n131, n3, n127, n116}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word1), .clk(clk), .rst(n141), .createdump(createdump), 
        .file_id({1'b1, 1'b1, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_1 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({n139, n137, n135, 
        n133, n131, n3, n127, n116}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word2), .clk(clk), .rst(n141), .createdump(createdump), 
        .file_id({1'b1, 1'b1, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_0 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({n139, n137, n135, 
        n133, n131, n3, n127, n116}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word3), .clk(clk), .rst(n141), .createdump(createdump), 
        .file_id({1'b1, 1'b1, 1'b0, 1'b1, 1'b1}) );
  memc_Size5_0 mem_tg ( .data_out({n195, n196, n197, n198, n199}), .addr({n139, 
        n137, n135, n133, n131, n129, n127, n12}), .data_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .write(n108), 
        .clk(clk), .rst(n141), .createdump(createdump), .file_id({1'b1, 1'b1, 
        1'b1, 1'b0, 1'b0}) );
  memc_Size1_0 mem_dr ( .data_out(dirtybit), .addr({n139, n137, n135, n133, 
        n131, n3, n127, n116}), .data_in(comp), .write(n1), .clk(clk), .rst(
        n141), .createdump(createdump), .file_id({1'b1, 1'b1, 1'b1, 1'b0, 1'b1}) );
  memv_0 mem_vl ( .data_out(validbit), .addr({n139, n137, n135, n133, n131, 
        n129, n127, n125}), .data_in(valid_in), .write(n109), .clk(clk), .rst(
        n141), .createdump(createdump), .file_id({1'b1, 1'b1, 1'b0, 1'b0, 1'b0}) );
  OAI21X1 U3 ( .A(n88), .B(n150), .C(n149), .Y(n1) );
  INVX1 U4 ( .A(n13), .Y(n14) );
  INVX1 U5 ( .A(\tag_in<3> ), .Y(n9) );
  OR2X1 U6 ( .A(\offset<1> ), .B(\offset<2> ), .Y(n97) );
  OR2X1 U7 ( .A(\offset<1> ), .B(n155), .Y(n93) );
  INVX1 U8 ( .A(\index<4> ), .Y(n134) );
  AND2X1 U9 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n103) );
  BUFX2 U10 ( .A(n189), .Y(n124) );
  INVX1 U11 ( .A(n105), .Y(n188) );
  INVX1 U12 ( .A(\tag_in<2> ), .Y(n2) );
  INVX1 U13 ( .A(\tag_in<1> ), .Y(n8) );
  INVX1 U14 ( .A(\tag_in<0> ), .Y(n11) );
  INVX1 U15 ( .A(\index<5> ), .Y(n136) );
  INVX1 U16 ( .A(n138), .Y(n137) );
  INVX1 U17 ( .A(\index<6> ), .Y(n138) );
  INVX1 U18 ( .A(n140), .Y(n139) );
  INVX1 U19 ( .A(\index<7> ), .Y(n140) );
  AND2X1 U20 ( .A(dirtybit), .B(n153), .Y(n101) );
  AND2X1 U21 ( .A(n17), .B(n33), .Y(n52) );
  INVX1 U22 ( .A(n136), .Y(n135) );
  AND2X2 U23 ( .A(n29), .B(n45), .Y(n76) );
  XNOR2X1 U24 ( .A(n197), .B(n2), .Y(n145) );
  INVX1 U25 ( .A(n130), .Y(n3) );
  INVX4 U26 ( .A(\index<2> ), .Y(n130) );
  AND2X2 U27 ( .A(comp), .B(n120), .Y(n4) );
  INVX1 U28 ( .A(n4), .Y(n5) );
  AND2X2 U29 ( .A(write), .B(n143), .Y(n6) );
  INVX1 U30 ( .A(n6), .Y(n7) );
  XNOR2X1 U31 ( .A(n198), .B(n8), .Y(n147) );
  XNOR2X1 U32 ( .A(n196), .B(n9), .Y(n144) );
  BUFX2 U33 ( .A(n148), .Y(n10) );
  XNOR2X1 U34 ( .A(n199), .B(n11), .Y(n146) );
  INVX2 U35 ( .A(n126), .Y(n12) );
  INVX1 U36 ( .A(n126), .Y(n125) );
  INVX8 U37 ( .A(rst), .Y(n142) );
  INVX8 U38 ( .A(n142), .Y(n141) );
  INVX4 U39 ( .A(\index<1> ), .Y(n128) );
  INVX1 U40 ( .A(comp), .Y(n143) );
  INVX1 U41 ( .A(\index<0> ), .Y(n126) );
  AND2X2 U42 ( .A(enable), .B(n142), .Y(n13) );
  OR2X2 U43 ( .A(n7), .B(n14), .Y(n15) );
  BUFX2 U44 ( .A(n159), .Y(n16) );
  BUFX2 U45 ( .A(n161), .Y(n17) );
  BUFX2 U46 ( .A(n163), .Y(n18) );
  BUFX2 U47 ( .A(n165), .Y(n19) );
  BUFX2 U48 ( .A(n167), .Y(n20) );
  BUFX2 U49 ( .A(n169), .Y(n21) );
  BUFX2 U50 ( .A(n171), .Y(n22) );
  BUFX2 U51 ( .A(n173), .Y(n23) );
  BUFX2 U52 ( .A(n175), .Y(n24) );
  BUFX2 U53 ( .A(n177), .Y(n25) );
  BUFX2 U54 ( .A(n179), .Y(n26) );
  BUFX2 U55 ( .A(n181), .Y(n27) );
  BUFX2 U56 ( .A(n183), .Y(n28) );
  BUFX2 U57 ( .A(n185), .Y(n29) );
  BUFX2 U58 ( .A(n187), .Y(n30) );
  BUFX2 U59 ( .A(n191), .Y(n31) );
  BUFX2 U60 ( .A(n158), .Y(n32) );
  BUFX2 U61 ( .A(n160), .Y(n33) );
  BUFX2 U62 ( .A(n162), .Y(n34) );
  BUFX2 U63 ( .A(n164), .Y(n35) );
  BUFX2 U64 ( .A(n166), .Y(n36) );
  BUFX2 U65 ( .A(n168), .Y(n37) );
  BUFX2 U66 ( .A(n170), .Y(n38) );
  BUFX2 U67 ( .A(n172), .Y(n39) );
  BUFX2 U68 ( .A(n174), .Y(n40) );
  BUFX2 U69 ( .A(n176), .Y(n41) );
  BUFX2 U70 ( .A(n178), .Y(n42) );
  BUFX2 U71 ( .A(n180), .Y(n43) );
  BUFX2 U72 ( .A(n182), .Y(n44) );
  BUFX2 U73 ( .A(n184), .Y(n45) );
  BUFX2 U74 ( .A(n186), .Y(n46) );
  BUFX2 U75 ( .A(n190), .Y(n47) );
  AND2X2 U76 ( .A(n111), .B(n112), .Y(n48) );
  INVX1 U77 ( .A(n48), .Y(n49) );
  AND2X2 U78 ( .A(n16), .B(n32), .Y(n50) );
  INVX1 U79 ( .A(n50), .Y(\data_out<0> ) );
  INVX1 U80 ( .A(n52), .Y(\data_out<1> ) );
  AND2X2 U81 ( .A(n18), .B(n34), .Y(n54) );
  INVX1 U82 ( .A(n54), .Y(\data_out<2> ) );
  AND2X2 U83 ( .A(n19), .B(n35), .Y(n56) );
  INVX1 U84 ( .A(n56), .Y(\data_out<3> ) );
  AND2X2 U85 ( .A(n20), .B(n36), .Y(n58) );
  INVX1 U86 ( .A(n58), .Y(\data_out<4> ) );
  AND2X2 U87 ( .A(n21), .B(n37), .Y(n60) );
  INVX1 U88 ( .A(n60), .Y(\data_out<5> ) );
  AND2X2 U89 ( .A(n22), .B(n38), .Y(n62) );
  INVX1 U90 ( .A(n62), .Y(\data_out<6> ) );
  AND2X2 U91 ( .A(n23), .B(n39), .Y(n64) );
  INVX1 U92 ( .A(n64), .Y(\data_out<7> ) );
  AND2X2 U93 ( .A(n24), .B(n40), .Y(n66) );
  INVX1 U94 ( .A(n66), .Y(\data_out<8> ) );
  AND2X2 U95 ( .A(n25), .B(n41), .Y(n68) );
  INVX1 U96 ( .A(n68), .Y(\data_out<9> ) );
  AND2X2 U97 ( .A(n26), .B(n42), .Y(n70) );
  INVX1 U98 ( .A(n70), .Y(\data_out<10> ) );
  AND2X2 U99 ( .A(n27), .B(n43), .Y(n72) );
  INVX1 U100 ( .A(n72), .Y(\data_out<11> ) );
  AND2X2 U101 ( .A(n28), .B(n44), .Y(n74) );
  INVX1 U102 ( .A(n74), .Y(\data_out<12> ) );
  INVX1 U103 ( .A(n76), .Y(\data_out<13> ) );
  AND2X2 U104 ( .A(n30), .B(n46), .Y(n78) );
  INVX1 U105 ( .A(n78), .Y(\data_out<14> ) );
  AND2X2 U106 ( .A(n31), .B(n47), .Y(n80) );
  INVX1 U107 ( .A(n80), .Y(\data_out<15> ) );
  OR2X2 U108 ( .A(n146), .B(n147), .Y(n82) );
  INVX1 U109 ( .A(n82), .Y(n83) );
  INVX1 U110 ( .A(hit), .Y(n84) );
  OR2X2 U111 ( .A(n144), .B(n145), .Y(n85) );
  INVX1 U112 ( .A(n85), .Y(n86) );
  AND2X2 U113 ( .A(n153), .B(n148), .Y(hit) );
  INVX1 U114 ( .A(hit), .Y(n88) );
  INVX1 U115 ( .A(n195), .Y(n89) );
  OR2X1 U116 ( .A(n106), .B(n92), .Y(n90) );
  INVX1 U117 ( .A(n90), .Y(n91) );
  OR2X1 U118 ( .A(\offset<2> ), .B(n157), .Y(n92) );
  INVX1 U119 ( .A(n93), .Y(n94) );
  OR2X1 U120 ( .A(n106), .B(\offset<2> ), .Y(n95) );
  INVX1 U121 ( .A(n95), .Y(n96) );
  INVX1 U122 ( .A(n97), .Y(n98) );
  OR2X2 U123 ( .A(n151), .B(n14), .Y(n99) );
  INVX1 U124 ( .A(n99), .Y(n100) );
  INVX1 U125 ( .A(n101), .Y(n102) );
  BUFX2 U126 ( .A(n194), .Y(dirty) );
  BUFX2 U127 ( .A(n154), .Y(n105) );
  INVX1 U128 ( .A(\offset<1> ), .Y(n106) );
  INVX1 U129 ( .A(n157), .Y(n156) );
  INVX1 U130 ( .A(\offset<2> ), .Y(n155) );
  AND2X1 U131 ( .A(n103), .B(n156), .Y(n107) );
  INVX1 U132 ( .A(n15), .Y(n108) );
  INVX1 U133 ( .A(n15), .Y(n109) );
  NAND2X1 U134 ( .A(\tag_in<4> ), .B(n195), .Y(n111) );
  NAND2X1 U135 ( .A(n110), .B(n89), .Y(n112) );
  INVX1 U136 ( .A(\tag_in<4> ), .Y(n110) );
  INVX1 U137 ( .A(n12), .Y(n113) );
  INVX1 U138 ( .A(n114), .Y(err) );
  INVX1 U139 ( .A(\offset<0> ), .Y(n114) );
  INVX1 U140 ( .A(n113), .Y(n116) );
  BUFX2 U141 ( .A(n195), .Y(\tag_out<4> ) );
  BUFX2 U142 ( .A(n199), .Y(\tag_out<0> ) );
  BUFX2 U143 ( .A(n198), .Y(\tag_out<1> ) );
  INVX1 U144 ( .A(n109), .Y(n149) );
  INVX1 U145 ( .A(n14), .Y(n153) );
  INVX1 U146 ( .A(n7), .Y(n151) );
  INVX1 U147 ( .A(write), .Y(n150) );
  INVX1 U148 ( .A(n10), .Y(n120) );
  BUFX2 U149 ( .A(n196), .Y(\tag_out<3> ) );
  BUFX2 U150 ( .A(n197), .Y(\tag_out<2> ) );
  INVX1 U151 ( .A(n152), .Y(n148) );
  OAI21X1 U152 ( .A(n150), .B(n84), .C(n149), .Y(n123) );
  INVX8 U153 ( .A(n128), .Y(n127) );
  INVX8 U154 ( .A(n130), .Y(n129) );
  INVX8 U155 ( .A(n132), .Y(n131) );
  INVX8 U156 ( .A(\index<3> ), .Y(n132) );
  INVX8 U157 ( .A(n134), .Y(n133) );
  NAND3X1 U158 ( .A(n49), .B(n83), .C(n86), .Y(n152) );
  OAI21X1 U159 ( .A(n88), .B(n150), .C(n149), .Y(n192) );
  AND2X2 U160 ( .A(n103), .B(n123), .Y(wr_word3) );
  AND2X2 U161 ( .A(n123), .B(n94), .Y(wr_word2) );
  AND2X2 U162 ( .A(n96), .B(n192), .Y(wr_word1) );
  AND2X2 U163 ( .A(n123), .B(n98), .Y(wr_word0) );
  AND2X2 U164 ( .A(validbit), .B(n100), .Y(valid) );
  AOI21X1 U165 ( .A(write), .B(n5), .C(n102), .Y(n194) );
  OR2X2 U166 ( .A(write), .B(n14), .Y(n157) );
  NAND3X1 U167 ( .A(\offset<2> ), .B(n156), .C(n106), .Y(n154) );
  AOI22X1 U168 ( .A(\w3<0> ), .B(n107), .C(\w2<0> ), .D(n188), .Y(n159) );
  NOR3X1 U169 ( .A(\offset<2> ), .B(n157), .C(\offset<1> ), .Y(n189) );
  AOI22X1 U170 ( .A(\w1<0> ), .B(n91), .C(\w0<0> ), .D(n124), .Y(n158) );
  AOI22X1 U171 ( .A(\w3<1> ), .B(n107), .C(\w2<1> ), .D(n188), .Y(n161) );
  AOI22X1 U172 ( .A(\w1<1> ), .B(n91), .C(\w0<1> ), .D(n124), .Y(n160) );
  AOI22X1 U173 ( .A(\w3<2> ), .B(n107), .C(\w2<2> ), .D(n188), .Y(n163) );
  AOI22X1 U174 ( .A(\w1<2> ), .B(n91), .C(\w0<2> ), .D(n124), .Y(n162) );
  AOI22X1 U175 ( .A(\w3<3> ), .B(n107), .C(\w2<3> ), .D(n188), .Y(n165) );
  AOI22X1 U176 ( .A(\w1<3> ), .B(n91), .C(\w0<3> ), .D(n124), .Y(n164) );
  AOI22X1 U177 ( .A(\w3<4> ), .B(n107), .C(\w2<4> ), .D(n188), .Y(n167) );
  AOI22X1 U178 ( .A(\w1<4> ), .B(n91), .C(\w0<4> ), .D(n124), .Y(n166) );
  AOI22X1 U179 ( .A(\w3<5> ), .B(n107), .C(\w2<5> ), .D(n188), .Y(n169) );
  AOI22X1 U180 ( .A(\w1<5> ), .B(n91), .C(\w0<5> ), .D(n124), .Y(n168) );
  AOI22X1 U181 ( .A(\w3<6> ), .B(n107), .C(\w2<6> ), .D(n188), .Y(n171) );
  AOI22X1 U182 ( .A(\w1<6> ), .B(n91), .C(\w0<6> ), .D(n124), .Y(n170) );
  AOI22X1 U183 ( .A(\w3<7> ), .B(n107), .C(\w2<7> ), .D(n188), .Y(n173) );
  AOI22X1 U184 ( .A(\w1<7> ), .B(n91), .C(\w0<7> ), .D(n124), .Y(n172) );
  AOI22X1 U185 ( .A(\w3<8> ), .B(n107), .C(\w2<8> ), .D(n188), .Y(n175) );
  AOI22X1 U186 ( .A(\w1<8> ), .B(n91), .C(\w0<8> ), .D(n124), .Y(n174) );
  AOI22X1 U187 ( .A(\w3<9> ), .B(n107), .C(\w2<9> ), .D(n188), .Y(n177) );
  AOI22X1 U188 ( .A(\w1<9> ), .B(n91), .C(\w0<9> ), .D(n124), .Y(n176) );
  AOI22X1 U189 ( .A(\w3<10> ), .B(n107), .C(\w2<10> ), .D(n188), .Y(n179) );
  AOI22X1 U190 ( .A(\w1<10> ), .B(n91), .C(\w0<10> ), .D(n124), .Y(n178) );
  AOI22X1 U191 ( .A(\w3<11> ), .B(n107), .C(\w2<11> ), .D(n188), .Y(n181) );
  AOI22X1 U192 ( .A(\w1<11> ), .B(n91), .C(\w0<11> ), .D(n124), .Y(n180) );
  AOI22X1 U193 ( .A(\w3<12> ), .B(n107), .C(\w2<12> ), .D(n188), .Y(n183) );
  AOI22X1 U194 ( .A(\w1<12> ), .B(n91), .C(\w0<12> ), .D(n124), .Y(n182) );
  AOI22X1 U195 ( .A(\w3<13> ), .B(n107), .C(\w2<13> ), .D(n188), .Y(n185) );
  AOI22X1 U196 ( .A(\w1<13> ), .B(n91), .C(\w0<13> ), .D(n124), .Y(n184) );
  AOI22X1 U197 ( .A(\w3<14> ), .B(n107), .C(\w2<14> ), .D(n188), .Y(n187) );
  AOI22X1 U198 ( .A(n91), .B(\w1<14> ), .C(\w0<14> ), .D(n124), .Y(n186) );
  AOI22X1 U199 ( .A(\w3<15> ), .B(n107), .C(\w2<15> ), .D(n188), .Y(n191) );
  AOI22X1 U200 ( .A(\w1<15> ), .B(n91), .C(\w0<15> ), .D(n124), .Y(n190) );
endmodule


module four_bank_mem ( clk, rst, createdump, .addr({\addr<15> , \addr<14> , 
        \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> , 
        \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> , 
        \addr<1> , \addr<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        wr, rd, .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), stall, .busy({\busy<3> , \busy<2> , \busy<1> , 
        \busy<0> }), err );
  input clk, rst, createdump, \addr<15> , \addr<14> , \addr<13> , \addr<12> ,
         \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> ,
         \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , wr, rd;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , stall,
         \busy<3> , \busy<2> , \busy<1> , \busy<0> , err;
  wire   n124, \en<3> , \en<2> , \en<1> , \en<0> , \data0_out<15> ,
         \data0_out<14> , \data0_out<13> , \data0_out<12> , \data0_out<11> ,
         \data0_out<10> , \data0_out<9> , \data0_out<8> , \data0_out<7> ,
         \data0_out<6> , \data0_out<5> , \data0_out<4> , \data0_out<3> ,
         \data0_out<2> , \data0_out<1> , \data0_out<0> , err0, \data1_out<15> ,
         \data1_out<14> , \data1_out<13> , \data1_out<12> , \data1_out<11> ,
         \data1_out<10> , \data1_out<9> , \data1_out<8> , \data1_out<7> ,
         \data1_out<6> , \data1_out<5> , \data1_out<4> , \data1_out<3> ,
         \data1_out<2> , \data1_out<1> , \data1_out<0> , err1, \data2_out<15> ,
         \data2_out<14> , \data2_out<13> , \data2_out<12> , \data2_out<11> ,
         \data2_out<10> , \data2_out<9> , \data2_out<8> , \data2_out<7> ,
         \data2_out<6> , \data2_out<5> , \data2_out<4> , \data2_out<3> ,
         \data2_out<2> , \data2_out<1> , \data2_out<0> , err2, \data3_out<15> ,
         \data3_out<14> , \data3_out<13> , \data3_out<12> , \data3_out<11> ,
         \data3_out<10> , \data3_out<9> , \data3_out<8> , \data3_out<7> ,
         \data3_out<6> , \data3_out<5> , \data3_out<4> , \data3_out<3> ,
         \data3_out<2> , \data3_out<1> , \data3_out<0> , err3, \bsy0<3> ,
         \bsy0<2> , \bsy0<1> , \bsy0<0> , \bsy1<3> , \bsy1<2> , \bsy1<1> ,
         \bsy1<0> , \bsy2<3> , \bsy2<2> , \bsy2<1> , \bsy2<0> , n9, n10, n11,
         n13, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n1, n2, n3, n4, n5, n6, n7,
         n8, n12, n14, n15, n17, n18, n19, n21, n55, n57, n59, n61, n63, n65,
         n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n88, n89, n90,
         n91, n92, n93, n94, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119;

  NOR3X1 U9 ( .A(n99), .B(n1), .C(n5), .Y(stall) );
  OAI21X1 U11 ( .A(\addr<1> ), .B(n11), .C(n12), .Y(n10) );
  OAI21X1 U13 ( .A(\addr<1> ), .B(n13), .C(n7), .Y(n9) );
  AOI21X1 U15 ( .A(n21), .B(n16), .C(n99), .Y(n124) );
  NOR3X1 U16 ( .A(err1), .B(err3), .C(err2), .Y(n16) );
  NOR3X1 U18 ( .A(n94), .B(\busy<3> ), .C(n99), .Y(\en<3> ) );
  NOR3X1 U20 ( .A(n92), .B(n99), .C(n119), .Y(\en<2> ) );
  NOR3X1 U22 ( .A(n90), .B(n99), .C(n118), .Y(\en<1> ) );
  NOR3X1 U24 ( .A(n88), .B(\busy<0> ), .C(n99), .Y(\en<0> ) );
  NOR2X1 U28 ( .A(\data3_out<9> ), .B(\data2_out<9> ), .Y(n23) );
  NOR2X1 U29 ( .A(\data1_out<9> ), .B(\data0_out<9> ), .Y(n22) );
  NOR2X1 U31 ( .A(\data3_out<8> ), .B(\data2_out<8> ), .Y(n25) );
  NOR2X1 U32 ( .A(\data1_out<8> ), .B(\data0_out<8> ), .Y(n24) );
  NOR2X1 U34 ( .A(\data3_out<7> ), .B(\data2_out<7> ), .Y(n27) );
  NOR2X1 U35 ( .A(\data1_out<7> ), .B(\data0_out<7> ), .Y(n26) );
  NOR2X1 U37 ( .A(\data3_out<6> ), .B(\data2_out<6> ), .Y(n29) );
  NOR2X1 U38 ( .A(\data1_out<6> ), .B(\data0_out<6> ), .Y(n28) );
  NOR2X1 U40 ( .A(\data3_out<5> ), .B(\data2_out<5> ), .Y(n31) );
  NOR2X1 U41 ( .A(\data1_out<5> ), .B(\data0_out<5> ), .Y(n30) );
  NOR2X1 U43 ( .A(\data3_out<4> ), .B(\data2_out<4> ), .Y(n33) );
  NOR2X1 U44 ( .A(\data1_out<4> ), .B(\data0_out<4> ), .Y(n32) );
  NOR2X1 U46 ( .A(\data3_out<3> ), .B(\data2_out<3> ), .Y(n35) );
  NOR2X1 U47 ( .A(\data1_out<3> ), .B(\data0_out<3> ), .Y(n34) );
  NOR2X1 U49 ( .A(\data3_out<2> ), .B(\data2_out<2> ), .Y(n37) );
  NOR2X1 U50 ( .A(\data1_out<2> ), .B(\data0_out<2> ), .Y(n36) );
  NOR2X1 U52 ( .A(\data3_out<1> ), .B(\data2_out<1> ), .Y(n39) );
  NOR2X1 U53 ( .A(\data1_out<1> ), .B(\data0_out<1> ), .Y(n38) );
  NOR2X1 U55 ( .A(\data3_out<15> ), .B(\data2_out<15> ), .Y(n41) );
  NOR2X1 U56 ( .A(\data1_out<15> ), .B(\data0_out<15> ), .Y(n40) );
  NOR2X1 U58 ( .A(\data3_out<14> ), .B(\data2_out<14> ), .Y(n43) );
  NOR2X1 U59 ( .A(\data1_out<14> ), .B(\data0_out<14> ), .Y(n42) );
  NOR2X1 U61 ( .A(\data3_out<13> ), .B(\data2_out<13> ), .Y(n45) );
  NOR2X1 U62 ( .A(\data1_out<13> ), .B(\data0_out<13> ), .Y(n44) );
  NOR2X1 U64 ( .A(\data3_out<12> ), .B(\data2_out<12> ), .Y(n47) );
  NOR2X1 U65 ( .A(\data1_out<12> ), .B(\data0_out<12> ), .Y(n46) );
  NOR2X1 U67 ( .A(\data3_out<11> ), .B(\data2_out<11> ), .Y(n49) );
  NOR2X1 U68 ( .A(\data1_out<11> ), .B(\data0_out<11> ), .Y(n48) );
  NOR2X1 U70 ( .A(\data3_out<10> ), .B(\data2_out<10> ), .Y(n51) );
  NOR2X1 U71 ( .A(\data1_out<10> ), .B(\data0_out<10> ), .Y(n50) );
  NOR2X1 U73 ( .A(\data3_out<0> ), .B(\data2_out<0> ), .Y(n53) );
  NOR2X1 U74 ( .A(\data1_out<0> ), .B(\data0_out<0> ), .Y(n52) );
  NOR3X1 U75 ( .A(\bsy0<3> ), .B(\bsy2<3> ), .C(\bsy1<3> ), .Y(n54) );
  NOR3X1 U76 ( .A(\bsy0<2> ), .B(\bsy2<2> ), .C(\bsy1<2> ), .Y(n11) );
  NOR3X1 U77 ( .A(\bsy0<1> ), .B(\bsy2<1> ), .C(\bsy1<1> ), .Y(n20) );
  NOR3X1 U78 ( .A(\bsy0<0> ), .B(\bsy2<0> ), .C(\bsy1<0> ), .Y(n13) );
  final_memory_3 m0 ( .data_out({\data0_out<15> , \data0_out<14> , 
        \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> , 
        \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> , 
        \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> , 
        \data0_out<1> , \data0_out<0> }), .err(err0), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<0> ), .create_dump(createdump), .bank_id({1'b0, 
        1'b0}), .clk(clk), .rst(n2) );
  final_memory_2 m1 ( .data_out({\data1_out<15> , \data1_out<14> , 
        \data1_out<13> , \data1_out<12> , \data1_out<11> , \data1_out<10> , 
        \data1_out<9> , \data1_out<8> , \data1_out<7> , \data1_out<6> , 
        \data1_out<5> , \data1_out<4> , \data1_out<3> , \data1_out<2> , 
        \data1_out<1> , \data1_out<0> }), .err(err1), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<1> ), .create_dump(createdump), .bank_id({1'b0, 
        1'b1}), .clk(clk), .rst(n116) );
  final_memory_1 m2 ( .data_out({\data2_out<15> , \data2_out<14> , 
        \data2_out<13> , \data2_out<12> , \data2_out<11> , \data2_out<10> , 
        \data2_out<9> , \data2_out<8> , \data2_out<7> , \data2_out<6> , 
        \data2_out<5> , \data2_out<4> , \data2_out<3> , \data2_out<2> , 
        \data2_out<1> , \data2_out<0> }), .err(err2), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<2> ), .create_dump(createdump), .bank_id({1'b1, 
        1'b0}), .clk(clk), .rst(n1) );
  final_memory_0 m3 ( .data_out({\data3_out<15> , \data3_out<14> , 
        \data3_out<13> , \data3_out<12> , \data3_out<11> , \data3_out<10> , 
        \data3_out<9> , \data3_out<8> , \data3_out<7> , \data3_out<6> , 
        \data3_out<5> , \data3_out<4> , \data3_out<3> , \data3_out<2> , 
        \data3_out<1> , \data3_out<0> }), .err(err3), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<3> ), .create_dump(createdump), .bank_id({1'b1, 
        1'b1}), .clk(clk), .rst(n116) );
  dff_212 \b0[0]  ( .q(\bsy0<0> ), .d(\en<0> ), .clk(clk), .rst(n2) );
  dff_213 \b0[1]  ( .q(\bsy0<1> ), .d(\en<1> ), .clk(clk), .rst(n1) );
  dff_214 \b0[2]  ( .q(\bsy0<2> ), .d(\en<2> ), .clk(clk), .rst(n2) );
  dff_215 \b0[3]  ( .q(\bsy0<3> ), .d(\en<3> ), .clk(clk), .rst(n1) );
  dff_208 \b1[0]  ( .q(\bsy1<0> ), .d(\bsy0<0> ), .clk(clk), .rst(n1) );
  dff_209 \b1[1]  ( .q(\bsy1<1> ), .d(\bsy0<1> ), .clk(clk), .rst(n2) );
  dff_210 \b1[2]  ( .q(\bsy1<2> ), .d(\bsy0<2> ), .clk(clk), .rst(n1) );
  dff_211 \b1[3]  ( .q(\bsy1<3> ), .d(\bsy0<3> ), .clk(clk), .rst(n2) );
  dff_204 \b2[0]  ( .q(\bsy2<0> ), .d(\bsy1<0> ), .clk(clk), .rst(n1) );
  dff_205 \b2[1]  ( .q(\bsy2<1> ), .d(\bsy1<1> ), .clk(clk), .rst(n2) );
  dff_206 \b2[2]  ( .q(\bsy2<2> ), .d(\bsy1<2> ), .clk(clk), .rst(n2) );
  dff_207 \b2[3]  ( .q(\bsy2<3> ), .d(\bsy1<3> ), .clk(clk), .rst(n1) );
  INVX1 U3 ( .A(n54), .Y(\busy<3> ) );
  OR2X1 U4 ( .A(rd), .B(wr), .Y(n98) );
  INVX1 U5 ( .A(n117), .Y(n2) );
  INVX1 U6 ( .A(n117), .Y(n1) );
  AND2X1 U7 ( .A(\addr<1> ), .B(\busy<3> ), .Y(n8) );
  AND2X1 U8 ( .A(\addr<1> ), .B(\busy<1> ), .Y(n6) );
  INVX1 U10 ( .A(n13), .Y(\busy<0> ) );
  AND2X1 U12 ( .A(n3), .B(\addr<1> ), .Y(n93) );
  INVX1 U14 ( .A(n101), .Y(n100) );
  INVX1 U17 ( .A(n103), .Y(n102) );
  INVX1 U19 ( .A(n105), .Y(n104) );
  INVX1 U21 ( .A(\addr<5> ), .Y(n105) );
  INVX1 U23 ( .A(n107), .Y(n106) );
  INVX1 U25 ( .A(\addr<6> ), .Y(n107) );
  INVX1 U26 ( .A(n109), .Y(n108) );
  INVX1 U27 ( .A(\addr<7> ), .Y(n109) );
  INVX1 U30 ( .A(n111), .Y(n110) );
  INVX1 U33 ( .A(\addr<8> ), .Y(n111) );
  INVX1 U36 ( .A(n113), .Y(n112) );
  INVX1 U39 ( .A(\addr<9> ), .Y(n113) );
  INVX1 U42 ( .A(n115), .Y(n114) );
  INVX1 U45 ( .A(\addr<10> ), .Y(n115) );
  OR2X1 U48 ( .A(err0), .B(\addr<0> ), .Y(n19) );
  INVX1 U51 ( .A(n20), .Y(\busy<1> ) );
  INVX1 U54 ( .A(n11), .Y(\busy<2> ) );
  INVX1 U57 ( .A(rst), .Y(n117) );
  INVX1 U60 ( .A(\addr<4> ), .Y(n103) );
  BUFX2 U63 ( .A(\addr<2> ), .Y(n3) );
  OR2X1 U66 ( .A(n15), .B(n18), .Y(n4) );
  INVX1 U69 ( .A(n4), .Y(n5) );
  INVX1 U72 ( .A(n117), .Y(n116) );
  INVX1 U79 ( .A(n6), .Y(n7) );
  INVX1 U80 ( .A(n8), .Y(n12) );
  OR2X1 U81 ( .A(n3), .B(n96), .Y(n14) );
  INVX1 U82 ( .A(n14), .Y(n15) );
  OR2X1 U83 ( .A(n97), .B(n119), .Y(n17) );
  INVX1 U84 ( .A(n17), .Y(n18) );
  INVX1 U85 ( .A(n19), .Y(n21) );
  AND2X2 U86 ( .A(n52), .B(n53), .Y(n55) );
  INVX1 U87 ( .A(n55), .Y(\data_out<0> ) );
  AND2X2 U88 ( .A(n50), .B(n51), .Y(n57) );
  INVX1 U89 ( .A(n57), .Y(\data_out<10> ) );
  AND2X2 U90 ( .A(n48), .B(n49), .Y(n59) );
  INVX1 U91 ( .A(n59), .Y(\data_out<11> ) );
  AND2X2 U92 ( .A(n46), .B(n47), .Y(n61) );
  INVX1 U93 ( .A(n61), .Y(\data_out<12> ) );
  AND2X2 U94 ( .A(n44), .B(n45), .Y(n63) );
  INVX1 U95 ( .A(n63), .Y(\data_out<13> ) );
  AND2X2 U96 ( .A(n42), .B(n43), .Y(n65) );
  INVX1 U97 ( .A(n65), .Y(\data_out<14> ) );
  AND2X2 U98 ( .A(n40), .B(n41), .Y(n67) );
  INVX1 U99 ( .A(n67), .Y(\data_out<15> ) );
  AND2X2 U100 ( .A(n38), .B(n39), .Y(n69) );
  INVX1 U101 ( .A(n69), .Y(\data_out<1> ) );
  AND2X2 U102 ( .A(n36), .B(n37), .Y(n71) );
  INVX1 U103 ( .A(n71), .Y(\data_out<2> ) );
  AND2X2 U104 ( .A(n34), .B(n35), .Y(n73) );
  INVX1 U105 ( .A(n73), .Y(\data_out<3> ) );
  AND2X2 U106 ( .A(n32), .B(n33), .Y(n75) );
  INVX1 U107 ( .A(n75), .Y(\data_out<4> ) );
  AND2X2 U108 ( .A(n30), .B(n31), .Y(n77) );
  INVX1 U109 ( .A(n77), .Y(\data_out<5> ) );
  AND2X2 U110 ( .A(n28), .B(n29), .Y(n79) );
  INVX1 U111 ( .A(n79), .Y(\data_out<6> ) );
  AND2X2 U112 ( .A(n26), .B(n27), .Y(n81) );
  INVX1 U113 ( .A(n81), .Y(\data_out<7> ) );
  AND2X2 U114 ( .A(n24), .B(n25), .Y(n83) );
  INVX1 U115 ( .A(n83), .Y(\data_out<8> ) );
  AND2X2 U116 ( .A(n22), .B(n23), .Y(n85) );
  INVX1 U117 ( .A(n85), .Y(\data_out<9> ) );
  AND2X1 U118 ( .A(n118), .B(n119), .Y(n87) );
  INVX1 U119 ( .A(n87), .Y(n88) );
  AND2X1 U120 ( .A(n20), .B(n119), .Y(n89) );
  INVX1 U121 ( .A(n89), .Y(n90) );
  AND2X1 U122 ( .A(n11), .B(n118), .Y(n91) );
  INVX1 U123 ( .A(n91), .Y(n92) );
  INVX1 U124 ( .A(\addr<1> ), .Y(n118) );
  INVX1 U125 ( .A(n93), .Y(n94) );
  BUFX2 U126 ( .A(n124), .Y(err) );
  INVX1 U127 ( .A(n9), .Y(n96) );
  INVX1 U128 ( .A(n10), .Y(n97) );
  INVX1 U129 ( .A(n3), .Y(n119) );
  INVX1 U130 ( .A(n98), .Y(n99) );
  INVX1 U131 ( .A(\addr<3> ), .Y(n101) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_267 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_266 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_265 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_264 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module mem_system ( .DataOut({\DataOut<15> , \DataOut<14> , \DataOut<13> , 
        \DataOut<12> , \DataOut<11> , \DataOut<10> , \DataOut<9> , 
        \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , 
        \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), Done, Stall, 
        CacheHit, err, .Addr({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> , \Addr<10> , \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , 
        \Addr<5> , \Addr<4> , \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> }), 
    .DataIn({\DataIn<15> , \DataIn<14> , \DataIn<13> , \DataIn<12> , 
        \DataIn<11> , \DataIn<10> , \DataIn<9> , \DataIn<8> , \DataIn<7> , 
        \DataIn<6> , \DataIn<5> , \DataIn<4> , \DataIn<3> , \DataIn<2> , 
        \DataIn<1> , \DataIn<0> }), Rd, Wr, createdump, clk, rst );
  input \Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , \Addr<11> , \Addr<10> ,
         \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , \Addr<5> , \Addr<4> ,
         \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> , \DataIn<15> ,
         \DataIn<14> , \DataIn<13> , \DataIn<12> , \DataIn<11> , \DataIn<10> ,
         \DataIn<9> , \DataIn<8> , \DataIn<7> , \DataIn<6> , \DataIn<5> ,
         \DataIn<4> , \DataIn<3> , \DataIn<2> , \DataIn<1> , \DataIn<0> , Rd,
         Wr, createdump, clk, rst;
  output \DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> ,
         \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> ,
         \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> ,
         \DataOut<2> , \DataOut<1> , \DataOut<0> , Done, Stall, CacheHit, err;
  wire   \CacheTagOut0<4> , \CacheTagOut0<3> , \CacheTagOut0<2> ,
         \CacheTagOut0<1> , \CacheTagOut0<0> , \CacheDataOut0<15> ,
         \CacheDataOut0<14> , \CacheDataOut0<13> , \CacheDataOut0<12> ,
         \CacheDataOut0<11> , \CacheDataOut0<10> , \CacheDataOut0<9> ,
         \CacheDataOut0<8> , \CacheDataOut0<7> , \CacheDataOut0<6> ,
         \CacheDataOut0<5> , \CacheDataOut0<4> , \CacheDataOut0<3> ,
         \CacheDataOut0<2> , \CacheDataOut0<1> , \CacheDataOut0<0> , CacheHit0,
         CacheDirty0, CacheValid0, CacheErr0, Cache0En, \CacheOffset<0> ,
         \CacheDataIn<15> , \CacheDataIn<14> , \CacheDataIn<13> ,
         \CacheDataIn<12> , \CacheDataIn<11> , \CacheDataIn<10> ,
         \CacheDataIn<9> , \CacheDataIn<8> , \CacheDataIn<7> ,
         \CacheDataIn<6> , \CacheDataIn<5> , \CacheDataIn<4> ,
         \CacheDataIn<3> , \CacheDataIn<2> , \CacheDataIn<1> ,
         \CacheDataIn<0> , \CacheTagOut1<4> , \CacheTagOut1<3> ,
         \CacheTagOut1<2> , \CacheTagOut1<1> , \CacheTagOut1<0> ,
         \CacheDataOut1<15> , \CacheDataOut1<14> , \CacheDataOut1<13> ,
         \CacheDataOut1<12> , \CacheDataOut1<11> , \CacheDataOut1<10> ,
         \CacheDataOut1<9> , \CacheDataOut1<8> , \CacheDataOut1<7> ,
         \CacheDataOut1<6> , \CacheDataOut1<5> , \CacheDataOut1<4> ,
         \CacheDataOut1<3> , \CacheDataOut1<2> , \CacheDataOut1<1> ,
         \CacheDataOut1<0> , CacheHit1, CacheDirty1, CacheValid1, CacheErr1,
         Cache1En, \MemDataOut<15> , \MemDataOut<14> , \MemDataOut<13> ,
         \MemDataOut<12> , \MemDataOut<11> , \MemDataOut<10> , \MemDataOut<9> ,
         \MemDataOut<8> , \MemDataOut<7> , \MemDataOut<6> , \MemDataOut<5> ,
         \MemDataOut<4> , \MemDataOut<3> , \MemDataOut<2> , \MemDataOut<1> ,
         \MemDataOut<0> , MemStall, \MemBusy<3> , \MemBusy<2> , \MemBusy<1> ,
         \MemBusy<0> , MemErr, \MemAddr<15> , \MemAddr<14> , \MemAddr<13> ,
         \MemAddr<12> , \MemAddr<11> , MemAddr_2, MemAddr_1, MemWrite, MemRead,
         \next_state<12> , \next_state<11> , \next_state<10> , \next_state<9> ,
         \next_state<8> , next_state_2, next_state_1, \curr_state<12> ,
         \curr_state<11> , \curr_state<10> , \curr_state<9> , \curr_state<8> ,
         \curr_state<7> , \curr_state<6> , \curr_state<5> , \curr_state<4> ,
         \curr_state<3> , \curr_state<2> , \curr_state<1> , \curr_state<0> ,
         Miss, NextCacheUnitSel, CacheUnitSel, NextVictimWay, VictimWay,
         NextCache0En, NextCache1En, \NextReqAddr<15> , \NextReqAddr<14> ,
         \NextReqAddr<13> , \NextReqAddr<12> , \NextReqAddr<11> ,
         \NextReqAddr<2> , \NextReqAddr<1> , \NextReqAddr<0> , \ReqAddr<15> ,
         \ReqAddr<14> , \ReqAddr<13> , \ReqAddr<12> , \ReqAddr<11> ,
         \ReqAddr<10> , \ReqAddr<9> , \ReqAddr<8> , \ReqAddr<7> , \ReqAddr<6> ,
         \ReqAddr<5> , \ReqAddr<4> , \ReqAddr<3> , \ReqAddr<2> , \ReqAddr<1> ,
         \ReqAddr<0> , \NextReqDataIn<15> , \NextReqDataIn<14> ,
         \NextReqDataIn<13> , \NextReqDataIn<12> , \NextReqDataIn<11> ,
         \NextReqDataIn<10> , \NextReqDataIn<9> , \NextReqDataIn<8> ,
         \NextReqDataIn<7> , \NextReqDataIn<6> , \NextReqDataIn<5> ,
         \NextReqDataIn<4> , \NextReqDataIn<3> , \NextReqDataIn<2> ,
         \NextReqDataIn<1> , \NextReqDataIn<0> , \ReqDataIn<15> ,
         \ReqDataIn<14> , \ReqDataIn<13> , \ReqDataIn<12> , \ReqDataIn<11> ,
         \ReqDataIn<10> , \ReqDataIn<9> , \ReqDataIn<8> , \ReqDataIn<7> ,
         \ReqDataIn<6> , \ReqDataIn<5> , \ReqDataIn<4> , \ReqDataIn<3> ,
         \ReqDataIn<2> , \ReqDataIn<1> , \ReqDataIn<0> , ReqRd, ReqWr, n81,
         n84, n88, n89, n93, n94, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n133, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n170, n171, net62999, net104345, net104354, net104374,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n210, n211, n212,
         n213, n214, n215, n216, n217, n220, n221, n223, n225, n226, n228,
         n229, n231, n232, n233, n234, n236, n237, n239, n240, n242, n243,
         n245, n246, n248, n249, n252, n253, n254, n256, n257, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429;

  OAI21X1 U90 ( .A(n323), .B(n391), .C(n81), .Y(\next_state<9> ) );
  NAND2X1 U91 ( .A(\curr_state<9> ), .B(n323), .Y(n81) );
  OAI21X1 U96 ( .A(n323), .B(n397), .C(n84), .Y(\next_state<12> ) );
  NAND2X1 U97 ( .A(\curr_state<12> ), .B(n304), .Y(n84) );
  OAI21X1 U101 ( .A(n323), .B(n396), .C(n272), .Y(\next_state<11> ) );
  OAI21X1 U103 ( .A(n323), .B(n395), .C(n88), .Y(\next_state<10> ) );
  NAND2X1 U104 ( .A(\curr_state<10> ), .B(n323), .Y(n88) );
  NOR3X1 U105 ( .A(CacheErr0), .B(MemErr), .C(CacheErr1), .Y(n89) );
  XNOR2X1 U110 ( .A(VictimWay), .B(n93), .Y(NextVictimWay) );
  NAND2X1 U111 ( .A(\curr_state<0> ), .B(n94), .Y(n93) );
  OAI21X1 U119 ( .A(\curr_state<0> ), .B(n423), .C(n99), .Y(\NextReqDataIn<9> ) );
  NAND2X1 U120 ( .A(\DataIn<9> ), .B(\curr_state<0> ), .Y(n99) );
  OAI21X1 U121 ( .A(\curr_state<0> ), .B(n422), .C(n100), .Y(
        \NextReqDataIn<8> ) );
  NAND2X1 U122 ( .A(\DataIn<8> ), .B(\curr_state<0> ), .Y(n100) );
  OAI21X1 U123 ( .A(\curr_state<0> ), .B(n421), .C(n101), .Y(
        \NextReqDataIn<7> ) );
  NAND2X1 U124 ( .A(\DataIn<7> ), .B(\curr_state<0> ), .Y(n101) );
  OAI21X1 U125 ( .A(\curr_state<0> ), .B(n420), .C(n102), .Y(
        \NextReqDataIn<6> ) );
  NAND2X1 U126 ( .A(\DataIn<6> ), .B(\curr_state<0> ), .Y(n102) );
  OAI21X1 U127 ( .A(\curr_state<0> ), .B(n419), .C(n103), .Y(
        \NextReqDataIn<5> ) );
  NAND2X1 U128 ( .A(\DataIn<5> ), .B(\curr_state<0> ), .Y(n103) );
  OAI21X1 U129 ( .A(\curr_state<0> ), .B(n418), .C(n104), .Y(
        \NextReqDataIn<4> ) );
  NAND2X1 U130 ( .A(\DataIn<4> ), .B(\curr_state<0> ), .Y(n104) );
  OAI21X1 U131 ( .A(\curr_state<0> ), .B(n417), .C(n105), .Y(
        \NextReqDataIn<3> ) );
  NAND2X1 U132 ( .A(\DataIn<3> ), .B(\curr_state<0> ), .Y(n105) );
  OAI21X1 U133 ( .A(\curr_state<0> ), .B(n416), .C(n106), .Y(
        \NextReqDataIn<2> ) );
  NAND2X1 U134 ( .A(\DataIn<2> ), .B(\curr_state<0> ), .Y(n106) );
  OAI21X1 U135 ( .A(\curr_state<0> ), .B(n415), .C(n107), .Y(
        \NextReqDataIn<1> ) );
  NAND2X1 U136 ( .A(\DataIn<1> ), .B(\curr_state<0> ), .Y(n107) );
  OAI21X1 U137 ( .A(\curr_state<0> ), .B(n429), .C(n108), .Y(
        \NextReqDataIn<15> ) );
  NAND2X1 U138 ( .A(\DataIn<15> ), .B(\curr_state<0> ), .Y(n108) );
  OAI21X1 U139 ( .A(\curr_state<0> ), .B(n428), .C(n109), .Y(
        \NextReqDataIn<14> ) );
  NAND2X1 U140 ( .A(\DataIn<14> ), .B(\curr_state<0> ), .Y(n109) );
  OAI21X1 U141 ( .A(\curr_state<0> ), .B(n427), .C(n110), .Y(
        \NextReqDataIn<13> ) );
  NAND2X1 U142 ( .A(\DataIn<13> ), .B(\curr_state<0> ), .Y(n110) );
  OAI21X1 U143 ( .A(\curr_state<0> ), .B(n426), .C(n111), .Y(
        \NextReqDataIn<12> ) );
  NAND2X1 U144 ( .A(\DataIn<12> ), .B(\curr_state<0> ), .Y(n111) );
  OAI21X1 U145 ( .A(\curr_state<0> ), .B(n425), .C(n112), .Y(
        \NextReqDataIn<11> ) );
  NAND2X1 U146 ( .A(\DataIn<11> ), .B(\curr_state<0> ), .Y(n112) );
  OAI21X1 U147 ( .A(\curr_state<0> ), .B(n424), .C(n113), .Y(
        \NextReqDataIn<10> ) );
  NAND2X1 U148 ( .A(\DataIn<10> ), .B(\curr_state<0> ), .Y(n113) );
  OAI21X1 U149 ( .A(\curr_state<0> ), .B(n414), .C(n114), .Y(
        \NextReqDataIn<0> ) );
  NAND2X1 U150 ( .A(\DataIn<0> ), .B(\curr_state<0> ), .Y(n114) );
  AOI22X1 U151 ( .A(\Addr<9> ), .B(\curr_state<0> ), .C(n337), .D(n341), .Y(
        n115) );
  AOI22X1 U152 ( .A(\Addr<8> ), .B(\curr_state<0> ), .C(n335), .D(n341), .Y(
        n116) );
  AOI22X1 U153 ( .A(\Addr<7> ), .B(\curr_state<0> ), .C(n333), .D(n341), .Y(
        n117) );
  AOI22X1 U154 ( .A(\Addr<6> ), .B(\curr_state<0> ), .C(n331), .D(n341), .Y(
        n118) );
  AOI22X1 U155 ( .A(\Addr<5> ), .B(\curr_state<0> ), .C(n329), .D(n341), .Y(
        n119) );
  AOI22X1 U156 ( .A(\Addr<4> ), .B(\curr_state<0> ), .C(n327), .D(n341), .Y(
        n120) );
  AOI22X1 U157 ( .A(\Addr<3> ), .B(\curr_state<0> ), .C(n315), .D(n341), .Y(
        n121) );
  OAI21X1 U158 ( .A(\curr_state<0> ), .B(n376), .C(n122), .Y(\NextReqAddr<2> )
         );
  NAND2X1 U159 ( .A(\Addr<2> ), .B(\curr_state<0> ), .Y(n122) );
  OAI21X1 U160 ( .A(\curr_state<0> ), .B(n400), .C(n123), .Y(\NextReqAddr<1> )
         );
  NAND2X1 U161 ( .A(\Addr<1> ), .B(\curr_state<0> ), .Y(n123) );
  OAI21X1 U162 ( .A(\curr_state<0> ), .B(n413), .C(n124), .Y(\NextReqAddr<15> ) );
  NAND2X1 U163 ( .A(\Addr<15> ), .B(\curr_state<0> ), .Y(n124) );
  OAI21X1 U164 ( .A(\curr_state<0> ), .B(n412), .C(n125), .Y(\NextReqAddr<14> ) );
  NAND2X1 U165 ( .A(\Addr<14> ), .B(\curr_state<0> ), .Y(n125) );
  OAI21X1 U166 ( .A(\curr_state<0> ), .B(n411), .C(n126), .Y(\NextReqAddr<13> ) );
  NAND2X1 U167 ( .A(\Addr<13> ), .B(\curr_state<0> ), .Y(n126) );
  OAI21X1 U168 ( .A(\curr_state<0> ), .B(n410), .C(n127), .Y(\NextReqAddr<12> ) );
  NAND2X1 U169 ( .A(\Addr<12> ), .B(\curr_state<0> ), .Y(n127) );
  OAI21X1 U170 ( .A(\curr_state<0> ), .B(n409), .C(n128), .Y(\NextReqAddr<11> ) );
  NAND2X1 U171 ( .A(\Addr<11> ), .B(\curr_state<0> ), .Y(n128) );
  AOI22X1 U172 ( .A(\Addr<10> ), .B(\curr_state<0> ), .C(n339), .D(n341), .Y(
        n129) );
  OAI21X1 U173 ( .A(\curr_state<0> ), .B(n399), .C(n130), .Y(\NextReqAddr<0> )
         );
  NAND2X1 U174 ( .A(\Addr<0> ), .B(\curr_state<0> ), .Y(n130) );
  OAI21X1 U175 ( .A(\curr_state<1> ), .B(net62999), .C(n261), .Y(
        NextCacheUnitSel) );
  NAND2X1 U178 ( .A(n284), .B(net62999), .Y(NextCache1En) );
  NAND2X1 U179 ( .A(CacheUnitSel), .B(n284), .Y(NextCache0En) );
  NAND3X1 U182 ( .A(n391), .B(n395), .C(n133), .Y(MemWrite) );
  OAI21X1 U186 ( .A(n303), .B(n413), .C(n302), .Y(\MemAddr<15> ) );
  AOI22X1 U187 ( .A(\CacheTagOut0<4> ), .B(n140), .C(\CacheTagOut1<4> ), .D(
        n141), .Y(n139) );
  OAI21X1 U188 ( .A(n303), .B(n412), .C(n301), .Y(\MemAddr<14> ) );
  AOI22X1 U189 ( .A(\CacheTagOut0<3> ), .B(n140), .C(\CacheTagOut1<3> ), .D(
        n141), .Y(n142) );
  OAI21X1 U190 ( .A(n303), .B(n411), .C(n300), .Y(\MemAddr<13> ) );
  AOI22X1 U191 ( .A(\CacheTagOut0<2> ), .B(n140), .C(\CacheTagOut1<2> ), .D(
        n141), .Y(n143) );
  OAI21X1 U192 ( .A(n303), .B(n410), .C(n299), .Y(\MemAddr<12> ) );
  AOI22X1 U193 ( .A(\CacheTagOut0<1> ), .B(n140), .C(\CacheTagOut1<1> ), .D(
        n141), .Y(n144) );
  OAI21X1 U194 ( .A(n303), .B(n409), .C(n298), .Y(\MemAddr<11> ) );
  AOI22X1 U195 ( .A(\CacheTagOut0<0> ), .B(n140), .C(\CacheTagOut1<0> ), .D(
        n141), .Y(n145) );
  NOR2X1 U198 ( .A(\curr_state<3> ), .B(\curr_state<2> ), .Y(n146) );
  NOR3X1 U220 ( .A(n285), .B(n326), .C(n399), .Y(\CacheOffset<0> ) );
  NOR3X1 U222 ( .A(n394), .B(\curr_state<6> ), .C(\curr_state<10> ), .Y(n171)
         );
  cache_cache_id1 c0 ( .enable(Cache0En), .clk(clk), .rst(n324), .createdump(
        createdump), .tag_in({\ReqAddr<15> , \ReqAddr<14> , \ReqAddr<13> , 
        \ReqAddr<12> , \ReqAddr<11> }), .index({n339, n337, n335, n333, n331, 
        n329, \ReqAddr<4> , \ReqAddr<3> }), .offset({n389, n307, 
        \CacheOffset<0> }), .data_in({\CacheDataIn<15> , \CacheDataIn<14> , 
        \CacheDataIn<13> , \CacheDataIn<12> , \CacheDataIn<11> , 
        \CacheDataIn<10> , \CacheDataIn<9> , \CacheDataIn<8> , 
        \CacheDataIn<7> , \CacheDataIn<6> , \CacheDataIn<5> , \CacheDataIn<4> , 
        \CacheDataIn<3> , \CacheDataIn<2> , \CacheDataIn<1> , \CacheDataIn<0> }), .comp(\curr_state<1> ), .write(n212), .valid_in(n263), .tag_out({
        \CacheTagOut0<4> , \CacheTagOut0<3> , \CacheTagOut0<2> , 
        \CacheTagOut0<1> , \CacheTagOut0<0> }), .data_out({\CacheDataOut0<15> , 
        \CacheDataOut0<14> , \CacheDataOut0<13> , \CacheDataOut0<12> , 
        \CacheDataOut0<11> , \CacheDataOut0<10> , \CacheDataOut0<9> , 
        \CacheDataOut0<8> , \CacheDataOut0<7> , \CacheDataOut0<6> , 
        \CacheDataOut0<5> , \CacheDataOut0<4> , \CacheDataOut0<3> , 
        \CacheDataOut0<2> , \CacheDataOut0<1> , \CacheDataOut0<0> }), .hit(
        CacheHit0), .dirty(CacheDirty0), .valid(CacheValid0), .err(CacheErr0)
         );
  cache_cache_id3 c1 ( .enable(Cache1En), .clk(clk), .rst(n324), .createdump(
        createdump), .tag_in({\ReqAddr<15> , \ReqAddr<14> , \ReqAddr<13> , 
        \ReqAddr<12> , \ReqAddr<11> }), .index({n339, n337, n335, n333, n331, 
        n329, \ReqAddr<4> , \ReqAddr<3> }), .offset({n389, n307, 
        \CacheOffset<0> }), .data_in({\CacheDataIn<15> , \CacheDataIn<14> , 
        \CacheDataIn<13> , \CacheDataIn<12> , \CacheDataIn<11> , 
        \CacheDataIn<10> , \CacheDataIn<9> , \CacheDataIn<8> , 
        \CacheDataIn<7> , \CacheDataIn<6> , \CacheDataIn<5> , \CacheDataIn<4> , 
        \CacheDataIn<3> , \CacheDataIn<2> , \CacheDataIn<1> , \CacheDataIn<0> }), .comp(\curr_state<1> ), .write(n392), .valid_in(n263), .tag_out({
        \CacheTagOut1<4> , \CacheTagOut1<3> , \CacheTagOut1<2> , 
        \CacheTagOut1<1> , \CacheTagOut1<0> }), .data_out({\CacheDataOut1<15> , 
        \CacheDataOut1<14> , \CacheDataOut1<13> , \CacheDataOut1<12> , 
        \CacheDataOut1<11> , \CacheDataOut1<10> , \CacheDataOut1<9> , 
        \CacheDataOut1<8> , \CacheDataOut1<7> , \CacheDataOut1<6> , 
        \CacheDataOut1<5> , \CacheDataOut1<4> , \CacheDataOut1<3> , 
        \CacheDataOut1<2> , \CacheDataOut1<1> , \CacheDataOut1<0> }), .hit(
        CacheHit1), .dirty(CacheDirty1), .valid(CacheValid1), .err(CacheErr1)
         );
  four_bank_mem mem ( .clk(clk), .rst(n325), .createdump(createdump), .addr({
        \MemAddr<15> , \MemAddr<14> , \MemAddr<13> , \MemAddr<12> , 
        \MemAddr<11> , n339, n337, n335, n333, n331, n329, n327, n315, 
        MemAddr_2, n306, 1'b0}), .data_in({\DataOut<15> , n202, n217, n201, 
        \DataOut<11> , n211, \DataOut<9> , n210, \DataOut<7> , \DataOut<6> , 
        \DataOut<5> , net104345, \DataOut<3> , n208, \DataOut<1> , n207}), 
        .wr(n287), .rd(n289), .data_out({\MemDataOut<15> , \MemDataOut<14> , 
        \MemDataOut<13> , \MemDataOut<12> , \MemDataOut<11> , \MemDataOut<10> , 
        \MemDataOut<9> , \MemDataOut<8> , \MemDataOut<7> , \MemDataOut<6> , 
        \MemDataOut<5> , \MemDataOut<4> , \MemDataOut<3> , \MemDataOut<2> , 
        \MemDataOut<1> , \MemDataOut<0> }), .stall(MemStall), .busy({
        \MemBusy<3> , \MemBusy<2> , \MemBusy<1> , \MemBusy<0> }), .err(MemErr)
         );
  dff_248 \state[0]  ( .q(\curr_state<0> ), .d(n291), .clk(clk), .rst(1'b0) );
  dff_249 \state[1]  ( .q(\curr_state<1> ), .d(next_state_1), .clk(clk), .rst(
        n326) );
  dff_250 \state[2]  ( .q(\curr_state<2> ), .d(next_state_2), .clk(clk), .rst(
        n324) );
  dff_251 \state[3]  ( .q(\curr_state<3> ), .d(\curr_state<2> ), .clk(clk), 
        .rst(n325) );
  dff_252 \state[4]  ( .q(\curr_state<4> ), .d(\curr_state<3> ), .clk(clk), 
        .rst(n326) );
  dff_253 \state[5]  ( .q(\curr_state<5> ), .d(\curr_state<4> ), .clk(clk), 
        .rst(n325) );
  dff_254 \state[6]  ( .q(\curr_state<6> ), .d(\curr_state<5> ), .clk(clk), 
        .rst(n326) );
  dff_255 \state[7]  ( .q(\curr_state<7> ), .d(\curr_state<6> ), .clk(clk), 
        .rst(n325) );
  dff_256 \state[8]  ( .q(\curr_state<8> ), .d(\next_state<8> ), .clk(clk), 
        .rst(n324) );
  dff_257 \state[9]  ( .q(\curr_state<9> ), .d(\next_state<9> ), .clk(clk), 
        .rst(n326) );
  dff_258 \state[10]  ( .q(\curr_state<10> ), .d(\next_state<10> ), .clk(clk), 
        .rst(n325) );
  dff_259 \state[11]  ( .q(\curr_state<11> ), .d(\next_state<11> ), .clk(clk), 
        .rst(n326) );
  dff_260 \state[12]  ( .q(\curr_state<12> ), .d(\next_state<12> ), .clk(clk), 
        .rst(n325) );
  dff_267 MissReg ( .q(Miss), .d(n280), .clk(clk), .rst(n216) );
  dff_266 UnitSelReg ( .q(CacheUnitSel), .d(NextCacheUnitSel), .clk(clk), 
        .rst(n283) );
  dff_265 VictimWayReg ( .q(VictimWay), .d(NextVictimWay), .clk(clk), .rst(
        n326) );
  dff_264 c0en_reg ( .q(Cache0En), .d(NextCache0En), .clk(clk), .rst(1'b0) );
  dff_263 c1en_reg ( .q(Cache1En), .d(NextCache1En), .clk(clk), .rst(1'b0) );
  dff_232 \AddrReqReg[0]  ( .q(\ReqAddr<0> ), .d(\NextReqAddr<0> ), .clk(clk), 
        .rst(n326) );
  dff_233 \AddrReqReg[1]  ( .q(\ReqAddr<1> ), .d(\NextReqAddr<1> ), .clk(clk), 
        .rst(n325) );
  dff_234 \AddrReqReg[2]  ( .q(\ReqAddr<2> ), .d(\NextReqAddr<2> ), .clk(clk), 
        .rst(n326) );
  dff_235 \AddrReqReg[3]  ( .q(\ReqAddr<3> ), .d(n401), .clk(clk), .rst(n325)
         );
  dff_236 \AddrReqReg[4]  ( .q(\ReqAddr<4> ), .d(n402), .clk(clk), .rst(n326)
         );
  dff_237 \AddrReqReg[5]  ( .q(\ReqAddr<5> ), .d(n403), .clk(clk), .rst(n325)
         );
  dff_238 \AddrReqReg[6]  ( .q(\ReqAddr<6> ), .d(n404), .clk(clk), .rst(n326)
         );
  dff_239 \AddrReqReg[7]  ( .q(\ReqAddr<7> ), .d(n405), .clk(clk), .rst(n325)
         );
  dff_240 \AddrReqReg[8]  ( .q(\ReqAddr<8> ), .d(n406), .clk(clk), .rst(n326)
         );
  dff_241 \AddrReqReg[9]  ( .q(\ReqAddr<9> ), .d(n407), .clk(clk), .rst(n325)
         );
  dff_242 \AddrReqReg[10]  ( .q(\ReqAddr<10> ), .d(n408), .clk(clk), .rst(n326) );
  dff_243 \AddrReqReg[11]  ( .q(\ReqAddr<11> ), .d(\NextReqAddr<11> ), .clk(
        clk), .rst(n325) );
  dff_244 \AddrReqReg[12]  ( .q(\ReqAddr<12> ), .d(\NextReqAddr<12> ), .clk(
        clk), .rst(n326) );
  dff_245 \AddrReqReg[13]  ( .q(\ReqAddr<13> ), .d(\NextReqAddr<13> ), .clk(
        clk), .rst(n325) );
  dff_246 \AddrReqReg[14]  ( .q(\ReqAddr<14> ), .d(\NextReqAddr<14> ), .clk(
        clk), .rst(n326) );
  dff_247 \AddrReqReg[15]  ( .q(\ReqAddr<15> ), .d(\NextReqAddr<15> ), .clk(
        clk), .rst(n325) );
  dff_216 \DataInReqReg[0]  ( .q(\ReqDataIn<0> ), .d(\NextReqDataIn<0> ), 
        .clk(clk), .rst(n325) );
  dff_217 \DataInReqReg[1]  ( .q(\ReqDataIn<1> ), .d(\NextReqDataIn<1> ), 
        .clk(clk), .rst(n326) );
  dff_218 \DataInReqReg[2]  ( .q(\ReqDataIn<2> ), .d(\NextReqDataIn<2> ), 
        .clk(clk), .rst(n325) );
  dff_219 \DataInReqReg[3]  ( .q(\ReqDataIn<3> ), .d(\NextReqDataIn<3> ), 
        .clk(clk), .rst(n326) );
  dff_220 \DataInReqReg[4]  ( .q(\ReqDataIn<4> ), .d(\NextReqDataIn<4> ), 
        .clk(clk), .rst(n325) );
  dff_221 \DataInReqReg[5]  ( .q(\ReqDataIn<5> ), .d(\NextReqDataIn<5> ), 
        .clk(clk), .rst(n326) );
  dff_222 \DataInReqReg[6]  ( .q(\ReqDataIn<6> ), .d(\NextReqDataIn<6> ), 
        .clk(clk), .rst(n325) );
  dff_223 \DataInReqReg[7]  ( .q(\ReqDataIn<7> ), .d(\NextReqDataIn<7> ), 
        .clk(clk), .rst(n326) );
  dff_224 \DataInReqReg[8]  ( .q(\ReqDataIn<8> ), .d(\NextReqDataIn<8> ), 
        .clk(clk), .rst(n325) );
  dff_225 \DataInReqReg[9]  ( .q(\ReqDataIn<9> ), .d(\NextReqDataIn<9> ), 
        .clk(clk), .rst(n326) );
  dff_226 \DataInReqReg[10]  ( .q(\ReqDataIn<10> ), .d(\NextReqDataIn<10> ), 
        .clk(clk), .rst(n325) );
  dff_227 \DataInReqReg[11]  ( .q(\ReqDataIn<11> ), .d(\NextReqDataIn<11> ), 
        .clk(clk), .rst(n326) );
  dff_228 \DataInReqReg[12]  ( .q(\ReqDataIn<12> ), .d(\NextReqDataIn<12> ), 
        .clk(clk), .rst(n325) );
  dff_229 \DataInReqReg[13]  ( .q(\ReqDataIn<13> ), .d(\NextReqDataIn<13> ), 
        .clk(clk), .rst(n326) );
  dff_230 \DataInReqReg[14]  ( .q(\ReqDataIn<14> ), .d(\NextReqDataIn<14> ), 
        .clk(clk), .rst(n325) );
  dff_231 \DataInReqReg[15]  ( .q(\ReqDataIn<15> ), .d(\NextReqDataIn<15> ), 
        .clk(clk), .rst(n326) );
  dff_262 RdReqReg ( .q(ReqRd), .d(n322), .clk(clk), .rst(n324) );
  dff_261 WrReqReg ( .q(ReqWr), .d(n214), .clk(clk), .rst(n324) );
  INVX1 U262 ( .A(\CacheDataOut0<2> ), .Y(n190) );
  AND2X2 U263 ( .A(CacheHit0), .B(n193), .Y(n191) );
  OR2X2 U264 ( .A(n191), .B(n192), .Y(n264) );
  AND2X2 U265 ( .A(n312), .B(n266), .Y(n192) );
  AND2X1 U266 ( .A(CacheValid0), .B(n312), .Y(n193) );
  INVX1 U267 ( .A(\curr_state<8> ), .Y(n391) );
  INVX1 U268 ( .A(\curr_state<9> ), .Y(n395) );
  AND2X1 U269 ( .A(\curr_state<11> ), .B(n323), .Y(n271) );
  INVX1 U270 ( .A(\curr_state<11> ), .Y(n397) );
  INVX1 U271 ( .A(n342), .Y(n326) );
  OR2X1 U272 ( .A(\curr_state<9> ), .B(\curr_state<3> ), .Y(n137) );
  INVX1 U273 ( .A(n386), .Y(n309) );
  BUFX2 U274 ( .A(MemStall), .Y(n323) );
  INVX1 U275 ( .A(VictimWay), .Y(n398) );
  INVX1 U276 ( .A(\ReqAddr<0> ), .Y(n399) );
  INVX1 U277 ( .A(n336), .Y(n335) );
  INVX1 U278 ( .A(\ReqAddr<8> ), .Y(n336) );
  INVX1 U279 ( .A(n338), .Y(n337) );
  INVX1 U280 ( .A(\ReqAddr<9> ), .Y(n338) );
  INVX1 U281 ( .A(n340), .Y(n339) );
  INVX1 U282 ( .A(\ReqAddr<10> ), .Y(n340) );
  INVX1 U283 ( .A(\ReqAddr<11> ), .Y(n409) );
  INVX1 U284 ( .A(\ReqAddr<12> ), .Y(n410) );
  INVX1 U285 ( .A(\ReqAddr<13> ), .Y(n411) );
  INVX1 U286 ( .A(\ReqAddr<14> ), .Y(n412) );
  INVX1 U287 ( .A(\ReqAddr<15> ), .Y(n413) );
  AND2X1 U288 ( .A(n397), .B(n396), .Y(n133) );
  INVX1 U289 ( .A(n94), .Y(n343) );
  INVX1 U290 ( .A(ReqWr), .Y(n354) );
  AND2X1 U291 ( .A(n397), .B(n386), .Y(n374) );
  INVX1 U292 ( .A(n379), .Y(n389) );
  INVX1 U293 ( .A(n355), .Y(\CacheDataIn<0> ) );
  INVX1 U294 ( .A(n356), .Y(\CacheDataIn<1> ) );
  INVX1 U295 ( .A(n357), .Y(\CacheDataIn<2> ) );
  INVX1 U296 ( .A(n358), .Y(\CacheDataIn<3> ) );
  INVX1 U297 ( .A(n359), .Y(\CacheDataIn<4> ) );
  INVX1 U298 ( .A(n360), .Y(\CacheDataIn<5> ) );
  INVX1 U299 ( .A(n361), .Y(\CacheDataIn<6> ) );
  INVX1 U300 ( .A(n362), .Y(\CacheDataIn<7> ) );
  INVX1 U301 ( .A(n364), .Y(\CacheDataIn<9> ) );
  INVX1 U302 ( .A(n363), .Y(\CacheDataIn<8> ) );
  INVX1 U303 ( .A(n365), .Y(\CacheDataIn<10> ) );
  INVX1 U304 ( .A(Wr), .Y(n317) );
  INVX1 U305 ( .A(n381), .Y(n383) );
  INVX1 U306 ( .A(\curr_state<5> ), .Y(n384) );
  INVX1 U307 ( .A(\curr_state<4> ), .Y(n385) );
  AND2X1 U308 ( .A(n303), .B(net62999), .Y(n140) );
  AND2X1 U309 ( .A(n303), .B(CacheUnitSel), .Y(n141) );
  INVX1 U310 ( .A(n366), .Y(\CacheDataIn<11> ) );
  INVX1 U311 ( .A(n367), .Y(\CacheDataIn<12> ) );
  INVX1 U312 ( .A(n368), .Y(\CacheDataIn<13> ) );
  INVX1 U313 ( .A(n369), .Y(\CacheDataIn<14> ) );
  INVX1 U314 ( .A(n370), .Y(\CacheDataIn<15> ) );
  INVX1 U315 ( .A(\curr_state<7> ), .Y(n386) );
  INVX1 U316 ( .A(n89), .Y(err) );
  INVX1 U317 ( .A(n323), .Y(n388) );
  INVX1 U318 ( .A(\ReqAddr<1> ), .Y(n400) );
  AND2X1 U319 ( .A(n292), .B(n280), .Y(n290) );
  MUX2X1 U320 ( .B(n194), .A(net104354), .S(CacheUnitSel), .Y(net104345) );
  INVX1 U321 ( .A(\CacheDataOut0<4> ), .Y(n194) );
  OR2X2 U322 ( .A(n267), .B(n266), .Y(n195) );
  OR2X1 U323 ( .A(n311), .B(n197), .Y(n196) );
  AND2X1 U324 ( .A(n398), .B(n313), .Y(n197) );
  AND2X1 U325 ( .A(n295), .B(n297), .Y(n305) );
  INVX1 U326 ( .A(CacheUnitSel), .Y(net62999) );
  INVX1 U327 ( .A(\curr_state<10> ), .Y(n396) );
  INVX1 U328 ( .A(\ReqAddr<2> ), .Y(n376) );
  INVX1 U329 ( .A(\ReqDataIn<0> ), .Y(n414) );
  INVX1 U330 ( .A(\ReqDataIn<1> ), .Y(n415) );
  INVX1 U331 ( .A(\ReqDataIn<2> ), .Y(n416) );
  INVX1 U332 ( .A(\ReqDataIn<3> ), .Y(n417) );
  INVX1 U333 ( .A(\ReqDataIn<4> ), .Y(n418) );
  INVX1 U334 ( .A(\ReqDataIn<5> ), .Y(n419) );
  INVX1 U335 ( .A(\ReqDataIn<6> ), .Y(n420) );
  INVX1 U336 ( .A(\ReqDataIn<7> ), .Y(n421) );
  INVX1 U337 ( .A(\ReqDataIn<8> ), .Y(n422) );
  INVX1 U338 ( .A(\ReqDataIn<9> ), .Y(n423) );
  INVX1 U339 ( .A(\ReqDataIn<10> ), .Y(n424) );
  INVX1 U340 ( .A(\ReqDataIn<11> ), .Y(n425) );
  INVX1 U341 ( .A(\ReqDataIn<12> ), .Y(n426) );
  INVX1 U342 ( .A(\ReqDataIn<13> ), .Y(n427) );
  INVX1 U343 ( .A(\ReqDataIn<14> ), .Y(n428) );
  INVX1 U344 ( .A(\ReqDataIn<15> ), .Y(n429) );
  MUX2X1 U345 ( .B(CacheDirty1), .A(CacheDirty0), .S(net62999), .Y(n347) );
  AND2X2 U346 ( .A(n320), .B(n318), .Y(n293) );
  INVX1 U347 ( .A(n347), .Y(n348) );
  INVX1 U348 ( .A(\CacheDataOut0<8> ), .Y(n198) );
  INVX1 U349 ( .A(n349), .Y(n351) );
  INVX1 U350 ( .A(\CacheDataOut0<14> ), .Y(n199) );
  INVX1 U351 ( .A(\CacheDataOut0<12> ), .Y(n200) );
  MUX2X1 U352 ( .B(n228), .A(n229), .S(CacheUnitSel), .Y(n201) );
  MUX2X1 U353 ( .B(n236), .A(n237), .S(CacheUnitSel), .Y(n202) );
  INVX1 U354 ( .A(\CacheDataOut0<10> ), .Y(n203) );
  INVX1 U355 ( .A(\CacheDataOut0<4> ), .Y(net104374) );
  INVX1 U356 ( .A(\CacheDataOut0<0> ), .Y(n204) );
  INVX1 U357 ( .A(\CacheDataOut1<13> ), .Y(n205) );
  INVX1 U358 ( .A(\CacheDataOut1<4> ), .Y(net104354) );
  INVX1 U359 ( .A(\CacheDataOut1<2> ), .Y(n206) );
  MUX2X1 U360 ( .B(n225), .A(n226), .S(CacheUnitSel), .Y(n207) );
  MUX2X1 U361 ( .B(n252), .A(n206), .S(CacheUnitSel), .Y(n208) );
  MUX2X1 U362 ( .B(n253), .A(n254), .S(CacheUnitSel), .Y(\DataOut<6> ) );
  MUX2X1 U363 ( .B(n256), .A(n257), .S(CacheUnitSel), .Y(n210) );
  MUX2X1 U364 ( .B(n220), .A(n221), .S(CacheUnitSel), .Y(n211) );
  OAI21X1 U365 ( .A(n394), .B(n354), .C(n262), .Y(n212) );
  INVX4 U366 ( .A(\curr_state<1> ), .Y(n394) );
  INVX1 U367 ( .A(\CacheDataOut0<13> ), .Y(n213) );
  INVX1 U368 ( .A(n328), .Y(n327) );
  BUFX2 U369 ( .A(n316), .Y(n214) );
  MUX2X1 U370 ( .B(n223), .A(n205), .S(CacheUnitSel), .Y(n217) );
  AND2X2 U371 ( .A(n342), .B(n341), .Y(n215) );
  INVX1 U372 ( .A(n215), .Y(n216) );
  INVX1 U373 ( .A(\ReqAddr<4> ), .Y(n328) );
  INVX1 U374 ( .A(\CacheDataOut1<14> ), .Y(n237) );
  INVX1 U375 ( .A(\CacheDataOut1<15> ), .Y(n234) );
  INVX1 U376 ( .A(\CacheDataOut0<10> ), .Y(n220) );
  INVX1 U377 ( .A(\CacheDataOut0<13> ), .Y(n223) );
  INVX1 U378 ( .A(\CacheDataOut0<0> ), .Y(n225) );
  INVX1 U379 ( .A(\CacheDataOut0<12> ), .Y(n228) );
  INVX1 U380 ( .A(\CacheDataOut0<1> ), .Y(n231) );
  INVX1 U381 ( .A(\CacheDataOut0<3> ), .Y(n239) );
  INVX1 U382 ( .A(\CacheDataOut0<5> ), .Y(n242) );
  INVX1 U383 ( .A(\CacheDataOut0<7> ), .Y(n245) );
  INVX1 U384 ( .A(\CacheDataOut0<11> ), .Y(n248) );
  INVX1 U385 ( .A(\CacheDataOut0<2> ), .Y(n252) );
  INVX1 U386 ( .A(\CacheDataOut0<6> ), .Y(n253) );
  INVX1 U387 ( .A(\CacheDataOut0<8> ), .Y(n256) );
  INVX1 U388 ( .A(\CacheDataOut0<9> ), .Y(n259) );
  INVX1 U389 ( .A(\CacheDataOut1<0> ), .Y(n226) );
  INVX1 U390 ( .A(\CacheDataOut1<1> ), .Y(n232) );
  INVX1 U391 ( .A(\CacheDataOut1<3> ), .Y(n240) );
  INVX1 U392 ( .A(\CacheDataOut1<5> ), .Y(n243) );
  INVX1 U393 ( .A(\CacheDataOut1<6> ), .Y(n254) );
  INVX1 U394 ( .A(\CacheDataOut1<7> ), .Y(n246) );
  INVX1 U395 ( .A(\CacheDataOut1<8> ), .Y(n257) );
  INVX1 U396 ( .A(\CacheDataOut1<9> ), .Y(n260) );
  INVX1 U397 ( .A(\CacheDataOut1<10> ), .Y(n221) );
  INVX1 U398 ( .A(\CacheDataOut1<11> ), .Y(n249) );
  INVX1 U399 ( .A(\CacheDataOut1<12> ), .Y(n229) );
  MUX2X1 U400 ( .B(n233), .A(n234), .S(CacheUnitSel), .Y(\DataOut<15> ) );
  INVX1 U401 ( .A(\CacheDataOut0<15> ), .Y(n233) );
  INVX1 U402 ( .A(\CacheDataOut0<14> ), .Y(n236) );
  MUX2X1 U403 ( .B(n203), .A(n221), .S(CacheUnitSel), .Y(\DataOut<10> ) );
  MUX2X1 U404 ( .B(n213), .A(n205), .S(CacheUnitSel), .Y(\DataOut<13> ) );
  MUX2X1 U405 ( .B(n204), .A(n226), .S(CacheUnitSel), .Y(\DataOut<0> ) );
  MUX2X1 U406 ( .B(n200), .A(n229), .S(CacheUnitSel), .Y(\DataOut<12> ) );
  MUX2X1 U407 ( .B(n231), .A(n232), .S(CacheUnitSel), .Y(\DataOut<1> ) );
  MUX2X1 U408 ( .B(n199), .A(n237), .S(CacheUnitSel), .Y(\DataOut<14> ) );
  MUX2X1 U409 ( .B(n239), .A(n240), .S(CacheUnitSel), .Y(\DataOut<3> ) );
  MUX2X1 U410 ( .B(n242), .A(n243), .S(CacheUnitSel), .Y(\DataOut<5> ) );
  MUX2X1 U411 ( .B(n245), .A(n246), .S(CacheUnitSel), .Y(\DataOut<7> ) );
  MUX2X1 U412 ( .B(n248), .A(n249), .S(CacheUnitSel), .Y(\DataOut<11> ) );
  MUX2X1 U413 ( .B(net104374), .A(net104354), .S(CacheUnitSel), .Y(
        \DataOut<4> ) );
  MUX2X1 U414 ( .B(n190), .A(n206), .S(CacheUnitSel), .Y(\DataOut<2> ) );
  INVX2 U415 ( .A(rst), .Y(n342) );
  INVX1 U416 ( .A(\curr_state<1> ), .Y(n311) );
  MUX2X1 U417 ( .B(n198), .A(n257), .S(CacheUnitSel), .Y(\DataOut<8> ) );
  MUX2X1 U418 ( .B(n259), .A(n260), .S(CacheUnitSel), .Y(\DataOut<9> ) );
  INVX1 U419 ( .A(n342), .Y(n325) );
  OR2X1 U420 ( .A(n268), .B(n196), .Y(n261) );
  AND2X2 U421 ( .A(n352), .B(n353), .Y(n262) );
  INVX1 U422 ( .A(n262), .Y(n263) );
  INVX1 U423 ( .A(n264), .Y(n265) );
  AND2X2 U424 ( .A(CacheHit1), .B(CacheValid1), .Y(n266) );
  AND2X2 U425 ( .A(CacheHit0), .B(CacheValid0), .Y(n267) );
  INVX1 U426 ( .A(CacheValid0), .Y(n268) );
  AND2X1 U427 ( .A(n323), .B(\curr_state<8> ), .Y(n269) );
  INVX1 U428 ( .A(n269), .Y(n270) );
  INVX1 U429 ( .A(n271), .Y(n272) );
  AND2X2 U430 ( .A(n308), .B(n320), .Y(n273) );
  INVX1 U431 ( .A(n273), .Y(n274) );
  AND2X2 U432 ( .A(n345), .B(ReqWr), .Y(n275) );
  INVX1 U433 ( .A(n275), .Y(n276) );
  OR2X2 U434 ( .A(n381), .B(\curr_state<7> ), .Y(n277) );
  INVX1 U435 ( .A(n277), .Y(n278) );
  AND2X2 U436 ( .A(\curr_state<1> ), .B(n195), .Y(Done) );
  INVX1 U437 ( .A(Done), .Y(n280) );
  AND2X2 U438 ( .A(\curr_state<1> ), .B(n346), .Y(n281) );
  INVX1 U439 ( .A(n281), .Y(n282) );
  OR2X2 U440 ( .A(n216), .B(\curr_state<1> ), .Y(n283) );
  INVX1 U441 ( .A(n283), .Y(n284) );
  INVX1 U442 ( .A(n372), .Y(n285) );
  INVX1 U443 ( .A(MemWrite), .Y(n286) );
  INVX1 U444 ( .A(n286), .Y(n287) );
  INVX1 U445 ( .A(MemRead), .Y(n288) );
  INVX1 U446 ( .A(n288), .Y(n289) );
  INVX1 U447 ( .A(n290), .Y(n291) );
  AND2X2 U448 ( .A(n342), .B(n344), .Y(n292) );
  OR2X1 U449 ( .A(\MemBusy<0> ), .B(\MemBusy<1> ), .Y(n294) );
  INVX1 U450 ( .A(n294), .Y(n295) );
  OR2X1 U451 ( .A(\MemBusy<2> ), .B(\MemBusy<3> ), .Y(n296) );
  INVX1 U452 ( .A(n296), .Y(n297) );
  BUFX2 U453 ( .A(n145), .Y(n298) );
  BUFX2 U454 ( .A(n144), .Y(n299) );
  BUFX2 U455 ( .A(n143), .Y(n300) );
  BUFX2 U456 ( .A(n142), .Y(n301) );
  BUFX2 U457 ( .A(n139), .Y(n302) );
  INVX1 U458 ( .A(n129), .Y(n408) );
  INVX1 U459 ( .A(n121), .Y(n401) );
  INVX1 U460 ( .A(n120), .Y(n402) );
  INVX1 U461 ( .A(n119), .Y(n403) );
  INVX1 U462 ( .A(n118), .Y(n404) );
  INVX1 U463 ( .A(n117), .Y(n405) );
  INVX1 U464 ( .A(n116), .Y(n406) );
  INVX1 U465 ( .A(n115), .Y(n407) );
  AND2X2 U466 ( .A(n314), .B(n146), .Y(n303) );
  OR2X1 U467 ( .A(Rd), .B(Wr), .Y(n94) );
  INVX1 U468 ( .A(\curr_state<0> ), .Y(n341) );
  INVX1 U469 ( .A(n305), .Y(n304) );
  INVX1 U470 ( .A(n170), .Y(n372) );
  BUFX2 U471 ( .A(MemAddr_1), .Y(n306) );
  BUFX2 U472 ( .A(n390), .Y(n307) );
  NOR2X1 U473 ( .A(n309), .B(n316), .Y(n308) );
  AND2X2 U474 ( .A(n265), .B(n310), .Y(n345) );
  OR2X1 U475 ( .A(n311), .B(n292), .Y(n310) );
  AND2X2 U476 ( .A(\curr_state<1> ), .B(\curr_state<1> ), .Y(n312) );
  BUFX2 U477 ( .A(CacheValid1), .Y(n313) );
  INVX1 U478 ( .A(\curr_state<6> ), .Y(n375) );
  INVX1 U479 ( .A(n263), .Y(n314) );
  INVX1 U480 ( .A(n214), .Y(n318) );
  BUFX2 U481 ( .A(\ReqAddr<3> ), .Y(n315) );
  MUX2X1 U482 ( .B(n317), .A(n276), .S(n341), .Y(n316) );
  MUX2X1 U483 ( .B(Rd), .A(n321), .S(n341), .Y(n319) );
  MUX2X1 U484 ( .B(Rd), .A(n321), .S(n341), .Y(n320) );
  INVX1 U485 ( .A(n319), .Y(n322) );
  AND2X2 U486 ( .A(n345), .B(ReqRd), .Y(n321) );
  INVX1 U487 ( .A(n195), .Y(n346) );
  INVX8 U488 ( .A(n342), .Y(n324) );
  INVX8 U489 ( .A(n330), .Y(n329) );
  INVX8 U490 ( .A(\ReqAddr<5> ), .Y(n330) );
  INVX8 U491 ( .A(n332), .Y(n331) );
  INVX8 U492 ( .A(\ReqAddr<6> ), .Y(n332) );
  INVX8 U493 ( .A(n334), .Y(n333) );
  INVX8 U494 ( .A(\ReqAddr<7> ), .Y(n334) );
  NAND2X1 U495 ( .A(\curr_state<0> ), .B(n343), .Y(n344) );
  OAI21X1 U496 ( .A(n313), .B(CacheValid0), .C(n348), .Y(n349) );
  OAI21X1 U497 ( .A(n282), .B(n349), .C(n270), .Y(\next_state<8> ) );
  NAND2X1 U498 ( .A(\curr_state<12> ), .B(n305), .Y(n350) );
  OAI21X1 U499 ( .A(n282), .B(n351), .C(n350), .Y(next_state_2) );
  OAI21X1 U500 ( .A(n293), .B(n341), .C(n386), .Y(next_state_1) );
  NOR2X1 U501 ( .A(\curr_state<7> ), .B(\curr_state<4> ), .Y(n353) );
  NOR2X1 U502 ( .A(\curr_state<5> ), .B(\curr_state<6> ), .Y(n352) );
  OAI21X1 U503 ( .A(n394), .B(n354), .C(n262), .Y(n392) );
  MUX2X1 U504 ( .B(\MemDataOut<0> ), .A(\ReqDataIn<0> ), .S(n314), .Y(n355) );
  MUX2X1 U505 ( .B(\MemDataOut<1> ), .A(\ReqDataIn<1> ), .S(n314), .Y(n356) );
  MUX2X1 U506 ( .B(\MemDataOut<2> ), .A(\ReqDataIn<2> ), .S(n314), .Y(n357) );
  MUX2X1 U507 ( .B(\MemDataOut<3> ), .A(\ReqDataIn<3> ), .S(n314), .Y(n358) );
  MUX2X1 U508 ( .B(\MemDataOut<4> ), .A(\ReqDataIn<4> ), .S(n314), .Y(n359) );
  MUX2X1 U509 ( .B(\MemDataOut<5> ), .A(\ReqDataIn<5> ), .S(n314), .Y(n360) );
  MUX2X1 U510 ( .B(\MemDataOut<6> ), .A(\ReqDataIn<6> ), .S(n314), .Y(n361) );
  MUX2X1 U511 ( .B(\MemDataOut<7> ), .A(\ReqDataIn<7> ), .S(n314), .Y(n362) );
  MUX2X1 U512 ( .B(\MemDataOut<8> ), .A(\ReqDataIn<8> ), .S(n314), .Y(n363) );
  MUX2X1 U513 ( .B(\MemDataOut<9> ), .A(\ReqDataIn<9> ), .S(n314), .Y(n364) );
  MUX2X1 U514 ( .B(\MemDataOut<10> ), .A(\ReqDataIn<10> ), .S(n314), .Y(n365)
         );
  MUX2X1 U515 ( .B(\MemDataOut<11> ), .A(\ReqDataIn<11> ), .S(n314), .Y(n366)
         );
  MUX2X1 U516 ( .B(\MemDataOut<12> ), .A(\ReqDataIn<12> ), .S(n314), .Y(n367)
         );
  MUX2X1 U517 ( .B(\MemDataOut<13> ), .A(\ReqDataIn<13> ), .S(n314), .Y(n368)
         );
  MUX2X1 U518 ( .B(\MemDataOut<14> ), .A(\ReqDataIn<14> ), .S(n314), .Y(n369)
         );
  MUX2X1 U519 ( .B(\MemDataOut<15> ), .A(\ReqDataIn<15> ), .S(n314), .Y(n370)
         );
  NAND2X1 U520 ( .A(n397), .B(n384), .Y(n381) );
  NAND3X1 U521 ( .A(n171), .B(n395), .C(n278), .Y(n170) );
  AOI21X1 U522 ( .A(n395), .B(n384), .C(\curr_state<6> ), .Y(n371) );
  AOI22X1 U523 ( .A(\ReqAddr<1> ), .B(n372), .C(n371), .D(n396), .Y(n373) );
  AOI21X1 U524 ( .A(n374), .B(n373), .C(n325), .Y(n390) );
  OAI21X1 U525 ( .A(n170), .B(n376), .C(n375), .Y(n378) );
  NAND3X1 U526 ( .A(n396), .B(n397), .C(n386), .Y(n377) );
  OAI21X1 U527 ( .A(n378), .B(n377), .C(n342), .Y(n379) );
  NOR2X1 U528 ( .A(n381), .B(\curr_state<10> ), .Y(n380) );
  AOI21X1 U529 ( .A(n385), .B(n380), .C(n326), .Y(MemAddr_2) );
  NAND3X1 U530 ( .A(n137), .B(n396), .C(n385), .Y(n382) );
  AOI21X1 U531 ( .A(n383), .B(n382), .C(n325), .Y(MemAddr_1) );
  NAND3X1 U532 ( .A(n146), .B(n385), .C(n384), .Y(MemRead) );
  NOR2X1 U533 ( .A(n280), .B(Miss), .Y(CacheHit) );
  MUX2X1 U534 ( .B(n280), .A(n274), .S(\curr_state<0> ), .Y(n387) );
  NAND2X1 U535 ( .A(n388), .B(n387), .Y(Stall) );
endmodule

